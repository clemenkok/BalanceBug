��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�!��
��%Y l�׾�m�F��������2�pς���;����R9���e�����d�dX[|@C�ُs�Z�Ʈ�ڢ4j��s,3��E��.��U[��p�l�o��W&���B٥���Ǫ�6���9n�I�Sr�ˠ�[my�����IUgP�y�W ������Z��ju�䅈;?U�A��y�b&0,j;��oE47%��Le@+h	�Q�}��FQ{�3	��0�}JJ)E����8d���Yh�`�RNňa��Ǆg��	�C�m4���32P��9T�Tu�;?�穴��N��L�����#�����R�w:���ϟ��?͵?f�N�ڪ�i��%O]l� �Juh��GK7�_v��и��}\�9�"�k.���{U���	����?$��#X ��xI�DfG���fU�����o�� U����]8�X��IH����ۙD����V�U3K����Jk;�#��SRv �y܆�^��jH�<�����m֫Ң,�G��0Aa��z�Nw"����#�q/�aV��p���� &ŭ}*�>BNP���åC�S�nd�[�E����c���!y���|�j�O��PZ��k���ӡ�_}Ut�T�C��N����� 8%Ɉ	bgs��j����N�7e鿫A����x��f@��璩)Ӵ�U�k��BZt��cT�2��P�#�9���m�����3uq�&�L�e��2���ց���/�#���&����m�!�䍫q�L9��z�Q����XI�*{�M��Tky��M��%(u6�ިr���9a��k|; m)<�㛒�L�iSH�7ϊ�M{�i*ۄYk���#�$��P��5w����	U�4�Sg��S=��9eg!$}L�}� Kfn����7Q���(����FC����ƕ�$�����<!ʣ�Î,*�[��׵� �b����FluKM��32I5���ڴ߅���r,#�Q�G�O����fRZ�E�x�Ii��]C|�y}3���
�6`��
M�֙L�B���^s2�'�O�	���'J��7j�
 �޼f��$E�家u�W�L�� ��~,xFSW��T<,�)�szss[y��A�srҺNi�Zֱ1x��f��!ܹy���3��<l�l�F��?8m��1R�#|׊���
,�P\���^���/�����#=|�Vb ��)��o��q�R�U�c�����.�W�kP2��\��ŭ�Ȧ�(u�<�sC7�Q��''n��^��ڟ��q�?dں0�-�l�e����j���S4ZK��l�r���J��k4!��M�H�$�`�I��Ƅ�%?d�*�{"�8�.Q�إ�$Y�F�cE�����i�7�#\P+(��y�+Dw�H�\�)�㴶Q�2˃DT���^\C̢�
%v�H��2�N��t$�`5
s�!5Ş����{ �f6�v�Ժ�����g ���D�@�0]�Ѣִ�#1��?�L�fv�,Iz� ��Gg�5]�S��n0��aK�5�������@�j~�"O��T$�j��H���{��)��Ӧg��-C��4/��'0���H2)vɞ҂�r���tl���@�׵)�x����j���B/u1�HZ�%-��V�+�ܼ�vf3q�%0��j`�����^?���:�����I����uo���:���,T� X[�)�J�,(B��PU�J-�˂��X��$�R	_��)�J�݉3��EN)������Gw���YGe�WljC+(��}�)���k��~l(���/"��N�ǅ�'��
P.@�%� �`�����;d�<J@gx	�B�	�S���P�[w��p)���L��]�B����z���ޖa
��9G�]�d[���D�R�Ȇ�O���5U�@��O뺏c���(�e1$ �eJ��I�BH��Þߣ`F�M��k��TO�:=*�@��(���g���!���}��^��8q[ǄY�f�'$#ô����6ݡ#�=I��-$&@����H�b�fNo?u�]F��{8W�va�$@��&a�n�4ݰ��z��gIy@���I[@���H��$Nfvj7������`o��káė����B/�' �(ٲ�5�C�A�ej�Q�Xevd6��(_���(�?@��Ŋ��3y߄�o�y֋�¯̦%���ȳ(�D;5JRx�5�����d����L�������c�^�F�����T.a)~�7p��AH���I'�t(Ez��*�A�Ԍ,�<C���`����0FyHK�/W����-*�f����`6���Ӊ�dlW��j���W���]+Ge�+
���D����2��Mrz��~Y��?�LH���f�z2~�n�x�����g����'�Ng�͒��H�D�D_��{4��Xo)b���l�G:I3�@9-`�sG�"�8����r����y4�`���3f�G��V2I�?-$�	W����ɟ�Q�{\,�(BN��ti[.�S���&�I���%�H�g&�<k��t�u�0[��w����)/j57�?Ա��y�~�Ea�����<���٬䰣�CX��-h3�m-�$�H^2���pi���a����6���d�"��FƤUqo���*B�T���~xY��*��N:I��#�qJ�Kѝ/�%�����qu3�w�|l cJ掑���.+��䟣Q����l�y�1�[6G� ����p)WwO�t]��a��V���?v�-��)(�� �� g���^=���`��G+x48k�@7|�p���l7ĕ����x׵��Ȇ4�(��2��`R��{'���g瀝�գo�ї����o9L�2vs�W���'��b�>��e�\�hf�b��'�P�dM.o�]�$xN �S�Gp9xc���������Usm�HJ�M�op�n�ؑ�N�P��q����Y7
N�B������b�|$���Agj�>tn�1^���r�C�O	���(|�\����x��|�$����K)§\^�jba�.�?��7	�kϸ�$�<c>�
�����-�=pU/���P�!�%]i4" ��b��G1����)؁q�Mj�=I�L�w�8�T)�(>y��T�e檕���T3NQ�p���e}ͼ�9��<6u���b����U)u� K|=�4��,8گD.�� ��1L���z�Q�3rLv�i��	R=ME6O���aG��J�ue*a�p��Jk#��Vc�a=��ܔ����g֊�ޤ�8��y�E�^�K��JcJ�y2�0Sa�H�;�s��?��[�ǋ�3IC&�|��R��V����.�����r3���dR!��`�N���@���5�J�������{�	Uw�ld�H��b�6Đ<��t��_1��|�0g��WqUG|�$(ᢈܨ0�5�z�F��,�m��*�+�[�M��y�;Y�������Ύ�	y@�Mg�Bڦ��T���-�!W+{��ٕ��Tg�}J�A��v.׵��Y�U��4W��8Ɍ�!]�U�]Zyе�^�lB[��h������k4��d��m��;b�)*�F\i�����2�.Y�׉�5�-O��q�'�#$��p0�t�"�l¤Ɍ�a$��i�Bv7b�S�!��|<^=mlɴ}�T�v�Sy��M}8Љl��w�g�,�p�q�a��O͑����"�!�)5=x��uB@f�r,?kl���n�����#�M����9dyQ��˻�������V0�X��@(åmWr0w��g-���"�?8ƻ������E]������>�ED�ع�Z5�
�W���`1�V�����"�Hʊ(�����~l���t<����ZC�`f��<��]�ɦ$�[�֮��$s�(`u/�z�j�"5ˡ�0V�^�V��Ҟ:e�ss�!G��������� 5�-2���t�}5$�<x��i���;�b��3]�>��x_-/7	��ۍWC^PsX�2���X|d{�vXb_�;����>M�[��3'6r��h*�l���R ��E��q���n�5��h�����h�Ќ�Z�K��`�l!B�^YX���̱��*N8���^U
�
��!~�O���H���-^u1˦��_�w�wZm�m�ԳO:LGM|N#-;O�x��,���YѮbr�1$�O����9q�ޭ��xOɧ@��A#g$���}Y�?�è�@��/In� ���@�cƛ��ߗ�6�A�{[$�Hg�����Z��S!hAH�����#�b��8t�z!�7x�-_����Cw�3����^�1����q���4��Ņ�sf�܄ܤ Z-֕�6_iM�^�������V�,<��9yy� 7�Q��Fp!�U$�+
��{�)�@)n=��@��A�rY_g�^U��݃�Lh{KW��8J�A�r�};t� �JS��Ԧ0�B\���VԾ6$�S:7'��x�>�d���	^8ovZ�b��L�k|MIM<�<�"ĳ�pД���x%?T�Ϯ�^fuܔ�v���p>dU��X��ԯ_��D�	�XV�+~�q�	{]Ƕ-���3�LZ��q��<�z�*�;��$��\�\n,�ŠE���־q��u�f�/�6��k$cy�ҙ��D�!��4u���1돹�8�V:2�D���o�������y~dV��`�B��lZ;�^j�6��_�:o5x�֒g��S�{�?�	��d�.|�gB�(��ZF�N����3��"�]�GD�g�xg�������b/�(�������|��+��/��R[���J�\q��6ġ>��_u8QY�z�O��6ˋ���;����L����I,�aE�+��̨l�x(������HLF퍢�V	���t�_��|H�c{���������������tcĮN��Q���������ݱ{[N�=.n5������N�M�3τ���1�A9��;#�?r��P�Z��K�6�HeD��w9�Wo�����R�5����:�+w�[�{�b�Il�H��b@�(��e�ͳ"�92�	�m��( z�Mc'�� M�c-m{�$K��Z����y���}�*iA��)lGU~�*�9�{Q�S#ddv��=�[װ����95[a���3��/%B�BŮ������u�L���Ff�YD�F8�i��=�c��F�Q��E�cSӐ�9,��`��ث���*�����X�h�a;��iM�����)���'�\ah���Hy.ʼ� RH�d�Mv�/z��:k�t'.�T��b)9 $�n�F�	C��t��t�>���D�͖ʏ�%cDt��O��OF� ��TS�3�T�L6i����p��T���c4��ؽ� ���7������T{�_�t�Ь��ڪ�y�N�uP���\�d��o�󒻐���Q�>$��:����2]h-@�3��q��h�-��W�t�Z����B٢x,4�wKb���V���J�l�E�}�֢���sb��qx�Me��QRB�-����W�^wrN��O�G�3&����Vc3�b ��
�Ew6PXJ�xN�o��ٿ�0V�Z�^�Y�v����(Pg��<�D��h�e��~N�JR�H�&H� jv�B��%�g[<al�5�km`�[v~g��8)����4y�4@C9�/���QW�T�˓K<��(�1����৽/AI�����"�C�����D��̖����fA����ꭃ��۲���~f���CE=�-�6�7t���+a˩ab�&�ẗÚo�p���]旊>��R��o�.P��p*�]`���w��y��GK���&~��uC�2�Ҽ>=HOފ$�qu�K��F�,C��C	
����g��C��l��+d1dG��3�\�&?㊡ӽqڣ�W�l�"��W{CFC�d>�/1kk��Zإ�/��0EVR�.�!����@y��?� �t4�e�P���A.�-�a��w�&xS����4rm� e
>-n�:�j�=��,9%���COA�;/�j}ټ9�U>R*�Y2ȩ����E�[-p�b��.h��`y���\~X���8�p9�C�[k?[���C�x�o��in���~au�����+V3n���ә�N���V�������)b��e����K�K�Er��+���َxp�6P�ҏSd`��XS��s�wja�����ѼA�|oH��5y��f���RJ�X5Gr�H���p3�	�i�mL[���(4�;lE�ks�uA<�L�}!��O�[�myq��kX ���N*�{��f���X��j?DA�Y]U��|+�z��O�\x'f

�����%�=�9R �+U�)���@��Sp	��u&�m,.����CD�;rģb����m�jx"ő`f���_�$@G��?�H#���	��%�>�Z%�Ž�	/�_�=+o�K��wŖG��B�v�����K:֨Q�˅����\�cɶQ�j1�����X�S��$�S�v}���G����t��T]�Bs��f��)��گ��T�G֕�����-�������(�5ia'�c���\������O��d܆7����i���*�Rz������9�h5�M_P��o	�Ζ叚\��;Ѝ��|��п����~b8����s�qG�+9u��ױ 5S3�Q{����X�K����k�ѹgX�������t��?����,N'mӃet����V$n�닠gju�:,�����p?��w8V�κ�p4>e�����5/l�E�[��:�p��� ^����A���.�B�uz����/Xe�ur3�j�%?��>����	Zħ]M�$E|S#�ٺy�װ�������Ҙ(7�@����)�F	Kϑ�B�/7�{�UGѴR���姓��n�8#,鉋�6B��T3[6�mp�fdO��T�#���:���R�|b*���ZV���aUs��.�W���� 6���:�{М'�5ن��(%w`P���-�Y)J�ަ��L��UǛ1^��ȩ��QI�)p��w[a(��ǫx�����1-�ز1�X�+��J�|�E��m��Ұ4O�"�������;�YɥG�;�iӁ)6"�e���~k�B���C�>�]mXj"~+��Rdy[�������pWA��4c�ouV�O�2����],F��_O��K��[�)�!�
�H�M���� �5�?`ś��K�h�eY+�m�W6��B|rgT2�F��[����߆h�W��A�*1��VB-���-�Iamƈ,%�|I�H�-PN�E0�,D�L�
�T�%�eW�D��h>ɡ<�����4�� !j+ݨԎE���[���R��:�T�x�Bidxvꌴga�l+j�:�����l��(A1Dë%��jVčWp���}1x�1��O3^�e����٨�0D��oNd��ǘ�b�4�4���ؙ�t	'E�C��}ޒ�>*X�����W}V�?Fn��\k��G�¸��q��6]VG.a-ԫc%!-O�L�������9����p�U�tb����8.2e(�����#��́�0�܎c�H)Y��}�A �*�]ʀ��+��7ݘJ�����sģգ�<���"1�T�,��Ď�][;�etU�_��+�,�̀
�ϓ�F��<īp�L7(�n	�Y$
a[�5F���`��V�Y"\�ybFkQ�X.߲&��+/����^����tk�"TFA�����Hu � t�
E9~fl䞻�, �<�����1��R�EZ�hռEC8�g��Ul��+���|Hio4�9�y�<���[�cvTNOڏ�п�)CL�TZ��[Jr�A�
I:��7��\4}�
��$g[&?v@�z�3���	K�dbyT��c�X�ڮ��y�w�,Gίoz؏:���r= ���V?����8g[3q�'�]9����<js��ИҼ� 2�ڶ� �'Ն"�.-��A-Aq[
;O��"�H�KP,d�/B[��<Qȋ�gWK��:ޞ�n|L��8�<����~�&�J9<��v�0Bt�2w��[��F���d3�&���3݃�ݷv/�IhIfi˭��z��mt����k�E�mf=7etħ�Q����*��2r����"@�3=A�B�t�U�^x �����>d!��w��$C"���Y��Gm�\��&5u� M@m�nZ�3��1��ƚY~V���S�s�p���Ú)�.N2&���ML���$�!Ӄ~\`q����R�Nn.�}u������bc�D��$��~�$�lؾ}`S����n(������S45L�=*��o}5:��PJ��__m]]v0��w ��4o���+:�#���9㆟ө�54�9��7*��, �
�:(p<sC�@��dM���*���ö�D�������[\�x�P�	�|�K�N�hs�D����ws��l�q�q�����F�:�F�Y�`7 � �y�`{N�w�(T��l���_�P_R��ۍ���7��&���:�K�o!
��Q��<}�@}L��{��W�����0߱g.�o7�p�.��ļXĸ�v��j��1���a_�q���_�ÃB>ڼe�$�0�7<�m�^<����G�a%���&��hN!h��f���e����: ��yr3�6ioI<;_�%���A"�����:7i[��P���=���_C���H���"e��|.�	C�w��Gu��;@<�ZPÆX�NZbP�Q�K8��
����	oE��Z�G��1��U�rsj�i�6aoBy��U�tK珇@��-�;n�}�� `߁ħ��>}轭��Ӹڵ;7�u�N��pY��/wu<nB�O���)rp���l�f�d��-�qڠ^�h1����/��q8\���8l6;�KZo�'0 �Gb��ČKy����̕o$o�)YM�4�\pc�F.��b��C^�[j�y��zQGօ�.0m��e�<cZ�G��t�9mD��P_sCQ<��
�c���4��l�V�઻Z�zY�S��[]�r6G�e `I�ڲ;��qۗ�>�~��7�\Wʙ_�˾������~�j�xe$�ɜfc�H�߲q�gy=/�I�|�5 �����z�.�W&��;�V���Q�%�7�H&�\��(ڌ�_��
m�������.�]3��C�8լ��E�P�7���@��;9J"1����tP�lb�F{ V�īt ��ܺ]��>5�ƚ��g�垊�ȇ�B�&�,��عG��4���J����"2�C�ĉ���o0A<�"��I�@r�0+����5��~�ɑ@��J;Xײ�72�5"���ٞc6%�-�x�y�")ce��ѬƲ��	�}��.�4�ޟ�Ӏy Tx�W؃p�(�.L��fa�Z�ۢ�3��I���O�����'�8�#��?����),�b6Yx��"n���eÕh���p	�c�7�m��S�;��8��D�K��]�M�a�G�@E�U:I�D���2���1�v��q�n!Y0�gG�&�r&��� � �]wI+�1%.�߹�w�ػ�n,i������#<��!�E�\�y�U�;$<֗�k��`b�����`�ե_�U��&˨1̻$��e)��Ʃ���\K;㨞{�*݂n]����^jP/晔��]?@��;�k����Ĺ	�Y��'���J��t��*}�~	�w3s�[�x�]�G1w��q�f`r�2� W f����K� ��XdH��0M��!!F�s�va㸘�l9�����nW �b��D��n���X��X9x*>j�B(%	mB�3ȲJ�����:�8{�F�h�͖d�pp(U�"�TD��4�S�#Un�u�mI�aM�<*��_�z��?��ef0����@(��/��J�Dy��ZqJ�,"���-�t8��s2���/������{��v+�/��bpC/�6��y���&��e�h��q'S3t�	�MN+i3��$k5�u���5
����)bPʩ��"et�^s|6����Wz������U���=�Q�њ���S�<X��m�^��H�)cA7y��4�	�?�x(գ�:�˶��H�;�;G�{q�v]��G6a��J�aƞ���L0��b�j���	n�I��%_I�x�R����`1�hI�Xz ��;��e!�p����5�7�:�p��U8���x������9.��xIR�7�\ғ�H�d{��,����&�a��LOBAR���\Q���s��/��{�X����{>2L�I�ya$q8�Tne��v�f�??]��ャeJ�s�cA�b����{��*��D�� pf؁G:�Ǧ�A�P�7�N9c��`��;������$7q�A6g�F�������M�E��L]�}��v��4WB�Gbǵ4����2�)�~��9]|�B�Gj���_t���@Ƹ�O$$[��4d+�'z0���bG�g��SN�e����0��lH|�ʹ�1�!���솜� ^�Ѕf��|��/`�{92�dl������"]/c�@�^j��=�T���E����?.=�~��Y���V:p�=�-��L�w�8D����\*>2҇����+��#�I�t=+�gб�S�(m�%[�x�4˄-\�"
؊�>�`��ע=A$�ڠDG�*Q0q�^hnA9#�E��7�������X�[���ܶ"o\T{���	D�����2����"�3��3�E+�m����Z�|؊�t��M
>�c��7>���������CL�Q�~P����)ꘖ~��@Q=�Fi��"����{QC6�Hbmw	�0R�N~�������P寔K�f���v𙭪�pP9�΍3�6)C�i�HO%�j9tЙsJ�yu1���6��U\�� ٦��L[�%����÷wCA�A�vm�� ]�`�`K�%)瓤�xNJ��)D,ᒮC�^Ah��+l��)�$�Q������~���/��[n�&GdA�bc���h��&�tպ�~����(��ԪR��^�N�Y��ssz���S<���_�:N×U��G��t���쭴���0�
���;� �b~�X��@v���V����rV��2Z�}��=���Vab��D�X&>���������L�P���̵�"!t�^yVz��]�2�KQ}�?W��a���;e�͞m}�%����Y���+�l�/.�� �0��3��R2V���r��`֌��8ڎ{5�b�F�������Ӫ�yxUL6x$����J��P���>�kB�*#R�S�Fg��K��
���e_��'�J�8z7X>	I5qI�9r;* o��$�+ʠA�&T��F�H��|eP��XQ�psE�> #d�覒�L����sJ*EE;#�����nPAymx�TӉeK��7-vīШX�زB���C^���{&?��]�i�ku*VIV��KD$��ͩ�Ҍ����>��e�� ������vQgad~��pNojN v 6ka����is�z�Ʃ��|fO(����dw��I�5�s�F\d[O]��`)�q��
���|��B31�#�;c���Hwpd�J��`�.�@m���m��y�%	��9CՁ�H���dJ�?�Z�G�^@���̧7Rjm�Kס]��!��5�8χՙ��sT�V&;qH>�]���j�XW_n��>��.H���7y������da L�xgc�
ł�����,��%Y 4I}� �_G!���W �RLY_".�?���9Z�dL�LL���4��DO7����ۃ�P�k�.|��|	��(��mu5�a3���~�J����� '�s K=d���a�;X�܎ �`8A�i��e�-j��4"�^ϰ��65��)��
����ca������F2�eٸ��|yv�����v6}"7=F^�C���u(Lya�u3ʏ��.l%"X�����L��"��`�Ю>�o)2����������'0c/8
ǢGB�"1<�.�.C|��fU�-��q��2�LU�$j��sRդ4�vd��})8b�<�'����yo*�f��t��hx��Ԕ:]o�1gcӸ?ha"��;Z�4�	;�p�m�|޻�W=K{[sRXֲ8���v��!�0r�����/��-�v�SdIޝ��گ[|���{�F� ��0��)��ޓ� ��w�H��ggeBR�*h���(r��Β�3��.��<���+��*��i�s�8y�6�Wϛ7ЦMV3���o�kH��0J~��QS]��Ǌ��E1�r�)9��=�[O��ԠY��*~��@���PϺE���5�o��<>s��	����F�c-�]J �4.<&\O��k���7�5�UY�l���
Pc��y��7�t�T�V�P��/���M�J bc\�]�9�!o��yn�V��'j���3�zJ�]4�>���.�7Y~�	GTQ��HA-�W�TR� s�6���bo�_��rCJ����퐭	��WI �gk�}�&{�Bi�2K�9!��ONunU�щ�d��$c��zа-t��` �㔳���|�i0�#�o �c�63�M; �O��K�t�X���֫�u�L(͹P6��0�0�S�\�6���6�]Xg:�;�!F ?�ow��F�dt��<��V'�R`�B2���������f�o���V[��(�(��۷��k��Dɱ{�,'i\n���`bFK����W�X�ξ0 ��ɤPmRg�a!��3>�ޏkd�������?���t	�_s��~��J��������T5iL��K����S�YpAuA�i5i���2��|�0�3Ȋo�!��Gra��,F��}+�<�;��lo�Ѿ�}�N�z��]���&���JV+���4yy���EB^��#�m̔����܆�s-)�, P�P�R��OY>һ�5�-�Ŋ�>����|�����l6vI�Ҝ��71�a|��4��e�u�H�>��޸{)H6e�L�,�Jt��0D:�D��i�5+�E^�@�pp�[,�OY���X�!9'@��\������g<"�]8�A����M̋��أ��!.?�&j�Ǆ*T�3�?�Q
�ŗ"d�U��9eNp=;`���K�)'�鏕Y׌�.�l�����R��ʦ_$ca*��r���y����p�d���#F�[��$�౩�+����O�rbԖa��l��X|�g�)���W�%��Y����;��=pϔxy�:mK=�r�|u��>P����FH6@���˩Χ{�T���ݞ/�Pq�M1"q�N�Y��񸥨_�m�2���KZ�P����RY)Jn�P�
G;������r���Tci���"F;yܴ��^on#^�Q�K]�H'4g��:c�&'���-P�[��#��H��ݛ͓
��χ��W��/n}�l�_�X�5r�`	����"x�|���S�X��G�]�ƿ�.�*�sB�a��!��"X�Y:J�9�5L�"���=\ŕ������_if�r��KF��l�&R��9ߤ����_K\���c�+�r��Y���v�� @����´A��������E�1\@�>lW1��I�D�g��$C�A+[��]��?O�:���3��0��;�YCL�ΘEQ��6\�T��MX� ̩4��h�H�{��z{nh�$�s;��JDg=ᜑ|�v�}��j�6J��ʛ���y=����Nz� �
�b{�L�7���Mr�r {Bmm=��ҷW��rA�-�C]�YvR�4�'��}�}��ɷSY�]���Ld��^����sʕ����)J>�K&���M�<j�t�:��P��{�%����z�<L�����J>�h����@��+ˉ��0a�=�-��[�B,u�t.�;L�-X�Cp���0έH!|�~��Rx�(0_�N��$��\��~ʇ�kI x�/���f0��8B������Ò���Sv���y� ���>�x�n`���գ<�൦�� 4�f����Ӗ����t)A�A����d�;1�N�Dx�>�7���|� �� �&6_��R�O�D
�s l�ϯ\q fB;�j����{��Q�u�M�χ/�j��~�|���{�����ɘ�C'�din���e���n��N]d1� �;�d��Ү�L�i2;#B����&��Y��+��8<��y�([���!+OA?�2X��O�p��gO��i�P�Nã�q�� D�6�o�ߴ)�}��I�ïږ�e�q7B~H��k"vEAU����'71��a���]j1�,����_�9��+ٲ\/"g���L�;{Xx����1��TR���p�@B��W��` ����'B��|o�6����5`/~����:e���H���O9eYg�/�c~/�O.W��9�l-�9���7�̍�oW�?_������53��NF���T���虾1��2�kt0���,u��[{6��V�t/��D!�7��a�4e��%�����Cl���Z��U�㎙�RT��KX{�Z��{�	�֭����m�Ƶ m�9��)wG�*�����r��^����&��w:���+���翼Ȅ�׊��Rz��c����L=T�<�����P½y@�\�۱\b�9B@\�[��"�A���_�e��!Ҵ[p��}�Qk�W���W�=���(���������d�/������38�8t ��o�H,�g�V"]�y�o@�|�6��A�\�q���q~p���~,�£w�����h�!��Ğ��0���H����i1��ة�7���7<K����c�������0 kh�����\��2�d�M���83:��W�Âh�k��_0�iq�g�L(ar���<Y_���&�Ì�k"�В�y�<�#�wi�N$��Y��~	��s�׽�W�����v$u�>!,�>v��T�*�He�g�8_��ͦ����.T�nXޜ}����p>Y��:�b����lI�<������Y(�b�F2��zb��f�����ā�粲��1�}
@�{��4�lA<x{�>�7%}�彰ɵn��T�&4t�$T+�F󻥺�������0��4v����k�~@�n�e�@;��r:�D4?/�t�X��y�LXx���e?�d*���jl��v�-$�$�#����h@�G0�F�pd4+��*:j?�fGn��ˣ�w�0@lC����x���)ZƓ�M�<q]a�J�]��_��B,l|�J�)E[�YCxfT�*l샯�[yi�UX�`����h+�G��?2ڲ�_���g�!)s�2F=Uh}�+ ��e0��F�R��ۍ���M=R�<�m�nW�^�f=�)��ɷ`o�X�4^����S�����e��뻂�����Џ�g�]������U�E4�}48��Ww)�m�+pRIR�~d�����D�_I�
��D?���U��8�Y"-+���O��_�G��K)wBP+�Ĩ�G�k��n�ޏN����5M�2�&�x�d8:W�� �#�cH�ߧ�@b��'|���&<�8�v�LXf,��58dB�ႌ��n�H�|P�����@w�d ri)���y�-���i^5��k�jV���&v�q��l��Am�\=�MS\�9���Ν �N=�t�(�H��:l��������d� »*!
��%����i)�w.)03Q��\��ܽͺ%�k'�Ј)x��:�H�E9B��M��[�^`������2}�4�avأ�F9I������:J���5i�.y{%6��PC�hZ/�[=%�m4�'�z��< ���K�򚊒�2��y&1ݜ�;�8I������7���F���y��yu'}��3̫�n�7��-�ܧ�(���GGH� �Y�,(7*����@ɘs>�fn"���(�6���^F���B�q�0ᬶ�g0q�~q�������*�lq����h�l�E�e�\*��p�`�A����E�з6w���Qn|���GZ#蜈�ތ4tB���mQ��ރS������\i^��b�l� 0t��-�lT�&�-�E�d������FE۵�.!r�:C�4y&ڀ�O��6+�خk� ���^d���@C�qz8��`'V�eTˤ�ĭ�����8W3K����)�>�9pC(�<<�
����I�A�\�j�z�G��N ����@'�\��*R��J"gf�X	�	H�u�sL3b��b���Z=�л,�x>=�)\��}����n�k	6�eɟ�T���	}"
�3s	�"t�~&�jjfK<��x��R����ַ��譩bt��� ��r����̕��m�W�47�124Qs����u2��h[$=����+	�)��������#&,N�v}����aqu��"���<`HKz=�ϗ�l�O��u���s�~��K�L^N�k��T&���A�D���%������V} ���&��l
���J�AcE;@�7��U�M��/)�}��'NW[U����q��m��8Y�&����(��?��&�=��e?v���2^��S�&�����eG����N�#="�'x�C�
�u0�r�C�{�����-�2�/�C�=;��b �"�Ŗ
l�ڽ���eր̽�Olb&'�@C%b��[9d�v8��e����;�������m�� �4Xl�G�g�FLZѺY��=��(D׾�I�U�s�FjXp�34@F�����Y�_�C[�cy��ڼ�u�z�Fl�~!��Y�/K��6p�R?���=�]d��naI�����.�x�~7f���eu9K�6�Z��]"A�TåV����;���PFhzG�G0�;C���W���*�ٛ�t�»=��g�eyuh��z*�zk��h΅��K�(D0�R�����~�Ӏ���nk���"��'S$��kO�'PX���g�z=	\�S9��vFT�����l�g������ˢ��[�FG��s��e����3�6sݼ �i^L�5(�R<�9�x]�'�d+jҚM�����(ߖFa���`Aw	��NK�� ӫ�Vb[2�ޤV�1E?�1?���C�Q�ch�iK�~��P���-WT����f9v���e�l��T+� ��TNlP����=�:<����f=�F 7P)(g��$�H@���4�����W�O��i�D,w�+�a|,x�]�hyܲf�kX��h8�������A]~	;��u�Xp�4�V�~T�^����k���W5[O)xi�b���60?aH�j9�\��=�C���Ҁ�NT��d�v�M�`�5%��|{��:'�~�]IT�5l;��[�c��O�f���P�C�n�]�o�ˇۍxz,�e�}u�g���+F�)'���n�#��l�L]��+���o� Ť^��gC<30�zY�����w5��J��y�2��O$2�@�yԚ�GD�&� ��ty�'
7����bE��@0'%�M!�~#�E8��_������(���lޔ�a��G����� ��k��r��>���p�T�l8ߟ��~u�^�
��y�\��}�+���#��	H%�xQր�axUJ�k@{�2e�x!n��,������	8�_, ��UQg�,<¹B�W��#a_S���04R�9x�p� �|Sӥ�x�!Ϋi��H|�D���Ɨ�Pr�59}� �!%�,�L�Y<5��,��������V��Ι���5P�"JF����Y-��	О�Ѫ��L�O;C劣��6�i4Sʯ�N��?�n���\�$n����[��a��M9�#̱�+���`8��.�����k��Z�"+�^��7jp8�hr��G�ux|���f�s����T12n�𱹭�ڳH�(�"N}�EݨOu���WC#;�v��������lw۱r�߾*b�-��S��4 )"�ԫ;��(V
`v~�od@*��mM���MU�G�s�6ӫ�n�IR�u�7��mϝ����%���T_&%�6I�;��[�sK�zX�C#���v��^�x�����9W��U��=o`��\A�l�!b�Jz��*�X|tJM�5^���5�(y�qŁ���z!5��Y��<	�	�6�W�l�ZC��.+'ɝr�@�Rn���p��Y<$\p~���	�ᾮ)�9�iq��kn�9�*�]��an�������OUHO�OY!x�l�U�7��,뤹9��qޫ{o��>�µם��Y�WT,5��/�֕�#���ƴ-�-V���>�f`)�%oӪ�R%�蘃�u˄oY���Bt���dިEޮ�lY�/u����o����=ɏ�R�΅���sht���<���~�E�~V��r<���@�"�[	.���c���.(�Mr)�a5�,g 4�z�d�/b!*8�[u�I@t�����lt�#�x��"aH�O��d��;����9JȞ��k�2�������⑮�\MU��$�=��|OkYČ{{�/�,�P�2h^��?�2T�@I�@IϘת8������KdE�S���������3L3@��ݚ+�� �k���v�:��>��ͪo�ş:)��$TV�J�u�E�lS� �����-�g�?�)'晔�ǯ�����gXl�`ϱ�������!�$�ˀtg(xa}�|�w8a�䂫�S%!Dݨ�5�(����̊�R����x�D-�G�,�Իc������$1�kk�h�7�G�Rԗ��P݀�/\_"4\���E�+e?��a��~�!~K����=�*��=�_j���8l�>]���bA��b�6�Q6�\SI·�;n�e�FH�� ��l�����;�AQ�$�V�[O�Vw��⁹]�Z¦�U�Wut@��%�g4��4)Ռ�UT�<��f��N6�X�¶_�.����ĉyө�B�� ӥӕN@F0�;�Q��D|�;�O�l.!�6!Ep��a���B]�f��`�Q����O��3&>��N��B�����<(w��H����G�Q�,���ܶ[����h�-���~N5U�<LԺ��~��`-!/X����V��0��GQ����Q�D�l�V뿗�a��%�iD�V|�o74��A�$���a�{�-@g"��}�~wt�]�Д\f1�<,o��\���������e�@�5��E����w 2�|t�ݓ�49X#�%?5i�5S�y��f����YY��m�v�Ci=ȏ���G�.��[�g�}�K�0�������d
�7��=!�����A`A����瘪�AI�\$A��B���UO��.B�e�����i2�iCwy�p���=�F�\�l����~sǢ0Xq��v�ݽ�zmHrO�F��K��h��J��e"]x�<6\�����BJ�䊕{u*<�6����7#�*����������&ƪ�y����5���Ȳ��>��h��V͛l�I3^��"L����	�U��m���M�雜�Dl�������^����f�˞��b)� �ujΝ�i��a���������'nfgE��~�U����bm���'I 6�vV���"M��v5�d�	[ԯ�=�ԥ��M�@�����^Ĳ�8as��~�m�pq2]�=��*k���zKa�4w�"������mP2���B'�X�oT�%����Z�̭o��&�$ܾ���DP?M�����KO������o9�(�+�<]�,�l	��=} �ǖ �LːNT�g�5*�#9jeK&#�m�K-�PX�U�,�c��?O^�!�ҌA#��B�V:ʬ��%�.�jO:ћ�o��r�O����+��t3��t��@�$�,�;V���C_��g��VMq��Ș�u�g��&�_��,7C`��/�/��x�&�|��8�$!4����$�1�?�2梄HY~F!)�]�/�NsOs�h�,i��åe�s�N��pa�
�G�m�u?؝��~��PՆj,eP���� ���Q�i��Vg��t/����7�D�L�^e:��g����xd8�U�����S�n��o"��1-���NB�Fd����S�o�"YH�.�� ��r��S��Ķ�Qw��c~c����M��ecAR�x�ەk��Q���dX�I�Q�mP m���;����>��: 0,ʎ���(qVZ?�Jkj�w�E���� ,��������6Z����i��g-�r�r��h�'�)I�By�g�X�Q�rel�Iz�TT�P5:���C�̸���`��h$<FV��+�(�p"-=,�ATb��ҥ4_�]���oK��a��+�wC�K&�3�P"ZK8A- ����ڎ<2��9��[H�����i݉결`�:��k�@�?�~/7I�P�ܻ�[���h�̿s#��x�H.*b�C�J�����i�+��yb}��i]\jHc��~��I ����H�Kr� �*�1�mD{�`�B$�}��Xu�	��I%B��`�4Jwhx���A(�u3���f�Sy���2�?�'7�G�MWͻ�++��c�VIaY�����t�o�W	&�(+�_%�B�/�FT�$��:�$�t!�5������)�_L��@K���S4�b��2B��mL�V����cj�]Q��מ�YsE�hӭ��'��[�i�%�KQ֭#3�lUV ������R��Gyg���@�ib/�X�Sʡ5��7"��Jݓ$�|~�~�"�S�D�E��(�	a�E�����P��yD��o�����3��&`�]κ5��T�Q����I�|r;ְ�r2)�EV(تE�K���V�/�I��ӺO"�Y�ǐ0���|�&-+-M\��J'�r�K��_�I������C��)�~�*��wl���b ��{h�RH''HCsm����@�Yj2��j��B����UX֋/��H���/i��S�V�(�O#� mYkܕ��)W�5���ƿ��Z��~T�s�ˀ3ЂO�p��Yܣ���gE'��O?����:�� �~�"2�����2K�'jch�A���5����*].č��'J�?T��mT��#�cs�\6G;�A׊��^��,S��_�w�E��s�؀��St�w1��f%s�	6xL��j	�`@F�U��~�$w�;���#�P��I֎Ұ��������!fT1;�p_���v`�A1(�g4<�z�Rj%k��� ��C4�rɝ�3�|�����nj�gd��	e�!��׮���6C��/��S�n��N��`��B�t�dE���D��$��>����Iv���?����������� ������r�L���F�S���x0���:��nF@)[�%2�� �e�g�i5f�o2V������Y�RR�QۇUh��!;3$�@�s\	p/E��\UZ�l�
1a����X��K��l���#v���A]9����aY��b�gW����=�
��ˑ�Qu�1�O(�w$ӆ��7W.}�c�C�L�����&"a�Fm��T�&�X�t7B}���Qn���\ h�����Г�4�F��S:㉄ݏ����-��Q���H����Nf�'�x���$7����ҁ�pݲ�\ֲ ��K #� ޳�� {Z��i�<Cs�~J�Q�
�ч��k���s�=�r�\��"��V�g���Pgzk�,��S��e�^�H�X�gߊۜ_t�sV�SY�}�}6aP(�z
S%.��n���r�<;�RyC2�q��K��/�8aM�kx�h�E�8,�O����A9^� ��St�7�\I�V�i�Ř.��Bj�XH�����������~h<ڗ���޵}�Yr��;������CtG�(�:�c��\��Ei-���<,��nΖA��k�-��q�q��,����W�%���[��"�fB
�f�(��J�ɀ<A����#�j�^w�6FR�B�܇���u���W#��-��.�З��+��U���l��_���ם�7�rk���,�K$fS�y?�f��\�h��{��U�ѓ��\�'���Y�M�p����hU~?�6�?� ��(9�HdK�����<x�ͱ�99�$�%���t@���G��k���%'�.6�
-�<5�b�-�j&���?O���Yyh���6��Z3c�k���R&I`����3�[=g�� ����շ�g��1��Q�ҕ1g��^�h3j�B0a���rY�$	�ź�p,Š?_�'�=�ʙz�p?���V�e�gA#$[�σ�)館��$�	vy+7$$Yu$��FU��J�N�஧܋�*�ml9�g~�.i5e�{���ܮTi�oX��&�J����.ǶGQO3��M��d�}S�u=E��qdT|<�5ꊗu�Q�N)��b��ʮc�4���Gm'�w��zk/��W����Q4;̜Q��P	ޕ���?��z�읜N�,a���/��;�d���L���|�z�Z�Ͼ&��U� �*���Y#��Nn��C��[��&
�T4�����������2��S�|S�Ѷ?�Zb3�C/�5�#�Q���#����t��"��m���B����Z�hE�����ώ��<��y���40���L`����U�H��U��:�p"��&�����n�!.�X�n5���Z��	?�fՇQL�z��6���i�[A�f���و�~�|�t�n���i�߫�t�F��^�t�V1.(¾=B�����b�6�F����8�G9����P����Q{ӄ�&���OKnϠuf�E����$�3~�6dn�D�:4R�_�k
y+�*��|p��*�$Z�Ywꀤ�i[�X 5׏���e��#*����쭢���i���1f��t��Q��	���Q�a\߿�����>;��җ�_��-�r��`+L��-U���[���H�c�ڹ+L����_�D���)G�ׄE�-+�}�������;��0�
�q-c�w�R�~ǦV�G��H�H�)�=3Yn;]�֎%2$%W*;�u�qp������n_6kh�#��]��z���Dv)��b��,J������x6^���==����I�xR�O)g�I���s��H%h��&>s�YDր╜�DƣE�Y��H�����ֆ�1���k�_�P�g_�r����b������$S�黜v�	섎qoG�ڟet�b伶�p�z]�#�9���my��#�_�o��Dł�\��r}��}��p��{�0?��.G���.
�$usS�!��O�q!({�<��_|  ��
��(V� HS��23�,��B0�U�,�r]�j��>��n�}q�n�8��޲����R�S�a4t�{�<mF�%�F8��V(�ǧ8�$�Ƴ�"������m='M��g�g��4]���a�{��%����uh�����L���:��P�ƥ���GR�{� �l�ۈI�-��>��(wGl�����n§:ֻ,�8a"�ss&�H�cJ��5�Ü�DDq���2q|x�T�^��@�����U��
>��FUL�\�'*w���&Y�qW�b.�9&��q!ji"�#)577�dڬ�m��s�p��C҅�R �Y��$�?�a&���'�� r��]�.c�rvPl*�t��P�*��Q��*��J�'9n����HD�Uq�%�@xp�ڋmڥ9��jA�R��"���8������Kd�t�����S��Q�5��e�:����K��ӭ��=&C���1\�#$J"�Geh�,޶��o3\0��ܘ�\��BY�5BA�o��z�|���٦�KQ�h���9i���`Do��	id�d�+�!c�1���%�{�R�~%2�h�]��L��WEO�����@���N�tR��<���� D"|�Z��V�[! C���o��{����i��v��^�C[ �U�g��*ҵV��8{`����
0e8 Hy����p��Ѐ[�ϸ��VY���n�1ȱI���q+S�
Ƌ*	\5��f_�D�p���v�b���?%���a����s����w��|�u╱6^��I^��kud�'�A�Ϸ06���CØ�w���-�����/�T[xـ����zx�!?>�^6�?z6����-��xS�uD�QO�O<u�W�g-ڋ>�A� ��FJ0��5���~6N�gh/�@?Za�?*�BD��鮍�� �;��z*�K��hR���6^�5p�b�$�	!���0�{�Z&
�����C���jۆ7+^<����� ������047��>���of��O�F�d��@�%J+¬�)��|�: ���h�?��P��"Y�B��Qژ�V�b�)ULG7h[B�A�)I���I��� �
e7��o!��|;�4��yח���ZC��)��4�@���� ��c�M������ �ǿ��ZF3Y6�������ub>dH6��Xl����̼�MDS�Х��/7e[�&�/kz��?
��ћ!�����)�8��I���Ƽ��S�Y����E�d���J_��ُ���Y�P��5.����4)�q��z&܉W!a>�K�R����R��[�D '�E��J4)c�� �16Qp��>��$��L���XGʞ��k1;�������)W:�{;��q\�����*f���у*��*ϡ*�SEg�I6�bߒ��N�z<����U��h��Ս7��/4�¬�O��^b�	i!]�y8�3����	�j*Z�r9��$�`)�=̚�|Cz;�.��lz�k'�ۑ�>΋�lT0�7-N#�`{s��Ol�B�c�cAt\�LS$��;�h�e���*�f��=�P�`SN�w<�^oq�*>��[@�S߹䬏.mQ�V����O�	7���!����М3!�B���yM,��"S%o���HL�]��K������f)W��C�|�ᖅ�v<�\ڋ,�2�V����5��Y�i��}~�ړQ�ޜxw��7����bM�|�{Ӱ5����l^&<�$�NAv�8M����O�XUC����lX GA�y��Ƒ-�D-}}��P�:��@%����k$�n
�$#�)�'L�Od
��1K@�Yv���7(���8Q<�U]4��|��ag�Y���/�1�L�8"u�eb��c�����qhvp�C���ΗF���8�E��\�� 4+U�!�����_�4i��)&�!���⪃�Di8��o�G�^ ܴZ[~�ˡ�b�2��mi�Q�O�� ���?�	�.A9�h�^^���.j��M��u�Z��A���5
=�K�s�{���'���c�%W�T����j̓|�i�țy���Ρ��>������=|M��,o��K� �q2�����
�aYg����	R%0q<�m�G�4{I�Ҭ�%LwH���Q��:�+��'�6	|6c��6<�Ė-}K��D��[;�6�-��[jW��&�u��^�e@��乓�Z1��YeT����>��9#7
&���џ��-�tBhH�YP$m���-�%��bG��ㄅa������)s[�Sz����<��P^3�e�띣��.C��+cǦB� 쀕6�}�cl��M.�t�^[�ആH!��ǈ:l�蛜�6VGPP=-�>�ڮ���*�M��R�c�9H_�;����f3R��~'�ɑu�1���^�޸�H~�U�������mX�oj�`қ���1R��o=�J��}䃦o���⺻��Dz�?�>�`�ð��e@�O�����\mH�r$R8�XҩaS�Iu���f�n*{&��ԯ�$qi����Y`2K�#���W
��-t����r2	��J�-�k�ٱ(�
RE1�a"zwH�*Χ�
o�x|��k��'���u�E�j��ɚ���������ԯs��V(��i�E;��1�/ &��>���Y��.��"�<v������z/Z�hI�x�=�x/�8(s7���ҎL�g�#��k�o-ΐl$5W�������,��B����<�(f*�?@��aC=��о	rN_6GB�,��@�Q�����U)]�w���I����Fx%����������ةa��A`��F� �*����b`Ա�O��y%���$�ЫI}�n+c�	*bS
�:ʼ�)�j��f��}�J�[���E��p��R�+�<����=M	�I�|���ƺ��:ᄒ��i�qm0y&�Y��L� �0J�b�HՄ��� ���@� ��k �?h�����E��e�%h��m�s����_/ە5ᑸ�F8�xj��/:�o�E���@��i�g�*�K�Bl�vvGY=���#�������?�A���1�T��6b�dѺ�ұ�rȺ��rܸ�+"r���iQα�Bu�Ф�ߎ�B�Qbm{{���Wo��:(��y���x���VX�F�Ǭ_M��3o���i����h(���I�P��D��4ἠ�
���|�+�te���;G�WCHT��lˉ%�u��}��y�ũb��Q�Z�l��{�U�gpCJ�GW"DN�w��v�o	����)Rʺ(0�� �}���|)X*>&�-������8�c�����4��&3�Uګ�1cGr������؎���챋�_JU�pq7/o�v�e����q��z�~oP�)��q����AY9ֺ���\CfbwD��x�K���B�ܣ/ٍ���2.k ,(�����RM�#�qo�u�Q�'�ºh>[�7�נYe,��@���q�g�Q,�&&Y�7�0_Ke�U�>�2@E����:�p�b��/ݙ�p�8BN��X=�g|}{���d��ſ�Hn�P�e���K��oA&�?�'i�EWgEm�zMrH��/�yN�sω�9yK�>�˃LA�@6iY�$_ݽ�����M{�����օ%j�}�)��f�^��%IN�(����lv����q�ׯX�j�[uF*�m]vq�|�#�;�Wǌ��F>R���(^�9�l>_(hJ��p�}�3 �IC��������|�)����I^|��%��WF�=�t��S��A����5/)S��F 3�������;�ŋTʭۉ�������q����J������lޟ�XJ��Q|'ϭm����ѯp��������lWz:ԇ���VV��O��8��z
������s���)p��PY��K���8��#[��2=��p����@?�t��y�]��s��B&��Ӓ���d����RW��.
��fne6Z:z��Ѩ����M� ֺ�~��~/E6��I鰫��r'�M�6-���#�2��v���`A�v{�0o1����n���I�c�w���t �c�Z�O1�l=.��.�e��a���� �yS�_�􅿌vɲ�a��8�n��K����,�>�i�l@1��[j�Z��਩�i�mQ��	�R8j�ZY��'`�m�El2�r�$2o)��9)5��P(U�vr8��J9Ɓ�d���Hd,��P/Q�hX�Xa%�T�)�|iNJ{�bc��U2�� \4��}ǈM/�06�u&:=B��5���1Uv�nR��!�����BN$a�v���*�9�ݧ�⹲���,��NW�o��Ѧ9��VA���	�EN���tKa��� X���F��*·v�{_����!�����(
UI�5w3WY��"�J�M�{��%-� ���p�j�	Я�y}��0�{�Xɯ��&V}����\�b�d����y�غě*VN� �
I�vj�23��Q��F!Dd����Κ	u�0��y��-�q�g�(
cs�'�~.R
�Nv��:�q�8�a�U(/M���d�'צ7��˪��SQ�ҕ~��.!����`%i�����W��$lE��:�?��"�5ן�,�Pզ3�!&?7�k����-�\iT!84ohX��6�qwMx���gH�,�I�)N��uEF�ITW���Ri�[/K�i#Y�����8YS�BqD�{�]n����MI�ħ�l�x��<�	�B�8����ΉQt�ų��ql��HƸ=U���r�	����/�8-]��)뗫����9��#b�����rDq[L�$$�� �}ȝq�{O}E�I�h΄�ճcp˴mD�r�\/�>�B�� �^���by�Q4����kŭ�9�8�$[��V=ɻ@���}4�-��O��Z/�_�G��.��6��������Wn5��O�<�m�>�4�}=DԾ�������5�Ƃ�2j��c���_$�Q�p�@NU��W����)��`�L� 
v�R<C�@cM�t�T��F�JǵP�p��)�L(6E�-J�e8�E��N�T�a���5yj';%�&Ծ:�~��j�a��w]PR; �>��4띾b���p�"Ѳ��U�o���V�I���R;�.��h��6����P�������&z�� m�+1��ĘoW�#�ƙP(��Ѡ>�4�mG�P��w3���s�
(��uN�n���p$Њ葙�n޴����u<z�\l)�硃�鹓�j7N�c��N�WT�GZ�"��*�=�A���T�ߕ]�Y�G�G�nj�S\C�2�5Dr�* E�_+�|�AD��E���5s�"��A	X2N�644����iۣ�,�ȱ����\&��O6Qw^1���q'J!n��^[��HM�QחF�K�Gp�۩&���u��h��"�pd�]@���z*�Z���0l�1L�Ú�b���ӼXL��z��hb*W���.�I�c�����R���;nzk�Y�	W�ǧ_�ɝ�$��G��
Rj`��k��F@W5g�4RD���o�p�q|�����a�V.^:��-��aQˎ!�܍���w����e`Â,�'? J^j^6�.^]�PP�3��QN~�6�nk+��6&���-��S]���e�$������7�i�<��S�]͗�����wq�:\(�ޮ��}�y��~I�
�91���h3�@ ���BΉ3kG@+�&�黓ȏ>W�<��4�#�)7��'U�jgb�Dz�`tUc��?d�%(�l~STF�t���6��_�����=��B�N�>��C�U{�YU�M�,�z5(����:}���F�0����r�D����� ��hU�^S*Ÿ�3�o�pSY��@7�ĵ�����뫴xb	����'����}a*`���
�dWm�/���(]���P���Y��vfx���N����μ&}s��I�=�U<ET�	�  �b�_��n�=ƴ��3kEc��}_,�lh�@��"��)�c��l�>���Mk��#U��v���/�E,D�����ۀ��L�T� �c���ފ�ڣ���B�mG�ø�*Z��Y`;�1ODv�%�Ǖ9QA!�f�,*w\\���3+��N�+��^��H�����X��#u���^*��~��R�*+��c�K[� �e����{�`x~C��������|9D�uRg���B�`��u\u��ѓ�Rg��v�B�@�;N&tq�Fj�ɘU3+���"�T��r�p?2#U�4�<�a��NokZ�g@ݫ�EN!JS/���Sh��Y�����?J���LxA}l�D<y7N����ҩ�UZuW)5����XB*�;��3��ϐD�!�V��4]J��0 ��'4Oe������Ms���[�/�Q�h�&�-��C�$.��&%�^
;H�s��|� ��`@��z7M9lN�됀�-K���Xt�RѶy1b�Uo�E�`l���ё6F�u�;)����a7D�p�f�A>A�pNr9���ѕ塬��I�8�ڝ15��d{38��,3�Y9;�>�bϵF��ANЪ��N�Ai�.f8u.�L��.h!�x�-w"pj�	E�O�a�C���K���������]����4����� <�c�V�E>?�zf���z��+��8� [S���,ﵸ'jR��a�����ad3M �"�`��_��VV�ޔk<��֯�ه�FoQU풖$S��T��18؆�35��"fg� P���L���I��)�-��W�������ӏ8v��KL �d�.�\D0���0�8���Ck�]P�e�"���0���с�/��	VWkQ������V_����M�\ͽ�ea�$i��Z�ԃ�Y�g̶�{M;�k�^f�e���~��&�B�
���xG��@�� )���8c��g,n��W6ޚ�����RJ����[�f2y�TŐ�T��x�EЎ���̀�|�]���?L�<�B�exu>T�����~�͆����;�j�0vǄ�)�F���-).O�4���7qՌ�iz��"��g�n�g�neEy��=���_�j�V����6zu�J�*Bf�A6(��R����'���=��{+���my��(2��RU�ҙ���=h� ^����+�.v(I����o�R���H
�v�.�{.c	���31Ďɵ�n?3�Y&T���1A�%]��lR��4�B�sm�w����z�c�m�9#�v�}L$�ͩ��M����͉h7d�$O�Ղ�)���N���w�d�3��b��>��v�ą��r1ȗ|%�Y�P�̨V̈́(�yvyG����c�o_R����f����e�>�eUY�y����2�N����#��\���{LGR�e�� �����V!��2���",���t����#�K��t�:We�l��<��
��~Un�l�	lZu5>�CWH�Wb��l;e�ք�n�ئ�a-kjR�k�FO��G�D��BW?ͻu,l�&��Z�!�?��6��-� �lZH�����󁯦q4ʭ4	�j_��������z����/H�u�ɽd��
��6��k�4j��������շ�$�n�gK�}�E� B]IZ�n�C��T�p�)��<��J����Z���q��(u�9I|n [J�~:|g��"C��W,	<Q�R�C����za�m"c[[��.��P]��q�) v'5,��|JVC�n�bG�j�]%O��-��+r�f�\4�}O�</}H�H�E�hµI)6X����)�.�'؞�vSRY���L5:y��9��z�?�i��������y#��e��:ge�p��ᦚ-��P?����$������)�6�d��7?0�c�|���S�mj��ʔ��&{v�J�H��!
a��nI����Ñ���_�g�c
V�v����2�Ud����i>�IB���&��n�T�~�T3��6�x\�7a��X�� �v�@�k����Tl�N',��fx�1T'꧓���5 l0�)�t����G�~!߲uŤ�6��	����k��1Ж�R�]3�� ��}�����߅��ę�X�㨀R���,�@q�9��0��U�����ϱ���HB����ՠ�0 O��5j��2R^�h��3�?��^43(F˾@��039���
y��b���=ˈ(
��a�bĘ8���e���1��g������<�H��v�7-d�?�
f�����B����l�+�w�rw�HeY}�<��/7�h*H씕���%R0�?)�	S>Oi�5���-L���a2yEEԥʗ�����H8�V��c��vd`&b.������[l]D��|h�M$�B��^Ij�Tf��P4x�r����C��B�I[�A��;!��.����v��-,�S�s�̣� �	Ns��T�o"䎐l�����<�s[w���G/�?�������� ��6bӱ�R`����	��!j �@a��� ��ʽ���uo��X���jp�d']َ����!�n��������]���ʊNq!k=2
�[�Q�x<�������H9�tYkWW�����g@����nS`` uŠK�ʃ�*
t����c��
k���t��~eU6��_��h�#�2�nH�`9�S�����O���:�ǚ?D����ݯg�_��rH��$@o�n&Ô���-���)|��q��9�um�l�6�8;H��>�eF�����x" ƨK���q�1�\E�C�):���X���B�n]���וc�?[��ɫg.ӈ��e�יI���8H�;�k�0�yr������p&T����`v�D��qx�����됢�U��av4�IE ������i����1ئ�c4)ƒ��:$�VC�T��h�W�
ɧ`��'k��PSB�'n)�!s+vr�?fɱ�����9�YϚۂ�<i7�d����K��G���f���3,Q��|����_�>`��=Lb���J/�k�!w�$��`b�Qz������T-�����BR��(Ɩ����9��1�DD��^��YC�j���-��u�m�[��)��;�c0GJk'����0���#<���Q��|P�-@Ƃf���\�٧-��gL�O�49�C����8��cws�`��}Jhe�a0̣p�B�	Z�
�Hv9�W^v��6�ܒ͏�T���69v�����b	�����GQ\A�SX_��rd|��`\y���D�L̝$9���A5��==U��}>L�L�@	4AwLGv:"��(uY)�׫�������Yq���z�X^�Z��98�k{y�R��@!]dm��B*�=�����Ҫi���Ђ�-d���v������ԥ�N�c%ذ�N�ǒVU��I�M��T3��NW�:���R���9p��.����p� ��~��%<��<C�Z��Gҧ|���ZV�O�P<i����*�^d/쒷Ps���`̼�d��.[�Oѱ��V�p�����iе�֮��t8��(���!����$X��jE�oa�q��lH���fi]�4-���V�d�N�)u�vH��f��UZH�z(� �j��<������U��!Wf�N�J�x&��-c�h�n=R���%͐ؗ��6)w4���I\u02})��)!�u��dʩ,ֺؓ=�bͺ�o��.g��eNc��#����$E e�*�X�#��! �[���@~�_�a��RZ�8������g�n(��j�s�^mY�3Kj�=U�j���Фcۿ2���r�Q�ēGp.I}=O�J9μ�Zx-�򯯈DBB��"7�q�軓�C�I$e
�=0'4=����Xg/��2��r
�+sl�#��{�s��1�y�| 9�n�(�Ae��W3K��S��>1;�n�<����۪J�[Hǧ��(�T2= �31���<���,�"R�)�3�C�ɇM�k��IBcpΟ�慍R�K<� |�Qf��Ğ�oM��aoe!ÞK4���`���y��e������g������!�vq�K��~�Ϸ����/o�^N'���
B� �dc
�0k�������}�˥:rkم U6c���r�͞���m�`T��.Uv�X���QH}�`Gb�1��q�{,{v��1]�(��k����9e�n�>x�m�=���eivX�EO�Rz�^��y��?���pT�*��n�CG���$O�ߚ���`PL���/,깒�i�~i�	\��)�Rȣ%:�w @$0����Z�~fN�Se�gQ!�f��#L�@�! ����ķI].l�L	�+���-��I���e-�d�O=s�N�����P�>J5Ä1D�����)T����$]^�D��2�f��z�	�c�������� g��,h~4��+���7#p�bq��D'8Z�)S��{�~��^�l�޴��)�-�]����@�.s�jɣL���Č	-����ﱀ� jZb�$s�O:�E�쌘+��-���m�B/h~~RB޼��a���@9����'~�j�UW,2�˙��)��i��E�2��%*Hv�\���:(��W����V��U中�3��ɍ1^�S�0�fn�Rc�#���E�;�y�fڷ?f�3gA�d>��Ç?�;�2�a��S3_�NXq;x�s�(�I����~hT���y��a��̓�-��D|��x�S@��2��,w��i��덁t؈�у���-kr��ZR��>0Hi}=�(������i���zI�Mkq���ɭD����ƀ��Ķ�@�xz�t��A*���1�Z�ڹPi�/��kP���R@����r�K�)�^d�b�8뾯zl�����+`w5�� E�����h�p��B�d�^|M}m�z�F����G�+�'p��b�"�Q������Q]J;�n�,��� k�x5�x�s��K3�(�u�.�fa�iC+�����Vy5��M=�2g�)͛�I���Ic��Y)�����dDܦՀ1nd��u��ۓ]6��O�L��B�p������	D���_���d���ڗ7����� �k�';B��$��%�<i�J�*,�8��l�� ��B;A�u�헇�x�C9~�o���x�1�/���+\Z^#�����w�s���"ęڄ-����x�Ґ�d��=�ׯ#=��`B-G���H�u��i��'2��q����?\)p���v�9�l	�a󓯕�pqz$�?�`�9h�$lpA���H6��\��3�e�:�������t�*��he�er�g���<���pج
(�cn��eZ@(c65�hSF>+�q��P����aF]�ߑ	�F��{mK�؋C�����k�I�UMq�Nf��8a�É�D�����A��V(���^��6��{2�tR���[�^g�z�?w��
V%}�t����g�3G����62�X(��I����+�n`Ry�ƅL�AR��<K�){m�M��҅�ĝ�	���h��a��(�@^�؆�3c8�_'mf�?����>��������g�{�īP�l��v��o�q�[U:�k�������U���ý�[Z��8n�0R��?����$��k����wWd5�q�e�FVH6�3�ڇܡ��߼�0���uޫ+0������j^\ח:����g�����$,��q��1ڻ6W�9F���m'֓c���ܥZ!� h�(A �<�S5�`Z9����mBa�DW�2S�$�O*&���ꏹr+f��-.}Rb״�����g�� {m�3�%�wm�V d:4dz���f��x�V��7�w��{T�A�q��"w>�O0/>y�sd�}�e�-�!�#hsh�T�쁜5�M5�������p�M�H��A-��Twp�&5�EZIL�FZ�l��̀i�yᠾE3y�U��a?t4���J���l��e�gԾ?��}��=���c��!2FTBf� gS�#ἢ:��4p��\�	�o|-��93�Ob<aQ��<�[6�����;d]l�]֕�yX�q��t-zd��"U��&�0UM���V6�	\� �F�@&fN�@�o#H�c�J!��1=�WU9� �'��U[Rذɐ�I�}���^2�ܺ�7d?����l��O�-m!I�=�b۰@�oǦ#�X���q�����7��<~=w��Kh�-N"�s+�R���@B|ߗ%GPc_t����v�YbM7r9TF�hy�f!ϸ9��i<��[W�ԡ���� qg?�����[���&S�|3�4�i���<�@*s)��\~���\���Ҭ�&|Z��R�4�$���(�X,����'�vs��.�H����w��G�I����/7����9�N�X�v���c�ẓ%�������6��>�V�
��'����!�9Й*�0��I�ܳf��G�x1	�=[���٦9��0��{_�n	��,G�X��)0���]O6�ݫI������T�y���Hl;��އ���W���IdJ'�E��WJ�e���)}�li|+xsh��cC>����'�ʐ��f����9�ݭ���R~�*G�$�"��{�i'���,h���vb�-���e���U5P�vD��=Gs ��"k��~6��xf1�ܷ���)����9I������n�+w�_�	Ѫ�an��j����VA��e�� H����_�����|Q*�gh����>�ͼ�7i�ް���`�.�\^�0����t�:�����Ҏ+\������S<q���0B��ȸ[M䒵��M|��=�~���L�A�B�7C%�3�N��[�sX�vup[���+��8��M7ɰr��l�B�F��r��2}��lE��j��{;�������/��```�D�~7�0q�}�v)J�KV O���QB��w��;�÷�~���;"�qP�~c�u�ɦ�?����A�rG�r�*�i=5�M����P=��t��ֶc���t�A4f�m��-��+��V���E�6AJ�ߢ$��>������2.o/��F�b�H�"H�.�M��.	��nfx�3Ek��v�����l���	�h!�t��JbӒ�Ŏ1�.������r��}ܐ�֭� �.��EO��U���W��Աqb�y���0�����Wfi�1��^8Ș���rی��sK�"���`U(f����ټ\�4R�c�ԙ��cnX7�ma�Pq�2����΀v���WÞi��Eh;L%%j�ۼ�z$e�.�#ׂ}*�G^�:&9��&�-~���M,;�m�2FRK�ql��c��ՁC�2�;q(��8'�]�ϙ)�z\&�A�����*�7o�i�O4ѭB�N挆���BD�S�ڭ�N��$#��(�?��M�]0�*�&�h�K+���QsF�^�lQ2�1��H$�x����Ip5F��F�T�"�����#-�����q7O�=\r��x�i�l]�	���粮7 >�1k<_<�1<�������� jU��9�.���K4<_�NB��]ʾ�jV�>���+\�J��\0Ռ���,0pa~�<H˥83S�}�X^�@��l:~�q�����w�%�k<̶����M��ōQ�����F�!#�ģ�2x�̏)I��<f�j�P�U2���>�iTt�J�c@,GS���?��ͧ����P��V��ݑt	�Q�<6�_�i���,���c=��x|$����s<�W�dB �q�+�u�ہz�nF�>�c�Re�� ΏL')��S%���"��&G�F�֌[i_�W��=��$K�&Dգ������T��=�&��hS��V�xI�i�6}�@�����"��5#�J����-���������66�G�_��(�t��c��n�	��ŏ���ƾr]o�{�T�C��d�7�]:�6�X������w�[�� 12ǀw�ovn��y4�k��<;+j�V�N�U>@��cY��D��3z
dq5S'���c�@�B:�'��@PR>qf�W�-De]A�੭��KǛU�����ߠ����t1z6!��JP����o}8��b!12@1}���A��CΛ٫F�э�2ah-�)��r l]��%��$�)9v�oao�p0:J�F�Ecƞ��)�Z,�V��6�B���a����Z������R3C�I�b1�Fӏ�-E$�f�����2d����¸.��񦑹k]� (�8<��3�ǞU���?3�:�������6��g�yp��R���W�h:����*1,zv���*���js�v	L@����V�p��|;�r��vMڌ�# bk�hQ{@XSuc rmՖ@�y=;M���IZ���Z:0ʯ�i.&2h��Dp
(��X�ujShv� ��#�W�vޕ��
��gT
�'B����8�?��ӈ�z9m���#�{5G�G���gdyH��c1��?��łػ@3/^j1�rQq��i����I�	+�X�q��������F�U��&]�.;'��&���Qj=�C����S���Ͱ7�G�u�U\L�KW	��J�P�8�}���U�9^g0���_��K}Y�o�>ڦ��j� c^��I�&��������ꢚ^�ws���f�5S%V��	j!}Z�u}R�܁�k'a���^�IJ:`(�o�P���'�nf��x��,*��U�KW+�d��r�<��-�����!Ģ��M����'��	Ċ&�I��	���h������:'	Mq�-~�;�R�[���l��%4��~
�������غiL��.�U�kTFӿ�:�e�ɠ�E��ǫk�L��O�`ƅ-�p��B�I�^�W<n�'�(#<�j9=��m�����(�a!Lv�UF��
qviP�47��0��ߔ'�z��X���\`����I�s��1�k��/�>x��Ӻ���he6-A?p��gm�h +]�T�x��`��5/�͡�G�/�Ss��W��;�ͺ8`�
WS���q|�^h╈�\�L�����_tQid�s�Y��_�;ٕ��@�K�77���@^a4�Iv�g��_�v�ł�?�+�_�������]V����;�d�b��z��)���./�`yd\�ڑ���b��Մ�Q|e�]�;v3Gv�%8�r��ٳ5~z�����kZ�;�僿/П��y'c�ʟ#�w�!�B���^��ګ�	��Cn�9w�%��k�2Ёp�p�mƳzp����&�9j�2N�d���o��8�d�l�z�
���)E�:�p��z�����zy��by�b%��{L�Ctv��0�<��,�^������|��
�o^�˔A�LX�y�nϚ便��,�2����F%��]��F�9U}��R�e�e^6��a���˓�����Y�V�ɱ1�Jv������1��aar�ĕ g#�C����heA��D(�>��|k�	�R�&љ���{;��̋�6��V:6/ƪP�r1��Z�$�qҸ#�W�5����G!i�ąuD�T������-��\�3����l�	��^h�Y�ѵ�s^9s���'Cg2�
�ɨHn61)�z|a*���`����/�$i�C8�R=����`y�zx���n��Xl�Fro�L�^6"�d�%���<��r(J>�9��B�[Kf���(�6Ҡʒ�~��&��v�F���>��c�S��'�Ϙ�qb��:v�@�_�o1@�m]���1/^�|Ƹ,1Q1V���Jn�Řh�s��V"���B��v(��VD�jQ�oL'�a0;���2�K2K����E�tL"�
�E}.�.�����-�>����TU����Y��y��0:h�O�4y`��ڼ�u��!��p�������=���{�.�8���RL`"X���3'/Β�V�4�����]���!�z��8QCw3���C1NM����1�'�m`����h(��P�=P�n�BKo[����Nƞ���
S%I�E��Ψ�*>L,�x�����?��X�Й�����8.�P/X�]�gv!tR"���&�%\)�e�	�Z� !*�$��	[��)h(�t��������fWA\k�B]]6dP��:ec���W0/�Yr���A,���g.<�7[�����j!�P���4��k����CLP7|�`�N �&:m��TH�-b���ā�e�5���iH݅���<'��f9��
,���HݛMZ0�8��'4̔���m3�.�:��*��^��8�nqqqu9e G1�ڢ����vR<+�'�PE8m��M��\j�5��Qπ���j�3��ZB/5��6��D��j[�~Y�aҘIT9���6h���s�g����x��B�mwl����� ����EK۰ރ3g�
[����I`ӝ����,IR�f�GR󸯘�6�0�.(ۍ���m)��#��g��򯩍�-�yC�/=F�%�� ���'�ѯ���6.+�C�8�qzZ��HLBS�@j�5�F���2���J_<^qN��?�[T&O�֡ZV�V��>��i����Ye��^�P�Th@eY<���p#,H���7�#��0���I�����~���-�r�� }�'�K�W�߻�������IM��=�wo^�@��
�J��/;(`闃�=F��5�h����P*���>��Y?r�g����dɪK�� oED�OQ�ME��̽iԇ�I�<�df N�Kng�yQ�1���`!��%U��лO/r��?��.Y�S��J��odJ����%��%e�T@9�	�Jc`Q�¬��@�53�Օ�<���ئ�\�g��� hv(!AE�ֱwu�X�O�����py�f-'�/����a�_=�:h�֝2��xʐ�."
X�� A�7�^����[yh�12 ���V���yD+�c����V����ׄ���e|;��ZV��7��E������~s������ڪ��v���_@O����F�0L����a�OKG��)�j�}c^#1�0����A9J��8GR��l]�D*��ok*��+/h[4�!YzH>#'�>}d4��$&�d�}
)��N2��uo�|X�<X���*��b�[��U޴ᑂO�4χ`�HH�)����9�]�O�r�?j
��]RŹ��	�lؽ8��5��Pr��G-b8�:s�������?d؄���j�����j?�<=]��43�^x����N�E���^4���q�h,�E>D�t�h�Z/O!��<tPs���+~(�$��Z)Xؚz� ֱ�%��_s{=}��2��R�ps�D5�2��k��Cx��.=�(ޝ$L��P7J	T⸑d���:��<����I4���1�#�\n|�(~��i��5���7nP�N\K�7��o��Sm�]�5a�g3��?H��{�[����5Ɋ�;|qD� :`��D(�Q�lb���>��+��W��-:tm�G7����U�]t�e��Z�7� �;�BFGm��5����EJ��T
�L���dx��@��D�_Q~�VCu�̏v�����'(4�Q9 6x�f-�T��M/��Xhn��!Vߧ�ua.}q*��~̀@�饑���)���M�<�~�����:��cr��iM>'Ck�tWV�,_E}p�O	���.My��p�-6ŕ.�,y ȷ�%�C�3)���i,�}cL���X�K�����|�$�M�
tJ�	�'�e�F���]�f�+�⌙����5F�qR8��dZڸt��4��D%dه���� U3F0���,Q؍�R���Vk����h����)v^��ǯk�d��A��X-�Ғ��H� k�%��M����`���镦�RDT ����A*��gPBU��"�~�f5����<���O��2�ԩ�ۈl����f�󚈉���/�$m�H�{o��������A~lB����|w����y����d�h[�*4���EV��_�G�dd�n�`	.��c�G�`��HG<��~���PS�$aZ�9��-��+�)B��K��]�7+����'e�v�7]����������d�/D��ml�-�e�<�q�]U�opY��A*�V.��!�Q���h�t�cAW����_nL�|E���F5v���N>�F��.ω�r�
���r�9Zʮȯ�ľh1�ܲ�/�����=�����-�p�IO�^T�i) ���� z��ܦ|�E��YEn����s�X]��`�k_�� ��9%��Il�`ieQ;�_�H./��P& �%�:]��>w\\Q�Ju�U܇�w�B���8��7�vl7I��W0�Of��lʠ`2��fY{a���b��<6������P�ݱR�;�&D^�9 B���'�=�C�q5����;�N�t�T\<\:
�5@�}9>nj�[�[�!� 'Iĥ$~����N���:Q^wc�L���c/e�Df����OۧT��1��Q:����'z�f����c���2�w���^p�*\Mi૬4����N� ���0�	��t�R��7A��te�� �5��u�qyM	{C
�ߊz"s`3D9����za�p{8�{��'���� ���U���+74�YN�ҏ�g���+�v�Ł����íy�
f!���ј,�ti�:�|�ë;����d�m�x�Y�(�]..r
��~m���b�z�D?���֯*(�:�D�\�a��/̶\oءh\xC955߶0�(�����B���@w�Q��#��ts$W��]r3T��R����	@4��Lpl���v�"��PގM(�d'b�Ϸ������ji(���h��3>��Ot5�#�vn����V@9����7���	�4JoJ�Ln�����竧~�Р0�'쪌wSh~�F�fz����g����n����m&���� ���P�IY�g�~["�L�B�Ȟ{�?���b4c��%1��{�o��O����&�RG�}�o�u�Nm��̤�1:3� ��,D�CWa�>y2�Y6:!���Q��"��3��_��}L�kHH��մm�}�q�|j�$}�S�Ot�?__Fd���q��d�N����K-�E�3I~$�d��+CtEw<~�#�{5����T7&�Է:�"��G��۹l??j���~�d�l4�v�
>?���'�OPN����q.�z���\��ZS0ׂg�ܠZfv�3��S7mV��.����%��1G��00{?�ט��4���:=��5�������j-�����j?�r���z�+C2��̽`ܙDp�ޢLt%����v?��B�y���z�<0XY�,����b����hz9m+�n�jTD�����s���B�F��'C�zs��k�㈇P0y�q�l������r��-�l��M���{�悯��y7����8m��Vw�|�l]�8kĉiڦ�J���<`-�.���p�Y{�=M�q�K8z~�'��>���}:&��/��cH�6EQ
Or!�T���"��PPoK��X9QR�>��Y*��,5o6y	���HKͱ�݇b.n<_�y1���`�s����:gc)�9����$��fh�o=��H�N*d���2��u /3�[l� n���y+�@?X���ҷަ�q��-\r�݄m~�%뀰w�ȩ�V��5і��mO��ظ���iw�Ͻ=�{Y�a?8cX{��%��Õ�*ٳmh��6����b�����'P�i����ve�Ot+��pD���ۖ
�R��}tb�S��W�S*POF�F����(K �����]�&S~y�=n���G<���ü7�0M
��ɳ;C$�:�]Ḷa,u�*��i��[	&�Cd�%Ս���)m��r�b�[�[���CDW���nM"��(:yK�ʡQ+� ~��k�m��|�v,k���^���CwAvB���o��L��w�����*=�BHͭ��m����x��wh�Y�pX�4�؎Vo���n�5Z�W�t�H]d�i :�<�GR�H����t[�
*g�+*�շ�yS?]~͋u��VE��j�9W���g���B��[9�W2��<���ێ������qtF۽��HDE�<�үs��8�����	 V����[Ki�/K���M��z�ҐbY�S�z��=�2�,ƅ�C��u�������Ȑ윫�6�U�`|���aLbs��~a��ٽ!?|�
�C�:�m�i�&�v��HeK���!4sBHG��qr}A�/�y���z�Q����P��^j�BA;
ti��i�D�3���������/����.u�9Vdf4�ʂ��i	�����	[(�}4���>_��aE�KJ��娀z5�n.Q�THP���h]R��q;U�*����;��L����������<���{[��W�M���D7�F8��.3��+}���> �s��8�����Y�?�T��W�p�mOt$Sk_�Řί=��r�H��t@j��eEWG���9c���Sy�� �N0��y�_ŕ�>�]������5���Q2��Z̔m0�6^K�G��1w�ۃVf>$�iz>�K�;1�U@�:�İqC�P��9t��HΩ�Y����N����j2�,!$Jg�6�-w�`X5�( �E+�W�R����`��2K"�l~9i)yEf x-/�d-�2��w��������G���1+�T#z�Ӫa��x���K�P'B�x�!Й>z�C��	
y7���l� ����T�C�}�%���~�>�M��cjF�\�u�����gq������}�*U@?����6�D-�g�j��6�es|[��eP�ʒ�
�̮�����y��ztB��=�	s�����Q>��'[2q0 T�����f)os9���HJ-��j;N���^`|���e;�PfJ⎗(&m自:�I n�d1خ��J~�_�;�>T��>kjc~~ʹ�c��^�[{�4��#������o.������x���`b��dUׅ|�����`�8VdsWWK��/~�f��)�D�@�����"	t7��9��/jS�W�0��@�	8W|�U;�4WIh�1��"CMj�4�D��^GsVe�����8�0�����E{� ��p���ir�(3�P�K�4x�����{',cE���}��P��6p��y	[�V��\��:ځq�2毊b��kƝ���J��`��b]^�oG������{]�`�Nl����L��F��9�f�݆�iYn�Մ������U���	Dl�J��3_�V��[�[��0�	�r�le�CV�I	�:��;��xi �5 � )��Q�FME�c��ĤB��rW�i������s�O���+D��hH�����M��?'�ru��"xe�	�$����#1spP�B��	�[%�Uc�ڤ��{�%܍4/�C��:�ͬ��hr:�-g��XyUЯp�� .�
Ҕ���v��r��cx�����V�~�_�x#А5iG��c��e^��j�!2�8�A��b>@��G��薋y߇zD��4!N2(�s�7{���yL��H��|fW�D�7Ԅˬ�-d�U�y��7<� Sy�"�D�k�!MQ���e7��76~��5ُnFo��Cd�����a _��{�gu�Ox�I��7\��kq���u:����-�(�ޒ���������F�8{/�o�)��>�ۏ<���S����{\���-[�r�%�4�n�/hL�1�k��`ive���8�D�r��zK�0��e��d��a��	@b�>ҿ�}����\���z.t�x`4��_$K�Xj����.%
������'=fɱ1g��1�u ~�c�~@O��d�x��Ӏ��YAܖ��>L�-��
Gb���]q2Rb.�dHBS�2�M`�T�C���<��5B�R��*l*&"�#����wd��KnHƙS��t�g8z&p�=˹��h�=���h�qZR<�������F)k��sr�D�Vưz�+����[�����[���k�=�qk��V���s�7����[3�-c{0<mr1�l��r����Mlם��>@��$�çR�����I������O���K���������d#*�<��Q�;�=��|��5�D����j��� �쳏��:thg!��f��lW8��a�*;��w�O��;�����R3%R�ŰǄI��U�G�ѻ�㽱�׎ѺN|�ܖ)NY�XP�Lg�9Lw(�9�_�>����!%�-�&�]�(+3���r8���L+C����/�8�����@� �\�2����pD��.�\��5^8����]�ᚳrԈ�Vj�+N�6�#�y����s|�u^�������ВS�ߖF�df�:�Kmd�J}��yM�Z+z����7�Ks��Yv�5�-)���[����}>ݷ2�b�_N%>�S����Ű���$�Nq|��K���<K� �CX*ڄe;�S_�|5���O!C��p|��N�*�2x�|�=`�l����)��.��s�w����k$�r��xI�?�i�Û8r��0���g��Z�����]h_��k����7.���,��LP�њ�s�o�� z,�͊q5:p;Q�J6��X�B3�o�tS��(ahY���g�)]�@!��<P��䄔8c�c������� �Dj>f�2���M���
^ �'?0W�Blk"��&h޼i���	��Hl2ngY9^�P�B�Ј��c�?;�Q�'����:�FR�א�M>������}�;vF�)����t�8%��ړ�Ք��-��n����lmD�	���X+ʻ�W���2b�7%�]Ѽ����c�x�f��\���8�:ɲ,N�,ᑴ�j��������"���ݑi�����kOe�A�2����U$?�*8WX������n%]�4od�[*�nA�O�|��6 ���Z�"͒=4Y�J�>e�Ÿ���h���7]hz�HN}(w�r��D}?��w��p&ob=9��s,�ǤG���J���P|�v�`���9U'R#���w�.�[���L�B����Ik�˙<��W�8���dAe~~Ö,�~�������#�+-��n�x�?"N\���p�>N�=�l��Sk�M�p��N溉�^&�nc���#:S�O��V�b�rQ���؞��4�a$��5��"������jf��)��;�k88�O�Ŗ��X��~v��x��$N��J'![&�`�w�jT��_����f.�ߗ���-�!����-R��..��)e\m�\F�͞��]iR���_�� |�DO`=AY�g?\KC�$�6���,z��O�/W/M0�ۗ7�Ѽ�ھZ�l\QO�T��a�10�6̻��n=�'�#��Y���c�D|c\� ^���FN�.��A�l���M����� L����K�CZ�l���$7���8��5���C4�8[�&o�v_dXo6��Ad-c��@�e��=4�P���K�*㿍���`��1�L�ja����m�?�C��(�:UP��y�̴��b�v���K�Mnu��gVs�}��Q��i<4�ۅ��\>�J�rr&̶��|���ķx�K�<K�?��'���ZʌU:�:��6aa��H�@^.f�X3�p����,��ȮX4T����u~�D�z���Ch��6,=jĖ����{�\B��C�e�������I�R"��=1NuT�}�K��ުYb�_�|{�,c3$%(��q`<C�R��6�h�;����gdW��`�NL�Q�������#��$�y���{SVG
|R��_�0?�XK�F'd�aKR�֋PIґM�t��
��=8٧�O�;;Zݣ�41�	����P�x�0���ʁ��X�����J�j��q@ �#�ē�φ�Y�����6������؊N1�Z�B�W���\�,�Gx�m�g�g��|M�+@L�Y��F�����:1�:³c�����|��([�6����ux=�^��39!�*�2��-|ɛ$�����+1��rP�A$�M�.���T7�_?���ӫ�����]&-I�w�o1�W|Q'j ���e�h��<�O�Cd���r�<&f����r�7�(����镝=�*<{��׷����l�l��P��gB������3��"�*)21;wxakG�t�����-y)U�T���C�l<���)ZT>W^X!�0Y����F�x��O ��]���(����$r�F%/�rO�l�y[<|�N������Y/j���U(�uB'5���!:�?A�p����ʯ����Q/Y+=�|��k<�%߼yc@�X�-���{i۬�U��' ��Ӷ��2 �`��-�#��� �V���3(,��o�����{'3�7vѧ�#��� D@$|B���-�0l/7�U�7,�U'}��ng��VO�����������h��Po<N�7�l�����k�U�a�+Q��7�����o �Q9��r�h������O�7;�r����m7�^��#I�47�*�����!)��w��/������t��/a�܏�����gOs�[�v�`�8���h�"km�к2�`�<o��v�3�S��@Z's��@F��P=馧"�[q3�-PB.#�i�>�0����/��@u�ٲ�a�9Ԥt��&B5(�Z[���k}y��Q-� �K��jSv����栃C�4<�y7Ƴ��̖�ı|�N�y���Zq����q>gIy�jxr���Ţ-�.BHI@�v����53k0��|!~5 �kN�뚻����t�H'X��k��z���/����Uo0�Y�D��@c!�ն������=M��eW�r�I��8amJ�b0�����9$Ɔ�'[.�*�����Q��_�H��G-�Y����u_|��B��W	f����l�.d.��0�[�ج7��e�q�D6<3Ԑ�a>��c� �lT�0�r�]�Sz�pi�P��=F�`������U��4�XlH��o�j"�#�"K�+���G�M��3����3e�=H@��fG��۟�A����|~��ѱ���0pc�aO
�6н��(����/+}�2aGK��gM���fS��$�R�n��5[Q3*U�I!��0������$��|���7���=KxdKwu���}��}��\�+-�h�AY��{����4o���L����'�+�6~cJ+e)O�`��Ec�d�@4m��kh��K���X�T�B=g��}�^���H�lB�;�͆i����,�9z�w��Oy�g6���|�)(�Zz��Xv� �ۋe��+��'�(�d�)y�1�?��wЯ�l��2 ˓2y��� &i�Qr�߲�3��gPe(H��V�?�KQ�S�G��+Zk��.��35�Ma�1$:�Ȁ�=�Y@�T���@�y�v�3�g�w�r3���4z�&�Z�y��,a>�O���
��G����`Ȗ�u��Y���~���<*A���v�zhÎN��%k�YJ�P�J�{/�n���ɽL��EQP�b~�u^W�*.d��q���_�(8Rv���,���d�d|����ϭ Ǌ1�P��@�M��j��EA��#�I~���Q�v�Ĳ���)O[l�7i'��h�J���5YO.dJ���:qӛ;����Zt�Aw)�}��帲�&����`"_����!ۡ�A#���T���C�dN�+���c%�a(��ݴ�X�M)��^� `G���]'Hp�a����T��)�*Q�\��-���a���XfA<2�y���zP3p�X�����Lү�)�^Z�>��dμ+����t�=��q�pP�f��>�t�a�����nM����쥮8�cШ���Ya"1"��䐔�� �][	L4b-=`��[K|���s6��G��>����x��#	S~��L�y�7�_�}��6.�F���u�4u��;��M�h$�Ć7�9������2�d[�?��e��$Y�C'����P��؆n�<�K:#�I��W�Q��:ch_�B�A�lk�!��ni�bukm��@H~����Ӗ�K����ȼL>o�h����6E&�V���U���w~�?Һ.�\�,]1n�J�����dc��B������,��N7���0�ᤢ�o�g��&q�0���i�,>P�=9N=V�Õ�����"��)XX S�th<p -��^e2VG��h8P5���/�XY4gtL����Ȫ9�\F�w������]<���l���[I�_�	q�����rn����������0E^MQ��
�I�ʷ���Y-RH���PqO��ĢB
�f��r���5{/(��y�z��ɯ�t(!VU�,�R?�r��X�o¬�~�����c�X�,7�9�qG��W�k��|
��-)
�j�Age=�ŗ0 �2s�� w�A�m�@L�0�����s�`f r+�SUa������!�T3��m2jg�6�+i��D:xj�3��niޖ/��oK�;���r{���G74KϺF2��u�\���p��I�|���A�l�g��ů��4H~<z�) s��RYh�7嚲�q�̪:VVbS�m���\7rJ5�	��͜aFq���Qrx�M��1 �e��d]��g㩾]��NR�ϧ�7�\���ybDI��t�
E�KF<2�l?�%0��5��m;�����A>A���Η"<C�Q���N �Mj��^����H�S�hE�εZԉ�EԒ�$>>1��_�\L�ў<��*��HHʿ~��_�4
En*pQB/�d�m[�����ix��K�k}�;0�د�´�.���K�pJE�r5�v��TrL��q�t�e0%^�d�幂�4L:�R�.��(Z�T�KRF�&�_kQ"�"��D?B�ZZ��ߏ�H�P]��D��%�5�r�M�4m�R%�Ȳ��R�1D��l�QjNg�t��iܷD�F�Y8��o�������
H�Le���Ŭ�?�̒͙��%N��>՞�hҕ�k5%�S晿p�XL2/��Ċ����b+F�������j��}eB��߰Œ��/D
��t�ZU�>�6X̪4���Z��S!K�:Ÿ#z��b.�R@��e���n�	o���`�,�=�^�x��g�)O=@;�r׌8��^��c��}�}��5n��&\f�۹��d�9��M�d(�y�߄nչ�L�ϖo�^wr�ΰ��s�T&J0�g;��Mɚ��}&Z⤷A�+nᖒ� ��/������+�_��>�ːJ��_��p4�T=�M�r��զ�:�lkm�=�����?#��f)?;�����7�`Y����)?�r�h��F+��*��$���`a:ғbN:R������x%��c��:�k_�`��,g��`�/7��Jc:yr�3I�C�,*]��)RZ[SKʣ�3��#��6"�T���K\�Fs��7�YS��,���X�bKN���W�U�-��(�j01j4�Le��5?��K~��M+�����pS}�˻�0�K�h �o���
tU�H��;"��.���q�%~p����V��E���>`k0���4�ah��5G��
"���������_e�����`ygE2�B��ɺ
��<��a��RdAO�S�B����Z��Dz�%��C-�xMG-H��|��GS�O��V,��Xsu̮B��!6���;��6�2,�[�2B���hz�y��e��a�	�t�U.bC��v�s)�sS�!�Z*x�\xY>�!�~*_\�����w]�	g�1O�b1�/�L��V]����?� b3-���m��J�W�v��F`��De�7m�/��D9�l�����d���\F��ػ�K�����p�UҾڰ6��!���gJ0��֝�R/��F�O1�P�>��ܳ�4@3�ǀȫG�cN{�j�}}"V	��8�J|�:fk���L.O	�(GX+��>��K�D���S;N�̋\�Em���;'b���ߧV���EL'�HE�m01����o)<�t>���<�^���w+��z�m�oKjs�@
L9�׼�N���t)ޫE��ɦ���լӁ�	�#��'�w��iq?��fj��UR�)���Q��mͨz�f�hT�aV��B�s�Nc��xI��f苍p�]��m�$yۺZ�� 7���Nhs��`��[K��n
��X�ȩ�.,�I�Z ��7��g~����-o]����>^����霅I׆��a5�ņ��u�	�Oz�,���.�6�.saq���b�����%�ݜ�mݭf�!#�F��e������&�Q�S�MҔ� }�Se��L�/���ۖ�$�=2�h�����lF>iR��ך!,Gc��x�L�Y��*��Zi#=)��?��X5��o'c��RU��XtT�;��3�����A��joju+��h�}��ć9��H��.�������ޭǕ�F
������U_��Ϟ"��3�X�=���WS�W$�ۺ~@�6Ȯ%B��p�J̨\'qiaT����t��.eg����J.����l�@Q3�L����bQq���3(��=���&���&95��\�m`��V�R���Q��9��0]x�����Jࣅ�[W� �72��/��U�Э�ªO)8ؼ�i3�&��{F߁h��d �
��*p���'���`?e9���\������٠g­��pa�0G���H�b�ҦC�arϳپ"�H��QUk�l6f_��g���+�,�"]iT�|�|��>����Z��#��}��X�������=�έ�U ����`=��v�J?�
nu���o����vO}Bl{�8�n�����&-A(q�a �U|ԍ�C�������e����Ǚ���1_���d��]-G�v���Җxt�Md]y�%�XU$pWb��3�J� M5$��_ȪBL(^)�`X�`>��L��c�&]_�C%��SЀ~{��(-wD�Zg��/&��z6���k�ؐ%��p� j�9��4;��L屃2}��KCd��2���l,}**y���߮�"�ߩ��)�A�m[�#�9�F��C��ae���2����H�5�2H�`0N ����P
"o����jvN1�f6+XJ�ݝ;n��X���@˄F��r�O?WfS����
BE�R�Z�����Q=Q��	�Jg^�a*��im*�0�N��Bj՜��Ώ�O�>� ��~4	�3�NŪ)���孀#T����(��F�#Z픽���"1��� B1��ɹ�|�l
f:���Pq�,�~��J�m�%��'=�[��}�v@�߱�/��'��R�ģGt!��1w�)*��� 8�c�mSӑ$���[z�t�V� ���O��A���yc,+ƶ���>�X͢�dνO�����%<Mp��Qi��� J��p+���<<�U<#'T��%�͏��IvM�sOU=�~�K�I�Ub��y�DU��t�^4�u<m��qt��T��$?�D���oq:z��t�Z�!��q?��:�v�<��6f`nMV�����k�ӗ�T�M�gamM%Mɢ]��f��,hZ[?�c|=�����=¯�0GZ�Ⱥ���9Ej�̱�ί�r]OC骙­���y;�ZC��K�n($%d�_��)dZ�5����7+�Y�{�����3�mƺI�i4���J(��9� +3����+pW�n�Z�h8�àE��qUPo����%:��^��W���ft�2�M��k_#������cBX��a��&�R������θ(6��y�������?A���kQ
�B�!c��KρL��+}���3�u��u�|����&2�f�d�f����A���YKN�F�W��:C�UMެM*�(҉HL�8���
���$����2�����(���?��{���V<qI�����g�g�}��X,$E7�V�ƵO��%!�8q��6�i�3�߱i_BO��_��Ŭ����(L���S#Ix�?A�ާ��1Vr%�r�"��q�UOsܘ!式5��J�}������E75���O1�YG��o�8˃rlJ��hx��\~��ȭ����V^s�rڪ�F~#��e���3!٠�h;�u���RśA�E��o�M@�I,��^�4L�!~l�C�ex���D��X�W�&�;�쪸�$�[g�d��T���K�˃����؞1�A4el���9������Ԝ9��a�'ۭ��K����D�����H���o�p�� �n�*�OD���<��Gޞ�n�����:[��Q�p����nD�	���_�4��PcP|c�)��)�m������U�'qTԟZ�( �S.����2����{�"{ދp��1+`q�E2\�_@ǈ�ڊ
��z���_��<Lc��J�M2mK2�pDX�`��:-�:?��B�@�]X��M޳�=��la<�2��N�<��Q6Z��D3�[,ӉJ�2��7�� ��Iۻ(S�p��%�:���	�	+���Eִۅ{�/bɢF��z�'�H~�1Q,�*I�������k����ٱHs5�<��I�	�K�}��o������|�b���tî3B�۟���17Gu��_�u��'b��%�7�Z��I��N���U#4ݳ�V\�3@��Q_�e\�ڜ܂�	r��QRr ���d2��h�zǅ+L�6>߾:���KOU��X��o��̞rDw(�/�x�pN��"C �#��R?E/n�Ci85�۳<,7ط7��=k@�A�&��Ef�^6�Gd-���+�6�!���@U{�;�V�ۣ��'+�@�{�+�nuBi\m��L�a[w&[���l�_5�V��fC&<�ؐl�a�2.���5�����2c�����q���픃w�O�`�`���Q���<-8��i��gX�����O�*�8; T�~��~4t/�\�)���Gh��x��r�=-��R������\�b٣�3��%�k0�݆ڏ����tHG{�=X�~,unH҅�a��/�HM}cp"��P��[�f@X�h�f�WC]����F���Ž��	�o}�a+�����~y��K��'��V�T�k;��t�ˍ��#����u�Ρ@�U*r̨�u=��!���b���0qg��r��Vke~̀�჌��o�<^;��03l�����g3�d��J��ԋ�K�Z���
1AG�����z�D�F��W�f<�]:V��\�+��{8��VF4���k).�rSv�ZD*��Ah��&4�yB8���qSSQ�f-��jbv�4��3�N��6�����[�����E�׳���z���l�ơ��1>vBN��3v90s�S�؜���'�D';��p2�l�߱�|�D���B6�Jl#��<-�㹧�	VL �Y�PHm��^TV���"�R	����Y�X��wv�����Y��~�mOJYa���e'�����j<��®�̻�[��":ƴ�>c:�����2 �~�mdj{���Rc��A�?SFG-�ܭi���ֶ��3j��U���W�����+^��a>�p�����\o`&�F�@WM��@O/�-T� ��"��9O��@�(�P!����/���t��^�r��اҪ��')ߴ>r��F�%<=�|,gl|�24E��;5�#/��A}Y����(� 9G�|�fN=< D>�f@��Ƒ��d���#
��W�r�?��kmT�"봚(��UI�Ó��(���F��jⱶ)�e�N��.y���#��m|8m�M���K#�ȘG���]n]D�1�aq_�}k�sӞ�2D�i�C�ʐ1a6%$��?�S M�J�6̓*,U�E�3�����aǚ/g���|m4�L�@�ٔ�h	�R���=g���f�xvx�5����bָ�tл�Nz���.@��r���ী�5U���q75q��F6y��� �!vz^�ϖV���U�#|��z9���%B��f�c��x�	:��2�؂�oTF\�E�3�z�ɿ!�`
[��K����(Y�\��^���M�-�Oe]�2W���n�x��Ϧ~ �P��K�6<�,�P!q@�W�#c��Z�G0׼CIl`��5��
�����c�j�9��c��Lfj	g��;'����-X��3�0&���p����t���}r�"����i��gؘ�.v�QX�ц�<{ćA�B�QC\ay���@�FÃ�z� �z���j�/���Iu;��͡��)������1��$�u~�����5J��#H�[T�v���]�%SU��؜��x� n���M�*
"w���:kѣ���א���y�2�$	do'�܉��>9{f��3��y�J7����^�e3��CX��(�+�a�8���窬�h|pV�̼����Q�bwB�;��w)z�u�m�4�N&�v���V�Ƽ���vg��S� �@?�;��8���΀s��j^��{�oRb���B�'kvz�}�s�/��)EE��S1ܛ���ŵ�wb(��~ҧ���p��y�~L*�����T�u� �'&���j�Z� j5*3`�1���l����*�v��%����x#_�l%��ެ��K=�IA�y��#Y�E�	V��Jޜ��p�E��|c���=Ӑ[��ܧ��?A"��ƟZ���I5���ja\8��b���/nrZ�j[}�|{�SpX�k�*a�	�I���(��{Bh����M����{�.��������e�m�fǁ3�K�d����عm�s)GY�}�H���6!��f�3'�y����]�wJV˝E���z��џB=�Ŝ�R9L�|=3���D�����'R��g�I�������ט+~Z��S\��"�(�b_��ܛG��d�?�ה�cE���q_?ҀF���6�"(�PH�.�,qƜvjII��g��Q|�� Y�XsX���u�(��M��)�8!��k�p"d��[
�M��6���k���)��\�}�q��^4`�FŌKs�c.���5A��a�s8��O��W�ɴ;@4�u�s}+}E|�XI�(��L㣚�@$�l?�kES}C�!g�뎼����2l-��Jyz#Sl�x�.E����!%�W{���6�u�Y�H�4�J3X�*&v*M�����%H��|}���_�v�
�a�fZM���6`/|��J�$�lp������u��{w���w�:pP�:������BУ�QF�������/y��� '�<�tҬ)ݢ���e�-����h0�s$YH��,��U�\�R����md�p���ȹ]@>F��1��t�p:FS��Q�Z4���?�ˤNGY�9J=��f��ܜsE���\��:T&�x��x�z��jv�z���7+R1����`�RR�����?b�����B��ˍ��R�œ�j���z^hN�I�I��C_���`�����
��ߟ�K�\�Ł/B�l��¸�+b5%9��0C�Bv����tW��ë����R+ɉ�c]ol~"����ub� E���ަ-����iMI\�1L`d+F�h-!\�[q��p�UI���HR�:��-���fi�y;�|���7ޕ�ț7������	��Dz���Mw/�<��BQ�f3rW�X\ry�2_o��{�/��:1�����`0�ɣ=���u���T���uI�W+,� 0�#�A������{"^�@�$�n���R�ɝ��rL�����L�����:Tν��}ᆜD��uZ�n|@���6�~�&��؝�@(@C�"JV=nUd�5�c�¹o�O��Az%�~�z�Ƀ���������4m�>���Ȯ������3X4�"-F9*�4��I6T��ڊ�TS����/	�A�Z!^��daWfwT��!'���ӑD~՗�d�A��	�8�	�Ev�d��E�-XREc��hb�U5�1e�������O,��V���ŷʑL��)��x<bA/�W�Л� ԧ@"���I\�rvW�D�M��,������ҽ%Kv*|!��џ�*{��ֆ���|��V5�Z�Χ��nta��S}��X�9cE�4�@���N���}%�g1���0~i�?.D���u��_R���i���^��v�e��p ��t{�AZаs�,L�?f�� �n���I�%��HF�n�� ��{��4��5JZ�����m0���)TY�>af�"Dz�Pm18�-��D��2�8��Ux%c���}:�Q�\
�u�<�Ir �\m�+u�?�l��z�we�c����klx�9���,�%�_$"%x��$�r�!���cz&H�:h�"N���9q�JF�a�p�����{�q�0Jg��q�-�tr��)a�'�X�hsE�(Q� ��W�MJOULc�\ ���[�M(����bj�wWの[��s��<�L��\�P��𧡣�{g:g[]��F��1T��J��K�m��g���h"��@�7��������~cРS�� hb��U��rɚ������p�O������D�>&�E����gݸ�i��G��{8C}�����.�(�|��_�d�*��#|�d����Fh���}��%�Y�/�Ǿ�6��1%������u'e�v���`N���P��LD� ��?u��X���Uwf�Y4=�O���Pߕ�E����.U�,�I�����$?@��e8�=h���ob2�j�:��T���`�KNa��U^�
!��Ɨ~re���x�ץ��>-;�:V��g-dq��q�$}\vYs}<�ܺ�ډ/Զ��(��*���x[�������n��SqX�y*���O��R����h@6���篋��iƬ��m@0_��_���_��������u�$6#���bs�\����i������Y�,"ȥ9y�|� \!�/41 ՜d��x�QL��}u��S�lD��TSR'���6�䐽^H�Д/.гJ�aG�5����Q���@��d�M�Ă�Z�p>�+>��<�ԏ�I�S؜�?�@Yժ�y���)����(ȇ�NА���o�m�3�EB��:�گ7<^]� ꁁ�Ln3ݜ_>��<C]���վ�����UxC��ctN}��(i�F�g���eئ"6+Xv���8uC+)ԩb�SH?--�""��p����ߙF�k���1Zg�	�3ݔ���ۢ�k��*��[Ф,���/�6(ݖr9#����Hl�Ł����Dt�a8bS\�*!��-I��}�g~�m�u:�C���R
�A��R���e�p�'-
AG��}�z/۟9�v�����?c�IzELy�x�÷k� ��,�k\�{�ݳ��U��>=>�!q^�mrh'/Z/�e'��x�Ʋ������|4YCM���	���4jq�X9�:��O�(��Ʌ#�_�R�	�����Lx������qF���$�#���ʇ�r��qqU"�Fa�!1���R�ԙ�=4<Ϡ���z",�a�m}oݔ!G[{�=t�f��wԷԨ���u��ދ��<�-�r�ٹ,7�!p�M1#&�"6�)
�Ie���1���E ���[pB_.@��N�.�98�o0��kM�A�	��K*<0�tg��	lΩ���djY�Q�ٰR����[���;�p�I�S�dvkbY�4/�[���G�ֵ��4�������D8������dJ�_�� �sf%�4y
���w�����M 9��� �9MӶ�J�7��ٳ�Y�xrU���:�x��o�c�V�В�z�r�T)����˘��d��˪I��M13�~aq�N6��&�Fo���5��Y�{���|ȟl�`M�Rz=U� ����T϶�:T<Uk�' 4�N���C�����>�s�a��!�Ļ$}��63�LN���Ql8�x\�F��2\`գ���EP��"��W�����/�����D�i�(@O��1�KˁC���($�+FWw�����o�š��J+ӘQ���2ɞ���@�C5X�7:dW�YHʸ��JM�;�},�	5��s����Ȫ�R7^�#��_��@14�ϴ��	�(<G�t���8%s�B���(^z$�'C7��ܣ�{��O�R���Xz��}����*��5��d=M �������0ewt�B����������,�|ayo���.�'5�nT���|��*ns�qx��F%���g��hgX�rWg�sC�9���=n|(��t�Uc4�~+��{����3/T��Wk�f�g���!��6-V�a���=j����,��/V{��_�J��40����㆒4��(���StJ�}A��_��H�&�ɯՁm�^U�I���KYZٴkP�Xd~�i�qޫΑ#����Cۦ�e7��T`aO��+�uwF�* &��ܷ7[U�A��=5J�9�
x�����LK�Dk�&_~�*4��鍰r�����`��I� ��	*���:8Ò��h'�=Jă�<GD˟���`Rb�j���.�'�T�o���1���<*��v�$��}W�t:�kj�-(�|��Y�+�or�t,o��.pr�Ъ�d����uQ��/2�����ދ,�$� α��q��U��+��,t�|k��w����+�$k�-^FI�jzK�����59?��R��JK��}��2޻@G2����|���7��6�5)Ӗ�B4�9��X)�R�R��Z+�;��⏴�]B�[۲^�)\�`\�^K�(G~]:Mt-_����Z�)����J@�)9�Y}�ݭ1�t�����?���Ї(!�H�Ͻw�*�ʒ������ �#e�$�Jy,$�qւ�"-��
��M駷�y�0�]�Α|��zh��T�AJp^{� CqR�@x'!0(��M$<$i$n�k��� !C0�f�r����1k��r�u� ��5�t#QnMC���y:
1����5j��<�\bx�f��CzH��ޞ+�f[f���L��~/���]�6B��H���k���`S�v�ӵJ	Qڶ�([�����X�IJ��.;r�T��9�\�Y�(�<#�����ku,�����X([���#t2�0�uJ'����<���?��|d�(�j��֦�2��`����=!����/K^}���Ү�%��X\��7��a-R�E x�[2Y�g!n��& |��,�p ΀����\/́�{����.�\�n��j֚Ҝ�>7� "û��oA<��r�n�RCA���{Q�I��5��z:o�Q0��.J<i�V~�u��r��9����)�&奰��#���o�Мs��Mí���X�c�I�{�K/Lܒ�"�M��aK�%%Px���HV7�x�v�R%��<���g��\��Br$�1*ׅ�R7uځ�7�8#���	��s�d�s�����t���eg羦o�g%��6G�kr\d�.^�v,|���耟�Ո-#�YEw;���x���&,ܯ����2&�̂�~b�(h'<�mgzp�"8��?h4)���(8��?m�����x-�!P�)�u()-;��L��-��J�Ę�^T�|Sk��V�H�,_�ˇ��|jv��?<y�M�Qx���CX��I�����
����G�rS��3hu�H�yN3��w+M~?��A3z��(�X�c���}���ѯ�"?>rK�,D�A�	2W�r}f+Fł|��X~�n�
{��G�W����	Mxz�Pǻ��n���q#K�3(�*�5J��}���OL���5��$[���7��a�P:��+�������&������L�&�E!꫚A��ir�jm���Tg=�@�$j��!Ũ*���iv�y��| ��*Ϟ���{[uW��-�^�x�!����f3�^��y~�����%T�P��>�B�wEɚ��؄vȶ�0����某?�m�݀lipTUƗ��:��R�
���ɮ��	����߂;����Lq����M�
��4����96����6ಬ+ؠp2�A�ozUV����U�JЦ���j�����~j��A�YTT,a9D�k�@_��b�&Dt�s[��ͽ�J���[f�L*�qS��S�p���$�M�C��:D�:���+L��]q�Y��}TG� ���o.�� x溙T��!�b�׶W}xK�5=n!�5�B���I2L��L��)��2��u�mו�d����0����ǥ����h"6ɇ\c�M�db@-�p�}���$=��5]0iK����^��'��`���b-�Z���K߯�Jҝ�R7�_������A�W�GI�;{���w.��g؂T6�.h�k�˴�?b�"!B
,�جH�Q[���(!��)p�jH`)��
�v���h���V�p�]��a�%�R5t�^��� χ�G)[�ѓ]b�e�.��1��j�7��P����.��6�&@pK�l��0�e�n�UhƱ��ŋ�uѮ]�3�G�,��ؗ��:Xb=B�46%E<���HSt�ߨ7�{������0ٶ�N�߯��5����p?����Kq�]��t-u�'��qˑ�M
uT	�%��	c,Z
|�o�h@�7��y-�rn8�L��QW8����$�py�.aӡ�rHi��փ�����oB����$V�x�և�$!]-O[��j��e��H.#NM���1�ޓ̕�/%��n���Y[����9�����nx��\�U-�,��/����Z��!���L
��x�4&y�&��O,��/��l�U3��&��`P;l��A���4����	�Ό��204��tX������!m�t�E��-ϐN�VM����7�� {b�v�2�,�j0���z��$���N�M��0���%b����ɚ��$����բ5V������A�+�������,����\��-#��[h^�]W�J�_}��Lk��\LEE�hõ/CmF�I{z`�=��JJ �<�qM��z��j0�kZ���`_�",:{���z�)���b�U�<�Đ�^�Ѧ���[��9U0Y� '�w/Q)������ŵ0l[��W�o�n��]A_G`w0?��DuO�!�y
��>��]'�Oă�����f��M�bX;�0O`��N�m����Q2UX~���!T���m���Y.�/������]Z�������N+I��ӷ��&{�0�V��5��)R��~9�?ܸwU�HC��.�&�m"�G5]�C(���7�5�JE�>��&���F'���jq&��!� ���M�(�OM3��������:l��Q�a��y�?�,��� u�va�� �闚%Y�?��$�4$��yQSwP�{�v2:)�{C!��V�)Ƃ�&��,m)�7����9?G/֙:vE�*�d?BG���m���t+�@�X):b�n|��%�+���xA��V��P���SYGA9�ý�:2Y��1JAjE���O��1j�
\D�u$�K��e:��tv����	���EH�m�G�N>�X�4�˵qT�uj����x`Tǆ3>�M���3�4���Q��br4)�Y�Y]daݏ��$<�l�
���� �U~��JА��=��r����:��_:���d��� �>�f�@��%ܧ'LKnW��q]n8]���$����=��lx��:�t�߇��a�j�N�5�l�΁t�	,ޔ��vYFˣ��fx��靈�D����d�У!��Ũ��̷q_��b20��z02z:�̓�_a:�5�Œ(�%�x�y�;	Fs_�ke�n�=����u�l��R}N�\�_tTqs�w�
�C�5�=7������C���0�W�N�^�RX����9A�niv�B��5��Q�(����ނ��Eh[@���rS���M�1����9����0-R����p���y<�{��u|Rg&��5��bj�Q��Q������~����0���^ ��pO��r�5О�$��	\����m~FH��<�22����GCL��֯�+Aބ&��Lh?�8��ٓ֍���Y���(�����Y�n���/Q��J[����+��?�d>I�P6S��:���T92~�*�-��x�U�!��(SL3��\���y`_W>���\�'��1|J(B�7���Jdۏ㦥H���$�#
�a��(\�j��\��aG�0��U����*3���W����ڔ8R�7ѓ�,�+��s.pQ^��$F�M)Xm��G`�.f��=
��@�F��*�^��ں�O]�m-}N'�8���n����rіd��`@����k<�fY�b&�U�v@�������������QW�g�Y�+��.ZzШ�*_"m3��A��!�����l8LU�Fl�^FcV��1����g�V�9?�w#�q۝�	m+ظx����+L>M�L��M[��wh����P�V��:�|�Ȍ
a����#�y��g-��}0\}@mj)���[����,t��tޅ����O�+4�X�t�!����c�%ҁ�`�p��N�Χ�"&Y4!W1MLI�ش�2Q裭���:K���h� ��Rs�jU t�v�m�,�L�ʤ��<������'2Y�5���!u*%���:����H���l�^S��Fr����0s)�VtN�a��)�	9�7���Zd��AZ�Uv��ormEÍS)��3���M�R�9(�CM�ଋ5l��g?�y�8�(Ѕm�[�+b������\��ܯ����&E���DD�=E�©�޳Sh�gi�ӲI�?.��y�R*{��nW��&y���&�U&�4���Hi��O$��^J��H��ԛ�@���t r�����sS�$�H��q5S���� ����x�<m��+&Oz	�u�4�
�LZжK��W��k��^i�87�Jp��z�\�
��L�OLA�B����{���UX�};�G��1�f�����:,�D�~��9�>��Ƴ�.��ZA=s���C���AJ[�P$�S[/7��
��Ղ<�gX�����K_D? Y.e;7�q8��[?�i�UK�m���%6����d_>����GR�Y���%�w=����tv`�mGu5����j�픮��/[�}��i��,vM�w����O�|�����L�w��׌��)@S�� ���*�����p��F�x7��B���2��L�k��!09���X���+y��t
֊�0�����>�j�vS�Yty ��:[��j��3�>�.�Ogae��qy֙�L�6`.���$i5pM��;~>
���m�.Z�W����(\��"��"w��]2+_:G�^�i$ؚ*�ħ3ͪ+?N��U��Y�$~�+Ŧ����,���9��$w#�jZ�ɵu׭$�e� G|��1�\ȃƞ�"5�g78��B��?�̑T)�e��f�7�B�3�hGY՟ƍ
�3����|D�A����Rݐ�R����h�S��m�ě����v��cC4R������y�׽�<j$����0"���֝��W�
��ޭ�Xb��þH���y��9�(i.շ�����
~CrB *���z���\s��ʼ\���z�� �$$���ZHˆ��`���4n�H���I����;�zհ��>%�W��=9�H"@��`��iIBT��G��o��Ua �X� )$I*�:r�Ja��J񢂇u�����៼EJ%ث������V:"�1��8�U��#�N�*��o~h:��Ҽ=k�(�Y�*��D��ĕ�«	�>�vq���@a<��a�Y��DC{B���`�P��;p~�����s�0&��7a���� b���($��2�O�qQ{�QG": )��0���r����_����埿�\�{%I$��_���>�|�k�%��k���3xި���֊rH�-FI<{CgT���$`�^������1*�Zݠ	#R� �[�!a�Vq7Y��~�u��feAt�u�Hz��;+�d���_�YXL�]S�I�Է����Oh�	P�TK�����S
2�� �p��O
��7�\�)��7�xi���E�	a��,�XIx�C�n(��<��[������9���x?3_iQp!���%�w�5`��Z�����r ����G��r�Fi,���-�`�ŉ*�L:�0�y;�-����O��8�#l�6޵p5��jp���4K� ���q*eŹp*�׆_:n]8�:�f�A܍�,���۹�&��{O4G��;]2�޾�H���.�oA��o�O��!��/�(*?y3�\�
"1@nW�#�ت}�]<=3Δ��N���t|��x��^I�G��N����EΔ羻ϣ������+p��a�O�`}��v���h�18���d����Az%0���J[��\�\�\P�#�C3��z����>�0��<iG��_�7R R�4�~�7Sedh(�\�*ɾ���+6Q���Y1�Д�Uy*����y�hMI��	�����t�w���?Z�q�L�	)-��f�-sS���N3ԏ%����h�{����5z��m���@l��s�vi}jG6�i/D�iK���ƒ��jf/'�*v��/�az� 9��cLu�--��*o�rQI��ʵu�н �"I�[��ٔr7��E6vԱ��	0A}�<8ݪXPn�����%W��G;���]j�q��ǉg_� !�G͢�r���������`&mw��Y�g�������y��Gf�}8Џ|��n�P�[`ʚl\������|<��1(���Ԙc�o؛K"���Ś�Ea���y�F��ɗ�H��� &��]�AinJ�cZ�X���Mn���߱���q��5���?翿mD�Kw��ZѐZ����7$t6�!&��sJH�`�怘���.;��^�j#V�(�� $m���S)Ha	�yC���S]gU�d��䁉��fhG�eUM�r֞@S�m,��rD�����5l[��r��1F�!��j�5O^&f&jT`(�U�r�'x�@�����h݆n(��7n���ˇ4���3��^�&��]G��E�.zC�2�F�C��������1�$�{��8�7B��F5�1�s���u���έo �į��?�ǡ�¸��w�L�#�;�$���S8Y�b�j��0�d�̓�?HX��Xm���X���F���d!%�H�� <�y�h�1�(�t:@+���Fd������}?�t/	����F���lh���Rd@m�o�e���_w ���K�W=D��7�;�����(�����Q ��ӉT+���E"����V{�(�#��K?�]��W�-�Yʣ��4�]�^d14�~e7�.p7.���)~�q,�X8�"w��)�N:[�3�ru�BI1��ui!~V�Zz�%��j2#e[@�Cm7���Q��!�sP> iZu-���Z:�T��`di���r���H0��/ǲ���R��Z�\�,,�����ت���Zfw��#&��� x �(���/�=-A<K�_E�>���9�og�ۭ5�!�4Ĭ7����B���a�z�8fo!���ij�P��+�a�&�k�&���LK�~�PBW��bPU�l8KI�`� ��3����Y�Л���L���p�i�S&]�����������RF9��=KK7�"L���i����^��|�w�_��v�$Y�- �+����2���5Ѿ����=:��1C�	�E���lͻ�y�~%˷�ᔢ����/���93�C~m�'=��ߒ����~U��;fn����}�Z�3t�(R��2��*|��T���G��V_�8�3lɁ�t!��c�M�"���h��B榳���%E�)����#��r��a���U9@?u�";E_wyk��3����/'��2$���
0�8;_z�UҰ�dނ�rV�%���R��Γ�7d~��{7�*^)#�Ǯ�`W�j����kڶ!�t�-��];pX,����ta�Zf��-��Z��K1���im;K��G{� t�1蠍?����/����
�~+�~P����|;�%GZ[�.��&/]�ۖ�)rށ;r�s����8ˏ��u�i�]ȱhE9��5 �p��Φ�\����VH�L��\�6�~�4Ȭ��������/�Դ:���v�	m�מ�z�Oa x���z��lIN������h��R��h��Ol�C��s����W����#��D�7�,Y�醶k�����v�bN�%3��*��Tesr7�I4?��R�������3������,���g7�us���J��{���)�\!�dk�o���/1o��
�(jZ�M/4�*\,جt0��]{*��}�bď7p�W.���(0��Q����$��-�
u�Ļ�:�p��j�P�w�aF."����(��=�>8��< ���aꛎPf'��f�v�'cW�f��	7�q'��4q�|88�Ԏ�j��XȐ����HrߒT���K���U*J�72ֵ��$O��PM��c�|[<!�9WJbq]*V�J��Q�i�m��Ų�aH�v���I4�΄f�~-�?@gJ+���b�'$�@EX���&
%�j{
�
U��V{�R$"�%��k��M.�k�b�FA��M!��C/�"��i�����-��W��ӫ�r�f� CUrq��� V��.��!�[��c�rʈ\�C�x�J�_��)���KX[ ��%�_"�4Z��C��s�fg��cǑB<k�2��ٓp����l{*���@H�|����{˯�EE�f���4����Y�J%��p��Rږ��h{ƲQ�7��'(2"/�u����Ol0%/Y�3��Az���� a`K���v�@���{*l(�^�f-Yt�,|!K�Z�Gr}{ȈK��f�YD'3��naV��,��pqA��j����|�L��4r�2Qn�~md�l��wAZtw�MQz�PbN��.�G��Q�ul6L���a�c�I��*.b�S�``�qw�%H�V�Ԗ�|���Yd<M]OtfF����h
�f`�4{�o�	�,l׹ĺ�Kx�W���j�hԷ��a�gb�p��˝���0��@8���1G� �,��J��|�[�W{�͠X~�1"1s7y�퇇�9QSڍ����xƁJ6��sn��h�|��xF��.����#�ůMŮ�	���K�.���sT����n}�6�r]_ޢ�ZS�V��|��*�O��t* ��W��K�]����z�n�'&xp{���x�G�C��� |��Ȫ�h_�i�P���1�G:y���PE�F=��2-A2�fZ��i|}Eb��*����0^LSY��vhqv"^�a���-��z;ͦ����鿻ᛓ*ѯ}��i�%E�k�KW��o�S.�j�9��(a�L:c���?�6�,g�쒋7�f�L��Q�����Ķ��ϝ����/��I:'O-��X�c��\g��65�z#de��r`t��d�Re�+s����EhА.m?iU����J�$��7�k�o	Z	_Ld�n=s�߲�λ#Bo3O���f��z�_��#����ʚ�Q�ڰq�oi&�+�����Rs'Ioj7�I��KyU�4Q��F�%Gp�^Rv`6T�b@.��CB�s�N�����#J��Ҙr�k���!�Vm��8;B>び�S�;g���ӇJ�j0' ����9nC+�w$�4����XG9�ͨ#�&�6j���o��z5T�!-ĖQqc�
�Rߖ;4�g����`�!ȟ�� ����o� WHՆ
���Qr3F|f���*3O֑��u���yV�����{��P�� 35F��	}���"�MS�&��F�.D/��b�
ۥ噋y�^���J�2%�����_O%�B8�n~VY����H\+���S� !Ҙ�6����8�Y����$�CNh�Ua��?�2Mi�(A���`���^�/�@y(�Bx/��s���n�-���d��	��O{�6�������� �O��Apļ�(g����H�+!P����ܡ����
�t�x�4n��N�-�2VX}h��Շ��;�����
WԗB���e�θm��t�t�ur���>��>#x:��hG�ܶ༄�Ð���?���� ��AƱ�h�,�X���p��9K���Ęe��±������o�o�/rFnq�y	���ʼ3u��2Nt�Ѧ�R�ٳ���ލ��>	S��@@+���Cߠ�����
!���������ߢs�#��^5m~@h�i����ɾ��]+7��
����O2~��#PPXLg+�gh
Ċ��E)h�^n�O"c�vS�]�֏A^,�F�7��'�[L�n�H�,��/:�"�Bkۊ���;�)q,�y�f�S�6R3&����/�zp��p�Zqp�@��3LԦ	���>�ѫ՘댂`�l�4t�+g�#2����
�\�zp��(0�`��4	�����r7���{�'`��PB����+�ccf|���(��A(w�8o��	:H�\��;̨���ɨ�/�IV��F3�j�^"?�.�Đvq�;��8�X�e���s�<�7?8���#�����"���3�	{WÂ"2���hR�L��i��ܪ)�ْ�\�9ϼ-9�du�U>tQ0Sp-3�<p�5|�H��>�z����V<�"A�(��|9�s�̧k	����@��������z��>�M��5���ػ�Y��ς։�
s0:�i��免O�$)24��HM��3�}Vsmnt���u����}�t�4���:mΦ�@]U�ve]f�����U;��A��W�}s���f�oHwm�us�G�Q���\�c7D28���3Bvo���-1�h�WW>Ɩ�*��1�G!���������H��i�ҩMb��$���[MvU3�_Aw~F����!���Q	��rm�1�.O.b�����S	T�&�>��$��,��%!L��:��#�کBI�����ʶ��QOڤ���Z�blPǂ]��f �c#᳦�Q2[����G��H�%*�gv�������&;�-��k�mM���'l_�;6L<���`��Ղ��bg�"pn��x����������XQ���.g6�c�����h�m�)��*��T����V|�R.A�����ar�w������O]����<U5k�x1�V�M�^���Λz*'��sKmt�B]2ca�rw�J�?��Y��?>�5��ZT���O��bb��!��C�9nx�	� �*��龷E�?����x-�3�]d�)���vO˼��ȩPJ��=�N7�G2 n��i�=Rޕ`8����~��X�Q��������=rD���X�,��N�|2�D)/aqL;���	�y3��;�W���ZB�DR~�sz��@�]�e���r�}`�*)�����&���c6Z�'���qi�o��]ɵ�	��Jl[6�}0����W����-3AO�]��UE\zTH�0v�"p$ ���M��,���"�����oq��� �?C��!���W�l5Me��BRCC[�\�&oS��v޸f��7��7>Z4�-�ak�0[�t ��	��x]�Cls���@�@��'�𼢕�������͚� ��+'��)�T�(Z���d`�SdoϷ�	�պH��ts!d̔����S�V(8�6�H���Q,��j>��`T��=� ݟ!^�ݚ9wx�}��*o߽�����;�*�AP��xܛ�3�WG�)���խ��;cc��_"���ZIS�%٫��x�b��h5�२��T�x���a)�C	�T���]��h
�B/0�*ׇ
%`xL�f��hy]�)-l�!�Dڰ��[��$	��������p����	��gi�0��M�\�w���ٚ,Q3�%��| ��[t3=��z�6B�ڨa[��_�$Q�t�2�ܿdd� -�t~鎏���
E����nD?~����$�*�!Clj��H��/-ө�}پ|��LV�5��s��7N^�N����'�}n�b=4������;�z��R����06�9��NBS0�96Fգ~FK���6�
e�5�Y�>�o����{��Up9�Et��>T�-\�g&�4Y��ˬ�>��a���N{��^�ɥ��t^���n?^9�c��j�Q�u% @�v^t���J�j[����:/��Hk_��8O C��D-�i&$_�}�a�<�YM�9�K��r�
m{?�
��ͳ�nڣ�Z��/�� 5�L��'-��e`�
�rH�5��l��j�v}���RC ~� �����Q��S��Q�gѥܨB�#�O`ƣ^�kI��A�,[�2 ��e�ª�Z@����ԩ�]*D�"ڇ��MZ]mC���O��,���'����D*<V�J�5�϶��AnB��<�A��۲�^�V�~� ��b�c֐�1��QsF��V�2���"���a���},efD��-����L�j��:K29���dǭ&T#�d��]vꏪ+
}U]è��?e`�>�� y�N\H'���'�Vvק[��B= ��FP9��#} � �N�j�{���3��aqt8��ua�	��B �kb��r	��=E0�Z�"�S����RL��̦��e@՛?	|x��4��&��uV ނ,u�����$�kYȶ`d��-�W�?��T�-�Ge�k�r�����΅�6�L�b,*)&j>��9��#(�ڼ������E;pt�
1��ޡ �*��&�x�w�(�pQT�q��i�*2Q�U�a���^3��q�#���T�|�R��8D��~�NA����䳬����Bi�~�F`���-X*�L�^��]~������i5g�+{Nx��权��OY��TA��:�e.���ƛ������d��&��pPJ�
�z�_�ʃj �I����ތ~�8�
0�*�T� #;$D��y/��ep$�\V.Opd��$z񟞷J1�\�b�g�>|�K"��L�hh7l��s��̢�_l�d�|�?j1t�O����"�B|ģ���N4���g��1]��ol4��n=���t��N��}E��u6R�<ijy^|:�e=,�PE��e���~,��R,y$�?U`�.2�t#&�g#'2�l�涺�B|����$�P�w�j6!�p��m�8āpNN0Q�w@���g��"�m'7��RV���i�U�ТxRƵP`��Ye�붮B����.,ؼ��G��]��i]��a+ܪ�y��UeE"j�W�V��OG/.���8m<��TW�W�{!��RSu��|z��}D�k�j��G�C~\�I�CQa(%��
��1��<�^hT������݈�#�^#�u��@�NID���^ �:5ɡ<W.�a��i��Yzr���m"����aM�O���ʇ���K���f��R����f���o�����U�#������Hܚ
�J��(�*�\���{+c]g�������]V�8�g�og~�f�i l������@��n���@�}eQ?Z��,�gZP�ӻ���x���O�)|�~�0�Ӏt�el��鵟`���:�L�=��M�=څ�o�]�[����.z��n^���s՜�NK�^�8�D�WΠq5�0�D׋�7܃����T�X�֤��a��Fr�02/؊�QY��~'����t�b|���2kR_i�H8��>�+������K-��4A�w۹�%�:y�u)b�BfH	"'�e�0Г8� ���+Ö�zs������� [���!���ՙ}S�)Ɏmv�4���3^J7
�:5�ᮤ����q�\Yh�LC�=^�i�+d���	J�	<6�
9�����������E��"�-���W�!b�+��3�M%��u.Ce���������C�H:�1�.��B������\�}�EG�1��=s,�'��R#�:�o�ˀ'K&�Cj�?8 V��An�x�)#�e NO�<����;>�*r�6�$i�׃q��7U<��k1�(�?�Q����eaJ���_���t�;9�K�� �g���/61]�x;*B�n~�c�_�j���QP�e��4B*��˝㣲ؕ���$���;�������|ߜB��'��vw1�U��aE|K�KJ�7����;��M��nO�gv�}�,�l����R9���K/���GB=������0��8J���˩]�����������~��7����^W�o�dx�m�4�ζӠh����[��ud�� �a��ʾ�3��m�}~E-��G��`/��4<�1��G7�W��^ha�s[Z8=B�����`m����r<�]��R��`�2��q1�=�Sl�.[����'vf��Yw��
���c��4�܊�w�o����s0�2Y���@�*���������[I�D�c�.�BQ���O���q�.�8����5�ټ+��H�?-s���`�a¶L;�g����zum�Ȓ���p��T���T5��
Dda��4���X
��!�ǀ��U e����	���p��A���_D�"��� ���āST��{�b�&�~o�A-����G݁ș�N��N�O&\�;�S�[p������S��~YC�<���� �o4\/���G0�;B*�ݓ���{a��%>1%c�+q�߹������«�+	>�˥�F����%i���:�^Qy�7��D���$����#w�V�/��k��3J�~\T�djc]C>`PV�4�B&$ĄI�'as�h����5�w��t��^_�Gcz�Xh��d�~��4��~�ZuU�Y
�u�`z���]��6�	�7߇m|�L����g&�(a���ã�#(R�M��HZ��#Bj4��|i�!��W~p	�W׈���X|d�4��)�go �Xh�, ]͞��]�@���nb�[�ƅtmԅ�����y{Y�xҰ> ?�s�<�C[*h��~�ᵝz1����Q���9��4�p���1]n1���a�7ۃ��xP�����(�hL�v�������a����*U:jѸ&�?�0�ٱ:���B�T�
��h����=��'�0�J	�Ҿ�Y\���ۍ���:^��/�ڍ:��~�aѮ* �a��ck���ʞ >-��~;���G�w�i𒐩�eR��G��V��@�
���u�k�A�'�<�R�����2�Wb~�B�2�<oJ����v	���r�e_�(X4�x���s�:��E��9i�NU�o����'�5͆���	|���bZ&}�\���VUQ9��b�K`�3�d�v��u�<�����>���\-Zw@��ʇ?�)7�U�&��Hޠ�j��{r� ���E"�u fZp񃡎諯0�Z�S����A�F��u���u�'�q�� �!�NI�Ҹ.!"8/=�Im1d)�D�,�e6�t+������;�k�b���/�U���d�';p�)=.��.{���B��r�B�"=ԨL�i5��(˕����҇i�|��+�C���9�r}�1	%���yկ�g����"����dx�ps@H�2#�b-�����F����`��R���涞&��e� auV�J܏�{�B�d�.�N�]�Sh���#Z�E�Շ���/�9#�(O�r�kB���"�6�Q�7�F��/q┒˟�N��?��^�6��Iy@s$D� ���_��8����DKO����n'�~��Cv��Ԍ3�:@�mɜ���1�6-�\k��^�T��Zb#_�&:D�l���f5�u|9�ʷ6�s��~:T.k��<6u=�	��VΦ%5��i'�T��u�F{/H�0�dӱ�8��?�q.u� j�)܆�>Q!n�[�Á�*�]�0����#�5&N��#�BZ�,�����|�G��A��b癱W�������ʊ��7��n�Xz�
���-	"LkTa` �AoP(��t]'�E�,��oj�t����Z���O�1bA��c.6�7�rDAu�P|֮8T?�4�ƅ�qp
��|�{�	�tU�:�B�fP� b�{��@��7�Y��O1�&�����'�7<gJ�8c-%@�ͨsD!T���݄�5���q��m��U���f�Y}�-!�
:��[my7��b�],럔��S,�ޜ�T���S�FK0�+��GW�ڬ���VZq�>���ν���¶�(ϰoQ0g��+o�	�-�8TI�S|�^�2��Jԗ2��̍׳lS�k��?��T%#���5�� 8�^&E�1+��,P= *�bJ�'cܧʱ�,�y��O������ ����������mv��g�b"�)}����g����H� <@�YO�{W�%���ھ��8M�J�S�-{�*�!�|5�g:*�� �O�F3`׉�1`
�f���IԺ�(�9@�u5d������I ������?�C1���!��eB0,�iEf���]+���G�SR���҆G�\l�,�♀m�G����+F��)�Et돱թ-��`K=t�v�Ϲ��!�}4��<ڹ|�5��*�p�ֻ%��M#�(�p�&i��Cʸń�*�Yz���ٯ{�-J�'w<�\?p�L�,��X�=�U���ɨH[h}���z��F�R݁�*�@h{���5�kR�>�j5�w�w��fi ru���	�7*?��TR�2�T��Ru%&����u�c���nQ�* �Z�舉�����[T�]x�^�SI�k����y�C\J(m�+&wK�5~�	D���{�ƀ�J0#��ܶ�J3e����^E�\bs�%s�(���H�a�1,;��7��Cí{��.�*)��9�)V5�S{�	,M}��"�y���rZ7��E����V��jY{6��0�k���-î+1�1��ha}���!`jݶZ���W706<;U^��4���/	�0/C1Jb#�y����F�jk�闩�>����O�з��%hRl���$`6(�Bݡ�AC�6R}�������N�H|�ђoB�� yQ<��fD��8g$'k��="�C]���:V�^@�a�TJr�<�]C�p1����E�=E0�@r��o�q��l���BYNe�S�a�Q�^�g
�6����ekTRE�1זp�7�e+]�-��h�xQ dmH���#���{Ђ�~u���[F�]�Mѯ3 UL�d�@wM2���ۈ������緦��� �4��O�,X,	�j�����{B.I=�EH�SH�0���6A7<�(����z d%�)��FV�T�:x� [s'�7�m�b���F��R+c��6o��>۔Q�U�˴�kPoP*�9����d`�ۍ��B���a���x�S��}�U�Rx,e�p[���*�zD�pݬ�6���ڔ���-�)�IH5�� �%�v��|VO�K��"r����ޭ~IYW��B�2W�O"��
�����]�`�zE�]���:�s;�M�����n����ߜ���@��[��A�Ea\R}�'�I��%g����Ί�).O!-�f﭅�&cv"�Zx���M��)��A�1���?[��T�]���*��Y����iE=�O2�VEl�"n)�u��H~S�>�kjxd`P2WN�Um}#��%���AH־�/� 8!5u��`丞:���6���[��؁��%+��1]�9؎�=�`zU�YU��#j�D�\&�ڱ�Z����R�B`���<¿���u�K.����eS�E�����������UK��B+6�^�+�;��¢|~{��y`�<8-��v�h5�Qm�	�P���'?cw�����ee��.G$0sf�����.�7���8�9i��_|@�F϶� ��W<¢q8'7��E#��x��{�C��}|����(��O1��?��{bU��<,�z�ES�� �^+�;�	qC �\BT�܅��#c�˙M�|�P��Gz2E5XF1Sݽr+?)��w)Ҥ:D����\E��G��q��-�AWr�zD�w��W%�����G �Jc���AKw�sJ���U��$�@���-3�9��$��Y{iC xU8��y�c��e�A"eg��X7Ii����M�X�����{�k����*T9�
�/Z��B�[e���D.Y�"eSnS�Fό������z��IL �M��ƙ)|��8[�96hV�)"';:���K\~�bJ{�.�J�sW$8�P�g݁8��=o�hb��O��[76����e��4��DW/��[Tx
��@)F�{2@������I��c�!���&Á��Ɯ�kgG�R�ٞ�����z3Mġ���^gT�F���'<�5~3(�������5��3[���rI�=���?�w���
$_?�l�0���, ���ɶ�ذ�/�[,�� �ˢ�'�;��$	_Ԥ��%���躀yΖ���������-��§6d!f|�Jz5�������2\��?��h	��q����Qd}y��ĮL��m�E���8�=ܸ��c�u�����01X"��5a�٬v��^ٱ��Q��}���7��L�<w|e�x7�gպ-r����<ϴdl&����#S��;}��s/I9����啕9+ߣ5#L���N)�\.�"�(�B�0���szu�_]�!ŧ{)�Ο5�.�;B�G �_0����Y�7]�Z-s��d�|�BE��0�W(�����?��D6��iE'<�	r����a�����OmO��{]�1���y?.�jdIz��]�/���d[ٔ��2��9�B���g%��} �>�w��x���[�t|`�;����Bۋ�_���ӏ�Թ	�W�=[`�DGF7~����P�5q�3�j����^���v�mV��M�/:�Bލi;��5%�����ty��Ez��k6}UPH����'�25/�����XƽJJ���?�B��#�`$�q���zV�
��V���q��	\��cY�:��� ��� ;��e��r�4��@���������GKpr{"��"q�u�da��W�ɶ�G�Ϫf��*����]s��`���>/P�8Q�J���RJ�:����;"gF��Lb�?p�(E����㹚�PR5_�c�B4�{�s�h�(����ہ�O�޻b�b�HdpW�����J�����FWH���_V�:�?�٨�5^��g��i�v�HPK��>g���Jchn��_���"���R�p(�1�ë�6�굛QS�e�cY�8����� a�8v�%걪���GX��Kc���[1%w��Zo���ƾ\/p���!C�l��M������M�h=-��5��1�*�e(B��'��wEI7'�iz��pfr.t��[��7VQ�vC배���΄��3/�l_K)g_�E1���4���{�P��h�&�����`hy8�����$�~���0��r� }c�]%K��3�'+�N��74v����*�����U����-�2̥���ۡ�K�+���q����C@,��<R���U�+L��:�J ����9 w5R���w��r��m�|N_� 3����᎕��H��(�#�mN�AR(��|ػ�h��2�%�DZ@�E�#a�\iԈ2��Ҕdׯ!�
?�:޴�|�91��3�m�5���2����565
��'Y��	�G_>���h�щ�&�T���Q�'��ݘ �3v�g��B;@pcs��c(p^���S��m�����a���mV��������%y�Q)X�ί�v\����g㯩�D�s����.A��Ƽ�Y� ��Ԍ�u�^u��8���#���R
C�M!~�R�'s!��Ꟊ�O-�t�C�4ST��@#�8�źh�yF�D���W�'�v���+�nb�g�*�n��@��\�rd���~��iR�RY�3!.v�!>�&I���	ׁa)�D���#�)؞��u�+FM*'����
����B�tQ�1~7��kT�� d����ݽ!��RbL{W��뉊��~J�G�vM�vc���ݖx�/4�-P��ã�ue�wgw-�W��?�� �H��܂�O��%	Kܛ)��ҹ�d�r!���F��ɝ3�т\�0����r���3�m`ó}��U���m�n[�Q�
��YΛ��lmųԬ����PbLW	�g���ndn��@�5���ٸ��� -4�]v���H+s� �j5�KX/L����y�z�HC�|UH ������8܍��^3�"/���m�B�@3��gN�S��P<��)u�%��n� �b��e�%�W���)/ﾎ�q�p�//���K���	��Ԉ�S��?�uT��� r=p	 e��}EN����ą�a��Q�-�Ω2���Fy��r�3�6ڇ5��м� �[n
��8�Ή��-=�\˵<�ufL;�a*^E�Զ���
�j�f�^���).Nݔ6��n�����Xm`��t4� ������-Y�I"u���п��`2"H:��'Aע�D�21���O��9�TtX�a��@�w0��h���|���a��T������F޽����A��E�L_��(�ϵ0km��5i��u#���]���~B6=�Th�>�P�!z�9Nki�� �����@ '����T��Ye;�!���T^�!ɓ�&��.���^&������\#���kN2հ�:�࿪�j)~�i�gVY�C�������@�@tq+N]tŉf����LO��}�X�M<.��$��5�9�;Q�>~VG�
D��.I�J�ɱ}L��B���z��hh�����T����ʭ��j|o*�u��5����i짃���Pb.�������+.Hř���^5��Ub	X��7@']�)u�p�_,��U���а���Dc�U�l��T\�lZ�Q�p��+'(;H��V�C��Ld!0��2�#���`�J*@��a���'T�������Xs`��tnNw�Y�P���V���$�f�P�b ���G�_kܚz�6P������@�׆N&�����((v�Q{ץ��9a=�fƲ��(,�fY"iϾ#8��)~�&�}D���,s���r'�<�&��V��/����.]����#b|K����|�f�Nʜp ��-_?�PY@�cRC(� dX��� ۋI������'� ���!�a�2����5��y�Hzb����=��`j�-������ڟ�뱸���r�ݔ9��(�W�"�!�֠����χ1l��9��R�!X��OUS��Twvө�AJ��G�>�-4����g[�/ ��^�I�fSӡ?�V�w=��-]8��|�6��}�Tɧ� I���_���H�ϟZ��T6sQ�f���@�>�*8��B�I&��:��Gd�Re�^�?��e��6]#/��Vx�8�g��hV)� v�E��=�{�VYW�a�J�)�Q��z����0����%��:u��BG?1�	�;�ցΎ�:��6>�]u�j�ň-��?��_�qxn��	�Ñw�<
����njư��d)\�Zݒ4c<Lk+�	����)��:�9" �t^1KpI��n�?h��#N�`�7������Z �&��ܗ� �)� ٭xoWqll�wd���txe���Y���@|���F'R =�@�������f���@Zģ�L�y8tI�Eյk�A�*9?��b1�|�y��$�^��4�؏=
Y	�y.��m;.�2J��$�%�^�==^�}:��5������͚jAG��(���W8S��#�N�/p�P�|��$�廞�Ċ�e�|�K�W�����e1r�Sݝ	3_�D�6�} 1�a�0`��ϱ�C��yx��a��=����j�B�?�[_<�u�J��k�b��0M��٪���;~����+��QS�С#����j)-MK��3w���ё}��	��V7�A�)�,++D+ԯ��o.��^�o�C)�*7��"������V�E���ͽ5��T��>��}ڤ2��W�"�YSk��xc�vHO~GD�El?[*�k��j��F)������C�O�>#e�ԟi�k������V�v���Y�yS�2���m�%�w���N낮WW��'lh���t�>������(w�&�7G�k���p���̞ܒ��x*��6��Ǵ$ݞ���,ᒆ�D����;�G����o��g,�M�3&�x&�ٱ���vXh���Qȍ-bt��?II�&Q�@2$k�#!�_�`������[��Q�s���_;��Mт���]�f�πYO]��
S��Y�d���)�e�ª+ŀ�,�`{\���j4�����
�m�,�� ��f��K?S���A�P|<DS��@B���q`�����O2,����ï��)Y�(�����?.�X�|�����_}���1Ōe*eh�yX��M|yW���>h�S����. 8x��%�p��w�Q��b��N��.��mȑ�Z��R)+�n32�)$�M ���ђ�ŞwRےUd�p�_��H4|�8��=�D!��`ά�� 16!���1?��Ae6$<y�9��(B�8��_��Ǟvc�_ö��%śT��e�-�"=��5Ǎ�r���=,�&���Z�y�s�%���|�)��sk��L6���`���e#��3_$���V����vr�NX����<�P	R�ݙ;{��g��Ah$�t�
C=�n��k�#N�t����C�~���#�k�P�
N��^���~XXN[��D��.��^|�6��&0k�2^\x��_���x�Z���C'35��-j�"~�*��->��*Mˋ1#�����f��ffN>tO��J^Qr�uyEmG,���Ζ���ݟމ���c^4>��X��g�v	��r(K�u\Q��5�ӓ��B��euR����6��q����UE����x#)�|G�U�īj��	Wdr��ʘ�4��ڕ��ƺn�ѷV��b�O�X�����>T�Y�0�8RV#��^2	Xw��+D�)�'iƘ-n�t�V�=��^���]0�7bϵXnݭ��eR=�|�Q'�N"�Ym�2�H#,[�H�����=o
��9VY���xޥ���mv�@����3�ds7��9���:+&G0A �Z��Q�vj������Bzbk��+i��I8ӕ��S�������*�́�ѓ�wx����ps����A��D�{k������$�X�O��B�(3���X��H����J�[���O<nE��.��EǺ��AC��3Y�g� ]�&,Іυ� T.�~k�I�#g��J1J2`HRK��)?e�O�'f�=.����J���1���0 ?�b�]�o|W�j�Z	�����1שL�h1L钯~���)±�U��H&�u4�M��J��gM����[��&⊓�X�d3Q�ra9%���n-���|���8�G"�����۲�ؼ;�mq�2�����FJ��| y�i�����B��'Wb��L���v��;��ſr�v��mD���^��~�g�ʯp�	��'x[=�������(��E|�D���iL>7�<X���x��(;�1.�fQ�W�F��o�F9���X�3V�E�QLx[���CD47�����{s�]F��a��[2;���ė�Gr+�ŏr�C,�ǃ�ǘ�* �L��e#�X��?F���p�#��T��/f�ɴgV�����=���F���֤fFQp����n�d���R�h_�lf�����jꃙ��D�Pr�p��ʪ�p'j��\I/�ڐ�%�*�q��[h�o=2fb�$`g��Z����Xշᖈ��M$�1j�W�m@�����ty��b�ra�jѫىp�n:0ӝ����Pb�1�9��?>����1ޭF��'I_�=ŋ�xwFc�|Ln|L=����>�C�U���͈��nv7���yǨ��S"6zO?���]�r/�:hֵ�c�%4�R�@�Rm�FQ�}J�%u��nG�}bu����������]B��g���~�5Z�� ��� � t�jb��@so6=�Dk�;�/a�`���W.���c��KSߚMB-K!�I�0�A倫tT�����f�CIH�q�B���4jZ|��f-�@��m���� �������u���%x��a���;�y���|.����{n�b�+��`�`(���_�-U
�)���vrP��7��P���N��i�J�i?7�WIN �SѣIh�^�E�X`����n�&>�xJ�Z��yC'��&�%"��ǝ*Lb�����0�.��6�X�e2*৚x�C"�F���b;;��3BQ�	uU��0�c��Y!,B\D]�ڑ�.؂7�!ytd1���{�>K�]b�M$��F�Ӏ�'��� l��f� �`J6}�uTFH�Yrg�H>Y��ّ��Qɜ#��2ʕS ¨��7>��q�>̮�ȳ���S�ԇ%&�I��1�p��}��L��B��t��e��痌K�if]�0r|��8~ټt�7�3�& �7\>?G���=xzN�Sg �ϝvMS_���w�:b+Y��gwf�Mbz��dpa[�����M��Z��b��l�Av����,��`�o R��lu#2�c�ȝ�(�Ӯ�%��q��ly
�+��z<��_f]�-D���Ϗ��O���|9��K_O�Z��C���&�����`��]��(ӗT�XɄ����I�T,D?ѐ������B���&~�>8��TRB�-���Ǧ7-��X��pi?)nl�,y���T�-CI�����Տe��ѷ����q����p��W�	�؄�~�]ؾ(v�@��N�ը�;*ي�=��Ϲɀ~; \�U���7R���=��I)���o6�Q�Pz��D*��=2PN!O��Ub%��Sz���Geh+&�%��D:��qX�W�`����/��hv$�I�"�����_#��d"`�������Y���c���6�?4o?��#�G���9�\��g�aR�,8�!�0������0@����Ns���=���4$���PL3C=L���mFk�SYB}��b(gz˲q�5�q�[
���N�q�=x���1
�A���<6��?�D��3w����Zߓ}�ϖi�D���-��p���:c1�c:��E�j�y������$`���m�	T0ͪ�q�Q����z��ޜ��d�	��w��/N��8MU�p�Lz~ +YHgoϔ�@�� $�ўQ[}a_�R�EC�O��{�SI�	u ��0���T�gg�K�[y��[�鰩����HwRqC@��"ϰ�G#�Ac���H�l�}8B�����|�(Hr��QD}�-7�7� ӗ�;�f�i��1�V3�~ur%m���Kw:+*u�	����>-���O7r401�+���,�u�.֓�p�T��BZ�H�X4�e1����|<��H'�f�e��H�hx�����/��YoS|� f�B����妤�Y?A����G}6W$��/1Hwh�����Dܩ� B��h���Jf�Aq�B��Q#���L5�3���E��ȸ�����g�.��S0��谹<��sU$>47�;(���q��	�=lJx���B�.� �����8�㢎���qo��H(o���D��M�)��h����x����A�]�_;��&��HH MW@��R����7�>��Ym7��d�s�[�a[���n�%�i5x9a��P�ƁH'� ���J���T�Z��L<��jS����Iq�Mד�C8�JǇ��JV��_�9��·^o}W�Եj��G�i	����N����Rp�^���������� u�>�*�ފL��LIP��G���� �����Ep���E�A{���iZ+I�$]3[��c�\�u�`N���L�������秡�n�ed`IB�:�
˲����`�#�����:D{�&�� A�!D�9uj�Zo���7���O��ve*7��< q٪�Ґ8�u�������[II8�<Ym�+FE�$��o,���B�b���Cw5�c%4C{0����e��Q�|�S�x�}�o��*w2�Aɒ��:��o9\�g��*6
,$I������+��--�V�˻㈵^�x�m����T�~mʫ�d���լ�ꄩթ�d-L���p��E�z�+������$?�}튶L�V�w��.�J�3E[��XE�nG��[J��u0n?;����!��;����j��4�}N5�.��zO����g�S5�nB�e��HC�*���Zy���>]cb'��U��n��kn�|yǵMMk���
T��c�>�#�jc]r����0ح���GW
v���^����s1{��Ņ��W��K�_~���z�^������iF[lU��ר�,U�+)��i�Q$G>��u�s���9�5���w���23+�U�Z�o(;��:��7j� �J��?q�!%��9=����٭}=*��i��/��|3[T^�N�8k�ĥ�E�҆F[4G
#��I���+G#G�˺&���4	w?�C��?lg�h��F5��ff\9�� (�}_���J�4��].W�e�'W�}n��k��� �����&?ߜ��BBP��w��X��9�N/AX.P���b*Ѱ$9A�`�?�u�[���r��C�<�Vw��*K�-GPE\毱�-o%A���	��ǁ�y� v�҈�a��h����&�;��<��� _�@~a)�Gפ�Y��G�kp���X�jd.�c��D�f�+��ZM��p*��d�����i���O��AC�r#x�?|��Jn���R�h��s�
��u��.�i���G+S�`������Q'�'��7Y0�"�Ⴞ
x[�eh_�
��6�y��>_H0�ά�n�S�%ɿgYw�Dz���9������G�l4+�ω���HF��82Н?DS��#��"�
0l��3���Ef1F��Jn>�;�i �y�a{*�7�������s)�S�x-i+Ҋ#���Ծ(@�r~<��T�:&�Kn�k��~/,�v$��0|N��Ŀ�)7�f�Ne'�b6v�����*�J���e��D/?l=75l��}G��}_yh�"۵��Y'�S��#x|o�o�זo�5�Y"� q�~���;_El�jdUl�@/U�>)��Ӽ/��p=~q��>id�P%!M��OQ�&�b��8F�m_���|�d�ϹT�*~����z��7��fVm���y}^�i���f^�I�I�!���zh���H���C�Q��H��l��\,���{/O�����f"�N����ы��:d�:r%��2j�lg��xʳ懊��4	�fWaor\�1�'�]�!Oܒ������H��Ix��]�d��p�o����p_'�dc��hW촲0�$�c�/!`I��5u�ɋ��l��xТ|��@9���r"ۃ���D��������=xW�o3��.�z�NWX��T���
����F���?�v��A�T�0������E(i�$T�qiB[�S���A����AX�}ђ=��w4�����ҷ �[��	�;7C���-9b�"go[*˰a��L
���~��T2��q�}��#`9ǡ?U��UΔ<D�@�EZ����@��K#Iad3R'ޚ�ZR�fZ�~��K���>	�]X"�귑V[���x��wmLS7�Ay�
?��
�r߃۩$�	�%��^�5U F���Y,"���6Yd~3���J�/�ȧ���6��#�<pe6��B���W/Kv�o~�����S�I����,|.Ībj�jv02\P-S?u�)�F��՝�e<�.e􀹫��>1��{*��	��=r����k���ê�r�7ҚȎ��%;�ųg
�����ϵ9n���</z?�0���8pY��ӏ@#�������k���UW�Sfo{�����:t�|
��-+��9��m���8���éˉkB�����Ȼ�ߤv4s8��&<ˍ��` �<b����v���Vp�i8�>��\�'��	����XU��nY��i)[��A��هZG����.�e�j�d�AݶO;.� YJ]}�TN�G����Nos3bd�	Z��K>�
���El�����=���J:e�� ��L��N���B�B1	���&�C��u���ɬ+-�z<��_���#�j���̍p����zkG��dB�K,5C7M��!�x7zT�)_g�Ul{�ǚrb�q� �I�)"m�*�ݦ�����dg�H`m��ËN��/.3�u���	#@q�7��2'�g4��aCR W#�KV�
��A���W��h}�Ħp�jÃ°��5\1G���f�> �1eaYۂr�O_�2a���:��ՀKoROPv.cS�O����_�H?0��64�e�w)�����i׉(m��p/�`Qk�Y�z���T�-�0�SL��z��y���ώ2#z.X]v݉Uz?XH��Mvg�𷛦:�O�i�u�b��7���'�Xf)k����"���;8��͌�Ĩ��z��w�T�����#�����;��t��E���B߀-]��ĀRwǣ�b{%�����ЫTǨ|��	����hN�)v�:�f���k�(�t��O;�/�[k=����;?0U��T�4%�^mXcG>�s�L*��S���ȗA��5�o\͋Mv���k�1�R���(���t�E�ؼD�Fi��n/��=jk���d���;���䚛��>?���!L�@Z�>�,��@��;1lc�&\}��d�tړ���WA
�"B�3�f1b�۩&��� �k[ѳ@{��?���O�'�em=�EL�LH}ݯ��NwSQl� \��O�"� ,"�������S�g�|�P�3�~� ŏj������3b`��,��y�5R�갻��j���b��VI��G?'�&YBi��ai�r4"�!Z4Zy�|��c[���o���fJ�y>�{~T�>nA
��dkI=)��D�x�y�SXs�YZɳ�g�4]ݺ}�\��Kd�x�E.!ͭc��Ζ&�Q写���}i"�/�ħE���Kxi�=��5Dj��M��]�.�x�����/�W���$2W/��V�~N*�a����H��!B*�uC�)ƪ�)M-iT{f��7�7�sNh�l�	�֐�Ǧ��T�����|������q�@j��0�ش"�X���O����A�%h��q��P@�y��@����m�� �H��$o	G���&&��Û�<j�h��0d�3G�C�}��K�vތ�ϒ�'�� ��R!e�6S���)�gU�X�E	 U�v��՛��f
R�����; �wX��1�/����~�A2Rk���X��d�S��R����$eyLMH=P�4� �E�]�b(ώTr��%ڲ��8 ��3 �<�,�)�N�b��$5��8 ����z+���9�4n2����1��,�_V?Z�o騠-S�fWP�J���j�q9(��3d`=l[�y�n 1֩����&��v_�I��@kY~�J���K�P{��l�{cc����æ��}e�S9?͟sh����Db�B�pF�Z��W��1���MA��@��+ܽ�3(�ؘH�t����y�M�ݛ!�pJnL"|���@��'֨G�Ar��ew��,��}��a/̅�#<�2���d����n���
]oл�(�i�r�E��=T �Q�n#�]�R�K[�z���{��&,%F�����)��l�L!�/�7��S�=�"���>��K�woO����f=�Sz:������6�l�����j�4w�R+*� �Ml<��dh�+���;��P��D�7ک�Ͽ�r��:)��V�dq�������jsF��+/?�+Kj�,x�6\��Э?h��2��Xמ���VWC��(�&n4|�M�N��q�����I*�D_�����W�N�~솣����9!��VK�jU��V�e�9��wa��J඲՝����MRGo���y����;��zЛa��p"*\OMF���r���5�m��_S�� z���֓Z��d�=Τ�֌\�ݦI��]� �f���zKT�8�r��'�oҎ�W}+N�X������&�7�\�r�9!
�Y�N`�������+7���">�)��=iG�;v���V�I���V�>�Z���K���i�:�Z�'��܈ad=��:4�J�\�Ce0y#�;	�:(m�D��Pq2t?63'E*̀
�"Н$��@b�TB���[r�}"kR��kR��H��S1�#E]��UEy��_�*�
C��}�ޗo��nS;Ջ'����|T���F��!ݸ[T�_0�E��'!/���N�S�#���Be�2��%���D/�r;QF��XcF���f������Fwv�]ҧ��רl��V��AG�js��j+���N@a���N�ObFr����sV�Cin����u<vʱG/�|���e	����kQ����
e)�t���f{F��F��Bm�JN����q�X<BѮ2l�{6?�(�Vz�}	#�v{��f�c����H�^j��e�N�v
�AR�&�"%�Mj:�0��,�e��)}���gn�:#8�s�liP� ��� EX�۱���|�sm�(v�UjLW;�m���rvG�\�������ɂlf: ��n�����WUVpR����������vX��!2t�~jr`CHX���h�w���ʕ���@��*��9���>�Q�O3E��c�����8&�c)����
���6��}��.#��'���:<2̳`6%r}�� �I��#W�w���W���E�'t�8��7�Y�_+�'o�D�:st�t�g�T���d[hx����s=M(��ߤ�D�|�j�!C��!�fjA�Q��r�M��?���+����b�?��׎�m��%L�;�Eh����ݧo;�=�J[ ��w�m9�d[q��DYW�,R�H?1���X�4qO���dhMOw0�����0����ڒNT~٢��@Y���Ɠ��}P�1BA�_�����L?̓	��'ݔ��/�zZ�4�y�HPA����!Y��WQ�꧓H"n��Z��v��)Id~���-�Thd.����Ky�[Z)KV�R�c|k�����ak�ΓmA��������$t����m+j��X�'4�����H��V�1�X����o��Z�e���on;�?6��]��D��-�L���Ҍ��3�dR	���|IwDD��y�
�D�����pщ+�������7A���+>���`��e'�L!��m_�f?���0�G�����m��Rp�Z�������$�e]>͓fz��l+C>�*R�7�V��Y]��A��93+�<�)�tyZ�w�K�Sn)0����{�����@tV=��L4��RP��gc�b/!�?z<�P��h�w��] 3xʲ�S�*72T�
[l��l��ˉ�hd.G����sd
�N�w[(���k�*#�@s�� �����Y(j��6�131�yU8)�Va�~��.AVޮ�����Hhۛ �b�A�@�{��cӡ�����t9�D��?�3�;�����|��[�~H��[���À�)��t�ǥ&�#��&z�����,j�,�GS>a�7|�k����}��,t���(e��y�~|H���124�T��ik��� ��[�Bd�<�r&UE�g���l9M�J%�J�l[O���ZV�ǡ���T��%���Ͻ�cF�X�8�J3�_07#�|e~3\����F�s�?"�},��Y��s3Z)eW��]���C�z9ˎ/���HM(�J.���5/:�o�'�@"�&#�夗��7s������5	��&z�n�㉍<���_@L�}���K��y� �(�d]�ֶz{B���S;�&_ņ�ydV�������@���#X�����U4Lٜ��S�Y��fΚ�� ��[:���$-�|�����[�l&}�	����&�� �f�,��z �I��j���z�ݞjL.�b�.$x1�1d�Ikrl���r��aaF��x��%Q7��师��5o�+�irb~ �h��zDؘ<t,�C�"�5�M�v�D�s������&�;T��f=�4(z���D�cӼ�\�������p~��G0v$�����i?4��gg�)C�1Qqi)q�eB4�2�yQ�[bR�6F(Q��om��r��U[��$ >�~����"N���Ǝ���JҪ��JO4U�r�9�̩��F��8r ������ʘ�9�J6<)(����ŉ=}�xA7Vt���6)�NQj-��7�&���v��7ӏ$�}�inYGs�����v@��a��Ǩe���Җl�g����H<� +Y��wl�à�yIO���U��~h3Ӵ��8}�R�.�>g��5Y)�d��d鬵�2FL$ol���E����/"V����qXJ���[���d�͵�GM}�l\s?�r��S'��h��q��l8`���Β[��k����;:�)S�'X��ۋ��I��G�zPcgT��8�H��o@�m����>�vm?63�oD9� n�BHu�</ ؂�(�
^~�"m�#�.t�d��k|�ϒ��3u��0ب�D��̙E��)t�6���Tv��Ε<ڗX��:����>,S�o'j�������I����H|�'Ng/�A�* ���j�a1�2�.cr��8��R��$���r�!`Q�`Q��֚����ѡ��B�k8ƿ�/8�-E����ܷ�Y��ѱ9�5��
�dZ䭪s���_�\ٻXl��޷h�ٶ13)��5W{�|f���3p�PO+^�{������G"�_��CD�Wt�#��}�A��<G�P��L�qw��e��2�k�z�l�%03'�K��Y�����!G��.��ixD/�ɡ�lº��J��Y��iM���N�h��5lh#�� C#VR����X�R�>��lG���Ѡ����I,tL{��h���<g�KWB.L^F���n��������L�'?�=����+<��VD9�5C�2{K�	�$��ߥ5β@��M"�$-���V��**��d9t�?f��&p�O��a[D09��!�]������0G��c�
��oI��U������mG�� %�+2ʲ�q��fy�Q�"V�|�����(J�xI{<��Z�}L7�r$������H���X���
f	|l'캲S}�4����1�^�H�X���C5~���MG@XPڵa�=���Z�v��������"�\����P��V��6
�@���;��M
Bw��<���)���w�X����o�O{�8xшR����"��b�]h��p�r�Ӏ��r��)���Ǝ��m�Y|��#OO�Ѿr<��t�F�EeT��s��h��(9X�d��zM���5�
!~I@�a���:��hin���sG���>��'b�H9ȵ�(mN��@**^��,Q�@O�' �6��Zb�UJ�[���<�9绸��W�@��1��+��9գqR�9�s3��+�b���F�W}Tϒ����Rf�-��V�+�!���W����l/�%2���r��Hr���?�.��c����kN�j�i"��M�4� H�#�9@i&��]��⑋ �֪�,���������,`f��c K�Ӥ_��1�EdKℂ�4�t;濧�>\�<Q噘��յ��at�gc�X:�S��D�'h��i�ՠ�Ћ��i��?3�|��$v�B
>$u��� Ў����^L�)�&��/�u�GJ	���Zv6<�וJ�0��	���)���X�Zm��״�ru{�y(��nR��cU�|VxIx��+�L7�mt/����d�ض���>����'��b��lx#C�ȹ�{-c��0������|���̛�37��ߧv	*5e�M���o��s|�����u�R�����A��0hzx��?Bӹ��~q���c/�f�֪9�S�ʾ'p�A�#�����D)���S�f>%�[�#V��5v�� �ܿ�b���Q���J�`l��]]��L�'�B��_��*X]+�k9��Gf7[uM���=HZ�uD��$��l�_ti-��<��%FP���'�* c}<s�Q=@%�f:��E������ �CB�05i�6�[:x�l�\P=]('�ґ)[�������M�����G/����(KŞ��x���`��d֘ŉ{~�ADT��t�yX��Lm�CD%f`]3�xgf���i��>ŀ����e8��=0�{	0�vY� g��FY�.4_��2�kw�~7�O�q�q�=w�)'�s�>��K���j99̙MS��@4�q#�+��F��)6* �u�G۳�d��py�>�����%�R����@���Fxˑ�k��l����"�9]��t�˛����O	X�u�� �M�{wiqܼ�������ʡ�N�@��`����QI�=��}��d�#��\��%=�u˺`j�,�����]V`�	rRv�
ղƖk����hG}��(D['�戏�c<�h�����r��w!Ƈ�6q�q��}��X�Ql�j���X�����wU�-+meQ�	Ӊ���ʕH�W���n*�I�3�6g=$j��m�<��}��<��4� ��H�c+XZ\V=f:{ܧ~�zoxM��3uZ<��F.ƻ��'޴�1~�Zz���+˻9��II�̻�
�b~v��5l����C�6w�0�!�ni��O�feFֺoC���6���� N�������[�15\��$��1�uj7P�A��6�oX,�a��5�3�X���T���yN@�-D�Ǩ:��A[!ZyIs��j�#@k��Q305��|�[��\��kQx��Z�(�ܧ��)B�}����jP�Yb§N��Aښ��[D:�0љWE�m�u2c5L��ȘU��֗��y��*Z�˛]��>ʆ�k�J�Pb�}��&��ܛ�`U�eLm�� N#�gD�\'B�N�P��D�>M��.<�Έ�b�E_�b�,0�n ��:Ş��'�5a����*�|Z�!_��>g9�R��x�׆ü�w6x�P��$����Nٹ�α����oSzx�b�aߎ�Oп�#9���s�L�V�1�}�v�N��\뤈S�]�Gsnj~���Q�v�_45p�����չ�u�C�cb>�=p	� ��A}#ڝZ˒����0����w��g���T.�BY6�}l����=`���ZnM�~��C��Ȧ���� Щsx�9���U���#k���?��Ҙ�7�ϛ'��G5{�� 9���(ɝ��8>�H�I���[c�q:G�'�E��[`ێ��Ǜ@{(�.�	.����[#�+��$�]�ų�q�%�'c�d�k�$@�c�	g��DT���,?I�gl��Ҿ]�K*mh�@����(������4���\�JR�d�x�b�/�q �5�~�4��I��V*��Z�!zK�7�a��+�!_@��4�x
O�/�����ʓ$	h��	�ydY�]��x[�v J�0�-�3�իIe8���g	+�]G�`��F��l���YM�r"��J7�՝fԜ��������W��v�'���u#l����F���H�1�SW#��,[|N���X�#c�Nb�+��HX�H`}*|C7-t�]P{�R��-����0#b��l�ST�ZCޖX�Y� �V%`�����j8��,�0�O&u���R�`���H4�����*b��,�Q�OO��A��z[�2�KtioT��(F_���6G�N�Ms��{e#4|�G�
�xHagy[=<y־����}��q����6�5�25l�Yqu2���W%�ҭ��{����_���Z�G_�8��}��(ɫLɥ�W� �TY��K"����Dh����0k9O�������!�SЇI��B���S���h$'9X=��L���&�g������{�#"�{Z?�Pj0�Xf�v V$���ts�%�q���T8��4n����l�eU�r�6#lN�m�L�A�S�$b���wF��9�U�l!��k�4@1*�d�;Oۯř�Kʮ*xkB��������&�ʼ"$%o�"m���6,il�e��'�"��i>.�<MN��:{�@���ב3����U�>�ϱ�����R�)e����}�j[��'P��wN�I�'F/��+�$�O��`I�h�an��6�IͻTe�L]����1BjW,��9wc�u)}�w����p�x�T�O&;p�퍽�,o�R�8���;�g�U���`�|(�9\|A���2H^b���+�c�]��z��1��j��m�T\Uhk�7��>�ڻx̺Qz�LBWJs��%/)A�*�:yj FO��T�P�tH"f2x, L��Y��:�(Q�	��?�W�-֧>�1�)88��1�'�����d^U�2+�4�����.iܒ� @�.�������/Xs��D��3*���V]f��S��)�qw�e���S��0W��A�\����=���<�*=�e��2nF�)��b��"�1�gH��-����R�E[�/�n�#�RBja����������YT��cm�2�i��Y'0��K��ثO��3�ް�����N���7�@����j.NG���bl��{'�K�UeD���')��3W���ے�~�NZ����n��i��~^uG�["+ �E��p�L�)�r_8^�{!S6�>-x�~t��qs�er���1Nt�m9K�(嚵I�m$�-����4GUܴkiF��z ���r���C]���yTW����9`t��e����y/��u:�d)��c"�uv^��X�<�T�,��W�ފ���li0_��|u�u�����O1 H~��J� U��=*~���J�o�
:�ᮊ��sN��������|�9�ݯ��7J?w&(�bm���-���y��"����Qw����=��LL�x�R��2g��,�d`�$	X��>��L��=�SB�5�����VQ��G9U�`�ߺS����0��j`��Pr��%�$ZA�e�F�,�I�(:d�  y�����/D�7�=�Z=��S��Cu�;��5��夙J3��~r���	ZJ�Q�z�Y.h�������^��φ|��9tC���d�>z?�ua=�%�