��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�!��
��%Y l�׾�m�F��������2�p��X^h��@��[iKd���3sΆ�@���e)r�atVƿ��ߨ��d�_5����J�&z�<�ܮU�eM�%��fG���z��k��X�D�]
�*�M�������q0JE�JߒH^7�8��=��l���@�@�^�+5�;�=�����M�1)�o.�5Y��9wgW>RŹv���bp�\�A"
���z'E�T_���9���*��O�N`T�(Z���y�dw1>ׇ�����x/���z��J�s" �*~
6�g���h��g�xH�>�^_T8��0��o����lz�b87�_�9��(�= ��_E�t&6EUX��cB䏱t��ԓ%y;gy�%����FH� �HwQ����y8�9�ʩ�瞺Wk�&V؎�#τ���q=�!?�Dc�ИI7��d5���i	�2��¼�s��퉶N �.t� �n<V
�*�niǛ"�ڀЄ��y�T� ׎�U��mb����?��T���$��ňE���,t4$A�@V׵�wY��`rP5�b��x�D����!��ɱ���y�k������gJ<��Ѥ�XA�jJ��R��s5"�����j��.�U�b��:�{Bhv�m0!���;�.��6LFe�;Z�v-;{�W���6}^$K�
��E=L�5��P�WgL��5͌<�+C�b�\�%�G��#K%���E(�*/c�A�_0y�_���x_L��*��8�����P��cJ;y��4��&��ykh)����\��f�;�ָJmp���J��CY#�Ȣ�M� G����#�{#��yzFU$��G4�%�����z�x�A*�6��m��+�z	�A�n)�����烉����Y�t�<d>Y�L6�L�!ZF�t�c��̍ Ԙ���"R�Xw\��++���,-��
��{��`~���Ub;��?���.`��Yl�_�4����F��Uvͦ� ��u�m\�/�B�U�Hs1�7/�J��gFg5s���Fp��Ӥ32�Wr���o]����[!�{�my7>?>[E�3��p/1�=���E����ڋ �����g�ʐ�2�"�sds��^lO&^Ќ��^�`z®z�%�O����Ȩk��ц�Gw�R�Y1I8U^��xG�����s=z���u�.,_0ܖ�L&s\~)�<�gDf� �\����eBѯ(=�7��������=�h�HN�>���Ȝ`៏#\��h�!������v�ʣ�����	�:�R}��0�@���-]Upeq���7���s�y����TWn���+�<�c��Y�}n��U�9F(�/ص`%̞-�l�Kvf��i��� 4��-{�EB-�4�μ�>cJ��[L�0��=��2���Ú���L8�����{�X'��(�*�`���i][,�NP�ş(%��\_����(�������
��,���նv�JΥ'�+�k0ʧQ�U��-N�n��WQ��x�@A�Z	
���d��T�룍�p6b���e �YGq16Zagt:�`�D
n�+QhZ���π�#�!�dUCz%�ɅG'_�$(��
[�<d%��n��N۷f���>�����*F�c�o|�"?@5b�X�J;s�g^�땅#A��֋��k`�H���tm(=u-���(r	�����3�ƃ� �Lv�o|��1��(���$��'�y!��ڧ���� %C��L�A�1I��,�� of����j�� �����esG^�.�*�0�0$�@zs�m,��$�K}"#��+4%�*%!åӻ�1�{�j��=o"�X���}HV]	z�U+�ˏ�Ϩ�v�A5_y�D�ƶE��p��S�Mx'&�q�:��X� ��-�Tg�<7�3K���"�!my��i`p�G�Th� �J����	�%�qH��`�dO��i�Q\�2���������U,g�-�C$M%�ҹa2Ƈ�����T�g�F#����]���'e�{a3��6���O������.U��e��I=1J ��W!u$Ӊ|�@�X��%xu=M,����0hv�Z���A�TH�dVVİ��\�jc]��Y�������rW��?�=���������䴃����e
��XwA` /#ˊ��Es�?�D���3�("�o;�r�t��'�2�A�),@��b'5���w8��gR*m��7�gCP�
�8������C�)zF��;%f���O[5�*��}x�sQ��:�g���!eN���4#�f�`�}��31O�`I%=�� �Ӱ�zc\la���H��>�㖨5��˹��/�B�g_�2 "�iMKtI�pTU@�
��$��j�'��j��;6����`� �U�=�C��^���������)�Tp!\xhY�~�y�Pdj�?Ձ��ɒ��{��.��*���!��j�F����D(��:A�P�1z�N�.=ݸ���@��*�v��S�P=�J���u���]cWe�ەLy�����Y��Z�I� �/����XA�H�{���������do �@w�[P����(Љn����G�����ʦ�9Y��������q�p�z0��z�f@��+3�2�G���Rϕ��a�\o�2jo��`��6W�l/�CK��X��?��O�굋�Hփ֬4���y��̈́� �y�o�K��>��F�M�������z~z�}��d�J��w��r;��h��]�Ve�a:i�.�J��2:�M���4�hU�BCnb��=�9}�>�N�R�&EN��	!��ъ~�SRgG�q_�z�+���C��w��a0�8 G}�q�!o�����ߖ�6y��� 6�,����X �e%��,{^���K���Բ�i�ӊ%?G[M ��������ɀ���~,3u7MS�Q ��+�Z,��e8�(k-Y�)���U7+��Jh���+��Ty���$��T9?���1w�
���d��������/���_F��l���W.u��K�hR�rG�Ž����wv�ۏ��؋��I�ЮrU�3w�H5��� ����Z�ώܳ�> a�3��6��0a�%D\萚���
��~���^9������%'a`�	>:ʏ�p���8Iܹf�yt#\��g��P�ã��b����f��H.�����g�Z��-��B�\�`��q�6fb���:�|���6���������'���	��I
jxI��^c�۝S��e��K�g4�Ŵ&�{DZ���\���Q��/f�>�|ߋuꩨ�,>�,Ք��=LR"��O��T#:��I=�Z��lM�E<D�Go<PRE%����L(LC��[��X%0:i3o�!�@It�(K��b��������S<P0R��7�큘�ma�f������;U�ۋ�:oOZ�,_-�����y8����8�ꛖ��'9:{g�0����	��&�)&��鵌�s#L/?�#ֶg �����zm����,r�	G�@iaA��1��#����r)k�h���p՜�,��т�tF7����w-�އh7�a���S��a�M�ʕ4���3��d$Q������zk���Ң~���ևr߭�vɴ)a�ˈ*6��&��g�G:_��	Z�:04���w��"�?���N�>:��O����,馺|׭�����a���>ᩓ���-Cv�#�n�A,F?��U�F��ؒVO�)�P�딃}5%J�
v �+q��)���s��et�@��4d��F�#d.�\^��{>�͎"D`�ټ��|�@�
E�D��#*|�(ԡ˶R�"�5���3�Dx�\i�g�Yg���`$Q�ުOv��ӏ���U�nE�y�FE'��Q�8� 魟��$ RTp�	����H�n�M�|+N�@t���e�cC3r�S@���y�R���*�VjY"�������V�P>]nt�d�e_L4vռ<��aCy�>����xA�>���5��!�.в�±�?��( �p��8
�d-�TXHG�,�ż�携���9����kz9J�Q�	b�f�~��/��dr�փ������Q�4�$��H*՟��.�c�b��F�� �혙(�"�^nΊ`�u,���p��v�2�R1�je��;�O%t�/!����'��[�Ih  ��VU�.�������4�PZ`+XI`��F��pu&<��j���\7�F�y	�>H
=���A��)�ʞ�޾T����D�no�����7�������܇܏ �%!Jf�Ҩ/�-���7i��m��>��x-���N��x��}����X�3�j�vz����.���x���8�}�:��Z�f�ܵJP��
`��^�3��W�{d^+�s�&xZ��:Ĺ���(zI9!;K�ʻ{~oW+�ޢFU��z�67�:��&_���ESta�Y֏(��}���R"�\��~��#�Vi�*q�B�i�^�i0E��m���I��j��T4�t.^D�ߠy��54��1R�03�@^��HW�΀�H��N�(�56m����UfT�_�hR�hq��(�w͚�8���(�K�u9���SB}��
��31'`��\����'�Xw�"��S�ݣ6�2���&�x����$�=脑]6�
8�;�"���+h`W��'�m7!����� ��g�E�$]	����[�m���m����zPܓ�������I��c���bYL�(�nP8 �M�NO�� �������{6)0HI��RU����b���E�84q��.��Cd�W�ʇ^��>Yn��DD��_#=.�끈�`HV�8��(��I����D\�xEZ�l�/��?�J�|��L��8kMK2�ID�^���[�o�J�UI�r�E�Y��a��)��-a�	%�L;k:��Q��E\H��y�,��E-7�?�`Kd�͜�.�"ਔ�3���E��G�����S.� ����P��W��Ug ,�h/&F�
�+����'��D��D��g�A+�W���@=�Ƭ��*�1c��	�[ֺ�L�󔐓\U�·�4ދ�k�*�d��xk3�{I�d���|����R�?�5��!��vw�)Lx,�n*� �Ch�^�s{!*�;E�˗0�W��b���0�?���[|���+ZȽ������j Rqa��Q�E�,z�p�{Yާ~-��H���0h�'CˏU�2Wjl�r8�����"a��ّ�Z�.^��%���H��k;m���[kG��_u�^����l-9���l:csb�S|�(��I�J���<�x�9�TEIt�
&)f��)V��zP]ed������D���r&&�}�f�����3���SZ�%���J�zZ����4�B1`����d���V.B�!Js���#"C_%aن�=0�}l������6$��������ZF���_f�Y��Z�K͠�����U�2�[�>B2�}|�N�3�0��Ŧ��G��>|N�v�!�F��S?
�q��Dqڡ+�Y]�4d���J}9��p������lx��k��6y�c��?X�ݔ�HVe�Ԛ�c���.?�2j���2�թ�x�޹Uy��f�x����ֳ����p�����j�a2�ư�R���>$ʅ�k�a����������~���z!e�w康�OWE��sOp�i>Ug�A- (R��|���g٘�u�w�8�!$�u$I�H/�"�aI�f���G�]�8O�}��I�a�C.�Fp&N��JSe���$NPR��֌x��/��)�{�����`^R9ƉƪV�)ǰ�`e�k$��]o{\��&��2w��;#tԘ�p�淙dݨ���c��&#��|�(�S����� �JS�����%`�r#�|��X�O��9���
�X~?���810�i�S��m�xE��wۤ�A��Z-��%�a�Ǵ�.&mu~$�]l㿥��s���}��H�����ە!�Մ�a���p��ꬆ��z�qA"r�Q�~����D����߀�;� ��͢�r��.̹}Z�����|���3�i��ܰ�Nɘ����"�ȵ��|J� ���@!�����4wR����	 ���Q�
<�O�܋;�3l��+���d�p�*s�R��V���}%�ʄ����/G���:<�lt8��6m1��D WA����$�x�rL�Y�=RS�b�L�}�jy}ՍP��8n.]Zg�e\���Q*(�>���!`�8H�՛<��ο������b|����B�â��5�K"HP�k���&L�izp
&��9
�Q����9��t�db��ވ	]��nO|�`nH�ri[���wN�S����ۅn�2I��$u"XJ	 B��.yO�m�6��c���K��w0|��ӾRox�7��W��,�Ke�*������û�z��m���`�� -���Q�b�CK��@hP=��f*���_�S5 $SO���R���XG�N�D�
U��>�8(�"�zhSCi���sHD�NBv�j&8�<�b��5��Z�7��}]5D�qb<�?�Q�C'��v���]颧Ӟ��E��#{C"�N��f�ML::���Z������S��.S\2VػV�;��LK�ư	D�4?,�g�A�M7��j�nHUL���E�����g�]	�.� �R�i�Gs�4��:���P����}:��ϳ�Z��r���ML�Qr<{W�SrR5��MiOn����E��z�*FB�����:5f�,G�������b;�&�6�Ĵ,8���T��4�ȳ�ܴ����)��6���5�W�{*G%�I2_ ���LT�!�t��[��0�0Y��ly�J"W��/S4,�42k�*~?�7V�i?]	 nu͛� 'C2~�;4��9�#�dd��]������nl�*���i���}Q��a=U/CX۪����k���~�Ҟ���o�:~����+:/"�pq�~$Q]�Cײ"� [�n�=����l�҉jaCEJhF�ᛧ=d�u/�9����/��vw�E
����ڴ��X#ͧ���_��MuJ��-�1F���	2�E���w���
*VF���T5�K+�s�o�s���"m"�}dmQ`b��gS�(����^�L���bp.���pӱZ�%�?�NN�g|"�R����C`�~o�ō�åX5Ȣ�v��u�<����W(.��S���Pܜ�[����<LЦn��yzk/w����*.��!>���)�
�"� "۟�.@؇l��u�ejc3ӑ%���\Yd�.<_���!��4�kaI�G��
,$n�uO����-���
*���b�\��1r�k�oL!cghQ���9`�p.��A�aDh%��.�N��g�g.iu:8���\�#A�÷	|%���9>��jD�-i����]Oz�4w̐��,IY�����l�뗖ںԑ�����nE7<���6K2DNh��Z�j�����3@�sL#9�b@OY�V	�H�|��Zg��Q 2�1��"+ /�-g����*�CP�a�m#���Ъ AS�O�s� ��j�$�_!`lF[wfCq2�~\12^G���:��U�,l[���D�+S�",I��?���tfH���H�-�!Ú�Z�Ҍ���'横k�n��u�8�lp{[o�T�|-���.�(��-���d\�7+��e eR�������bʌ���8c�@s�<w���:�T��>�ۚ��rJ�'�Կ�+*��H�ď2g��#�$qPۮ-��&I�%7���\ ���u�`�\���[ڛm����%�k�Z87.�	�-��)/���db@aN���R�ly�iI�*k��jR���#��o�J���Yl�3Y79�І�<�WB�P��yd?--se	Y�܇�5Ϋ)��	]/?�1wG_�*v�'��P'�dp>�7Ć�$;~��'H���DU���1i�n�9�E�w��R,��qqU����$y�AD��A��V��^W+�8��#뿣9�BX\�����Ǥ����X�ԅ�?ҫp-�RO���J0���]\5��?Fug���BST����Żw��A@T��e�<Bzt��;o{��Wz|߂�]��rLR��0 'ڒ8�9W�
��R�P���8>��>P��p����/��/�E1�b�	B����B�f��P[89���p�I��Q1�-8B���*�D�6ןE�-O̝es�t�r����TU��bj�!�d.�4W�7대�����,�$�k6}:�nㆼ(L�G�R)P��N��]�K���9N\#6go��s;���f]T�[+wz�ڸ'5�U|��Cбc�dBt�J��Z��hrÒ��Ui��5���K_�cj�s����i����!��Ry1eC�P���ҹ_n4-BzR�ar	�ф{�~�{oE�OD�ty_I�H ��$c'*rV�"�+$�P�$���QE��t����2�f᪙�
$�	!p�D$%o̓v��{�9w����viO�]�@�Ji�������C���,P��OQ�0�/@HNF� ]�݊��:'6C\��<�"�;�Xv$�Ʌ����Z3<u��#�x�a�UT*��'��kH<�G�Uϴ�����}j����lKn��P��!5f��@8ْ��O~�[J���.Sz���zF�%r�[��;k�]�9vm�Rt��r���3h���3f˯أZ�ܰ��EPw��M�'��'M��,�f��XR�VM���V�+
;��8C;7�FX=yZ�xFe�,���[�Z���%QW�Hh�*I����z!?��� 3�����J�^�
��l�u3��:�|�&�-�����M�`rtl{�{u޸�D���K5f�r���X��W�7��ڕ,)�������]`ʭc{"�6V��;G�B`�x����!t|X����%A��D��O*�0�S��o��&(!z]��JǇ�`�l�*����k�tw�s�Kk�Q�"�$ze����~5l��g	�)B�t�M��n���I�8H��Ӯ}\Z�7�R �2�]xZ[�z�(�����uG1�<ؘ�qhT"�t򜪶&!zjS
�}{�7�Hfv{��|�&m�>e1��;c���޺� �A����B�<���vo�� '��@C��4#l��	ض*��}k�ئs����`��Jƞ���\�����K��G|e~"d;�&��P�� �۰z-�W�"�}��k4����U���������_��.vDe���E�MT�Un�b���-^9��0����?�ZF���r��(L��a�@�$����K\c��{",rǳ*~\z�6w���%?C�.4�&�`���!!���������\5\RZ�C;�՜^ �:zv��r"`����uG��t��Nl�����c	�9��������}[��8a�Mg�ю8ο�����t���
g�(#�dK�5m��U��nޮ�e Y�R�
�-I��v�w��r�݋yL���w�ŀ�l_V.�׽���pt��!w�}{������=����I�G�<n��R>� �.����I@ܭ�:�
�ý��֨��
�C�$���<�D<��y��F~��s=n0�P�hp�Lz�3�n�o��%2�B5`��YN9��6��yux�V�
�p��"�E�;�T[D���*e��#��P�\D�����"S��)[WMǹ2���/Q�>�N���aL+�����j�X]UT4�}�3q"�� ���H�*ؑ䟔�ɽ�F�b!ەTH�1�����󺨉�R4�F9���N0|���&��v�*�M����a9��	t'�	=�
�@����5@C�� kz�߄3>".�
c6�A�@DLq3���D�����Z	���Q[���	>B?����fL]9B���Őqwk�W���{��`|�mN�@��/�z`�J6B��������fAL�����<3��,z%R���E#Ҹ'�Y�8�p��C_l K��I���r^��k�9�W+���o����/tɅ�Ĳ|��5��[)J�cC@�Q��tU0�d�2X��Ǎ5V"���=�&���Ϧ/rI�U��m�_�h��I�W0�� `>IDqNW:j�Իy;|Ke?$������7WA�(h́�J�7��o��*b���0G�(�e��Wp�z�����I�V���k�]@��_::C,�~�zP��^1��4�{������adcpd7t1��d�	<���hW�B���%Z�t	�������M����pl�������Ow��Z��f�J�n�=�ߠmV��E�����z*�'S��ṗ�_	�*r����G�2cކ-$�:��*%���i�m�L4����ʉ�W%�~�ϊw���{��Lh����U�-��L<��:����k�H��.�8���0��D���qɺUԋK�h�>h�<Mɛ��R7��._!N�`݈K�'�޿�4*�e���K��\�密(��e	�xƼiK9�������0|�ܗ��D����H�"��(}G��xCq6�F����I7m�|'� 8@��t:���S�o����x�9�X�3{)��j_�"�M��Ds�h�Pm�(��I�P������3����:9F������i�SRl�Nٗ�JɊ��X��v:�{�Gy��Y}��s�e27��Pn�aɈ�b*�/�/�F�Ћ�F2���KJ�
`�?|N��m�f-���� x�?M	����Ke�@�a�-׿@5������W�Z�_�77�H�����T�7O��d�e�־�|7�A�C��qp	�Y�]mnNe����=5|��,aS8�R����:���[L?��U����AK�pQ���Yk17S�"]�c�:s!ru�O�kX���x�pcW����ཁ����d�Ԟ��������6�'truC,�\v7�*��u:ە~q��M�����l���4�|�Ե�O�)�M|�]����?H,I���k�ҷ"=��?�N
^�گ$��W��ঢ়�د����LX��0μ��'/���o{.���"��aj@��3�����T��Ql3��Y[�E#��E�֗�Źc���R֥:�Kf�)��rрI!i8��e�#��y 38H�h�J|���;��G]�\]�-n�V�Ω:͝M^E
��������J�r�6�����iMO��#J�W��m��4hǓ �u�S���1B��4v
�r�ű2�"�<�A�;�֤Ⱦ �=϶��V��ذ���ٶ���~B���Ʉ�9�wD�5S�oh|%@ѳ�5�}�?�W'���A���Wr����n�ϙU}$&0�<�8��~ɱX�͇v��yz�Q\
����C~���p�.�y%
��9� o���=
��	��fN�s��	1+�S&�C@��0)J�,Ǐ�4}s6��|�������K�jA��e,�va?^d�2��h�2a��|�=�s�h[6��sk�g8��l/��xn�˳"Kl�����T�'�qe�#ZDf�ꐜⴝ<X���C�N`�t�j9��]FѨL7d��^��]��?�H���2��/�)K�_ު��oNoř���XQB3�x��N�\$|w	Q�5���WL�*��9G�G��*�
��e=��9)X����{�:7�@/S3	�&r]/�hP�~�R_lzR�/���4���Xa�a�bnu{Y��:G<�=�+���
��9d�;��b�%����x�
����G<QƵǪ��p)� 񷚉è��>_b]>�I���{�C�O�R"N�em�D���b���u���$y�EQ7�"9�v�\�͓d���g��c��q&�`5q��h0� ,���A��9V�!>����0���N���"�I�m]��*�G�`���H��@`�#"n Qw[��)Od5[�ql;=�3���=��^wlR��LF�.�p�Z�5ZzS	}�Y���&,'w�KÉ�g�X@E�����%{j]���d�.��+n�K�f&�0Q���`lM��n5܁��n��\�%��@�U�7�q�0"����\Pǧ�]
D�s`n����z]C>�8�tV����勵��@�9��#Ib��nx8�A�ONͷ�#���S�6Yiڀ�5��$�qN��\���x�!�gG?�LZYt�����QCt繽p�VBV�]f�t��#����	���2xIo�
X�[��2�gݛ&��"���n�{	��B���v��.�`�i���D0�"/py�Y��x���s��L*B|��"��9N.�r�|�`������8�д�}<j)���*ͬݹO���9w��V��_�qx���Ӛ{�J?�̀� ,W|~����5!�us��d��
I2�f�J��+v���R���P��N�$q��#!Ʈ��ǟ(�r��T��[
��C�����4�K�gF)s�,c�i�o��m�j�"�k^DG#n7��ih�It:�q�u���&�YC8�
��)�4�`V�B�c�5'xr���ǾSχ��X��/Q@�7�$�a���^��_Y�p-�����P
&Q*�P����_�2eF	�[�ڠ���_"Ćg,8�Fq!_�ع'��@����b����`��w��B�1�/5�Gz�x�bP�0��]M$Ԗ������δ�J���^3��Ey!�<�Q�Q�C��&�nx��,����E�|�-`�#��ы
���j��e�K��yU����=[�cc��,Z_��Ͽ��w�
;���0���/Hs���M�����J1Dm�����>�c"O����%s�o�R`^|N�]�u��x�'�"�� �X[_��۝Wb8tHS�KE���k
G��z���� �\�@w��}���AKZ��ǌ�d5:t��#��+n�ڭ������n���M0ĬM��u�4���(-a_IB9���Q��.�ǅ똛{��Sz'�ĶTB���_�H9}��F�/��`F'ʼKJ�n����Z/���;R|X�`R� ��UY����߾5T� ��0J[��}��`�q�_hKP�+��@l����g�`2�<����<���><��,{0�=8��rqR �M�k����ƨ%�T���c��^�o+ZL}J�7�h�������C�us�f�B��&an
�뢶��u]��P�Ob�5b�S'�,��e����5pV�@w�t�新Ϲ=<�b�"k��}�nنB0�Lӝ-q�$C��g��ZZ#�1-���G؃��#���d�U���α�e�d��S_/�2��O dõT�:�?B���_�1Ǭ�8	��!�oWS���K|̐��U�r�0���p���E�d�iH,@�|π�F��;��P{
eSn�69v,�j8SGH�@d��w�w[�h���FX��Q;ǭ��P��Gx��2�Q)b�D�rimu�����w��B��^�ը'��D¹�ʤI&�%@�2#�%�plinW�!��tɪ�運/
}�p��Q���m.�eKx2s�הS���Dmx'$o��d��䒡V�5 ^�"�i�j*�;��Ї�,�ʪ7��ł��k>
�i�2���]7K[8_(=2ay�kVw_�xc�h�s�R-��#�'I16��[�t��C�[�����F��=�� !�����U�f�{E��Yv��\M���h�o��t<��Q��l2�m��~�]��g67ŶD��pj�}���tp�J�
4S�s$u=ݨ�T����y��)^j �w-@V��1�U���=B S�A�N ��wǌ����Y��c�$UJl5V�<��x�T��!��h�Lkm�,�Ҳ���B?�Pi,Q_�'��f���m�!�
yaM���ؗM!�ͯ��g�`D��Z�㼳��=L땼9�Ga���X�k�3=dJ��ՁJ(鄩#<w����ŬꪫOgF^\8*�]�z�Uշ_L�D-4!��g��l�e5a;�v�e
���%$�����Vj�`�o�a�S�Nd��m�yw�?p�8�3��i�ʵZf�6}u�2�ڟ|Bay�e+&;�Õr0��R���5� '��7!x ?JtKX��H�X0�B=ʅ�ܴ�-�);4ڋ�c�96"�f�Z���x�Wދ
��e�$�������5�X�
�����-·��	 �A����2�`'W���?��>����o������h�y�)�#B��Q�W�/��3���Ux̦j�G;�[��6Nӧ*Ю�v��mO_���"SїH�G�6!���^��L��d~%��ͬ���A8�����*;5i�r3��YH}9��2{Ȣ�)�&��Z(���R�JS�����3�8��1�C`:P	s�ƪ�y�?I*-���4�B�X���Toڎ�� h�\׫�����@�eژ㪩��*2Mø9o��3YV�l�K�x�� Qɓ\��R��B���ej��6�mh�J�6��WM|�V�W���r<��k`G�����WV�BnZ���	a��k覛!R��4���ۥ����	�˅�kR^!I䩼���$�q�����f�0%y oɢF{h��q���Q��?>v�?�F�OLB,X��Oz��\��3�V�P�9������	l�� ;zn,@��_T�ܫ��NWX�.0G��J�B_�/#�	G\�ި_e�#��-MŞ�H�������lH�>�'>`�ET{�� �y ��0�[�����i�qFd����,Tb�E�i��D8Gń�!iB�v̌ʩqP&�Vo7���!���#��⚺���m!�i97�|Y�&z!tܴ�z��tƘ�W1��{I�,�yr�}��0�c�{����X��sL��w���~B�zOG7�CF��t�V�F~O�WO�zG{/��ܗ�o+I��+;Tf�����ݴb����У�Ys�h��y@m�}�FhèaI��K�G�SN�%Q�Q7J�zI����FԒ��2�J��e�`���,�Ѩe�I��#�k�zM�K��3�s4:����F�Z��kF��Z�0�Ø��S!�hZ\|�`ӊ9�q5�1�,������o3��se�(�)S�b�E��D����a�m��lv�3�9	0]�wn����̧ �N��xY'�g鵱ʱ�>���!E�8���.$�ߝ��vd�%l�C�������t��gTzx�v���C���I.���%l��K�R7�q�)[��a��9���qoۈ:�S��x�g��NfY���a�&��$R!Z�������Pqȸ��Fw)S7�<�͞�{.D���ʞ5C��J|��I�==U����5k�z�2��n)�u3�#s�{e�5d��Saք���[�5���PP���ה){�$��]۠�� ��ҳ'� �;��H<mE��~���l}�g�k����o���N��2�o'0�Q{��ɋ���L�>X��e)�"g�y.����"O ��?�3����Ȉ���x�?�� ̄;&=J�|"X�xiC�˼��H��7��y̉��{����T8-q��6}ݡ=�:��xay�ر��)�Jow�X�������OZvhsxH�R4��d�uvV���2p��'-��|�ď�4a�RQ.č��N*�Wg</�����X��9�'�����T`X��<�|����R�5ˬ��7D6YI./x��/=��˛���-�H�i���q,ڽ,�f4^��e�����{ש�l!�`����p���0>[�"jCr�wRT�R���DP;o�N�Vi��I�nz�F��̶+��
 
�+��eӧ�W��a������J�J�dK���]Ԁ�
1���\�'�U�����}l�Rk�^�;w>ϻ+�jH���	
�q�D̛�]��y���føOx�S���z	TV��bJ@"K���&�G� �3V�%�J��
����ѯ@��҇����^�������Er�&�ә�_�L�
�6s[a���*0�Sa��ejI�5BP"��鵝��k��,��a|i�z��]���]��"T�ۤWu��ݬ�6�q�$?r~H�93fu��
�jeV�V-o»z���;,$�E��ڄͳ�mm2�������V�n�?�[�r%S7���G��ӆ����m�Ф?�|<�wMKzΎ�J�;x�a�N���A���N��������9=�4���\K�AY��Ӵ�.���|'���.�z�X]������}U��(��!�p��m�OC�1�r:O��,�k���\V�<����"t1�~U	��rճ�)/�ߞ��ՉCg��Ar��Y�?�-N|雋v&�.p,��-�7a&�z�s&�[:7Z<!��"�r/��lxE��
8YA�r9��&���9>�V[:�����/5�Z�(���Į���;�y�A���f=��چ��;�����vc=l_��S��y��<<Ƣ�ǔ�� ��Sx�y��<R3#Sbn����,��4�88�����qǥr?
�)ǻ��&��Gӡn㚑�u�ba�!�5|��I�"p��W������;��#�w+��2,uA�=8`<��ܷ���BR�sٷ��2�b#=´�P6�	�]ݞC�S��ʒ'_��\40�?d�z�-��)�tP�&�YK2�q�R��T��$���|�[|!�X�X�E޶3��S�p�k�άmH��O���l�"����Kt�m�>�}�Kh���2W�&������vts]�B��wm1A���13�)�cL'� pe��c�Z���L8"��3��f���&ա\�]�Xjٔ�çm�zGRE<�Qy5��'Bw���J-˒
�+���ps�4�&����&AҌ���ڦg}�}�Oh1@R��-�bP�����^?h.�:zJk7��"�i���*�[��3������Q�ʵ�ˌ�s�7ޕ3��^�v��ԑhZ�;ʑ�yˏ�,U� �O{�D��œ��έ�:�sTS�����'�Ӧ�J�CLٷ�`�Z�@�p�e�����%qh��� Һ�dn���F�n���t(h�``�Np�#&ဧk�E'�����{k�5��SjB�kƄ�scR�E���9w��yV�n:�B�l]��&Gz�q��	)�ݔk;Z�/+�'����Yq�I�?��c���-8+|^�U3[�Jor�D�
@�2��0���8O��jf����Xd�Y��ou�.A�Y��^M�#�p7E�H}��[�^w�LEFd^�kSiABӯl��v���^N���M*��j?~�,cq^yh)�Ғz���?���,�����C<�r����]@�)%T�\�5�W],��?(���_� ���
GsO�#�e�):'>��'�yo����{sԥ�o,��4�(՗k���/xש ȱf��(�<���!rKu�ٻh��c.i���+	��
(��<D� U&V]N�x����>^��i�qS�J��#_���&��|k���^'O���������o��ɼ�	��6���W�w�JP�?��% :���!�Fq>�����(=�z��L��}!f��w�U�qP��s�ZzI~��=��� �}�{�p���D��� 7��Y�QS���$����Y���T�ZuM�+E'�V�A���g����"�Hg����}Ǹ\	���I���N[���L���6�D�쮜��
D?�7��G:x� h�^�0��PN�~.d��G��e>�9՝���B�cE��&s4�=ԩŶɗ8��k��O�v�/�9BT��Y�-��\����g)āuh��(r`PK�TL7�4�A��l�S��
O�U�6ȅkEs�����˿����1��9K��1M�)Q����3@�`DXܾ�	y�g�%�N�7v�b�>��-#���4�|=��t���Y�4"�o�#&�[�.!�&΅p�S46��q.Ϟs/O��e��t�ћ�w�G����OK`���緔�>�Cq�nh?(j���@�����-%}�y���z���5��^��.9�G�S�l����f���dFF�|՗i�3a�C�;��������[�i�k�GR�]�b�����e���Yy3���>��e{
�f>���S��oE	Cڜ
�5:�;e9�Bf�$r���ytcu�G���>��֑0�"�[E�H�y�~Õ㙋C�Ag�4����Mc�n��Jގ9V��~�AH�T��C+�6��,�nQvܾ���y��� ��e-�v58�R�!�>|a�į�n��o��i~�(�w�=���E��5��VM{�FQ�ʻ�]�ѣa��g]��� =6��*�Bv�T���}���j��4��]�+b�WQ�!A8�z�k�n ��+a�ĥ(�CDYd�z�(��_^�=^��}fVQ�n�����v��N{G� ����Sǫg�>��3��C�*�h�ò����ץ� Ŗ���ǌ�I4�hZۓ����A&���=�{���e��uWB��Er$���%�T)u7�f���)�(M��*�M�� H���`��j���k3ֽH��jf��z_/4�#���n���3<��K�~,��C&�GH�D�e�.0��lÀ�c�������H��V��F!��v�߮�ܒ@�w<m�����a��$�J�jZ��F�ay���zE��1��ˇuq�-ڄ�IHL�>�0 �����Ț�����I�GX��L�%X �(XC��ՂGVdm������|��.�i���,����{#�yȃ��s�߷�p	��mco�r���$��]Q�Ћ�#���㝧bG�d��c�v)X��*(Q-�[�h�E]z���pټ_W�k�����r�1N=d��pm�M�ra1r��JB��2r����~)DY��v|�>�����ɗ�	��fw�BK�ә�b�,S1O�mYoO�;�Ӈ��JMa�H{�?J���q����/0M-������"Dw��	�	k�Q�ob��1%���I�՗Q�2���y�k(8Ň9����ԔNe�woJ4L!�~���a!H�ƏU��!�@m.�a^'�'�p��ª���v:�1t-Jniw�S��� �5����!$$�\� ����/�q2���.*ijO_�!�䧉�%LTz�X+�������y.=�q�.Л7a�Y]�l�������F̠�^��X��]���y����`8���@�
�R��Þ+	G��j��M꟢��	��D�3����10�r��H6��6T��+���j�ۂy>�ˆ�X��A�/�Lz�w��In�oSl3�*� 9��2�хa;��� ���(�s�K�0q�/3��v�Υ7����w�y.ih�Ӂ��֊c�S!K�Z�jWw�a��p�c����bY�R��&Q�� k?K��1^�ٱ\�8د�ʏҴ���'�Y���� ��J�9	�ۣ�ƙ ���]�P�e�+4�|\8��M
��},�z��~a/�2gu��� �.�;��w��#O�G�]��̫SW�|��>��l�I�_����B9`nR�z�x�v��a�di�/�̕�8O����|@6��Šj��g�SL��"�����(u8|�G6�#��b��_��S��A�<�4;����R~�&������y�(�^��Cy��0���A>��|����m��d�Q9k��s�[X�ȫ�> {�a�O������t��ł�[:+EH%��<������/9��X�%)3�|���񮵢*��_����� �1hCO��3�hL�Mm�qnH.�l���=P�M��ֶ��R�H�H	zc��L4�w+\�����%�>Z�>�7U����D3Ж����<bܑ�VUK�i,��oHβ��T�>������gC|_�(��]�����/��	���>��%1T��۸�]��Ǹ)Ok(<d%ǎcg��c���1�m>M5X�KGWIn5��J#�UEc���l̢�}��VZyXӞ�Z�_Yp�/��ɺ�ʃr�/���'������X��v�5bS����C��!4��>���5��k�)��|x74k[��X���9�pu�K*�e6`�hj4�Ċ��<��B��=�4�LP�Q+A$ت��S�`+��t����<K�3[1d���Ϭ�J�g��m����
��d�j>�U�m@� ��Ռ��S�6
��݆���J[]�k	������^��(*�L!��Tt�ډ�1J�P��#��_��<���_�NM�Oz9A���wF�p�ح+�O0<ބO�v.|]����,x�>�$%f	W�	���Yd$W�����K�|,��AM>;�AmzBO���=��ͳ5��\1��4}��e8�[9ʻ{,��N����UE�zn[�S���Cӳ_,�|��c�_�
G/�����;
������h������*�_RB-��^���;����Q��]�翷�,�<��!@%?,+R�n�"�`����-˺�=:��f��/�;��g$+Rr� �i$��x*"���״C`#!_7dY���WT�W4�]NF�������ɒ����>��ϯ��wt�0�iw%�@*ؽ2��tx8׆���4G$	9,aʽ���^��Ƞ<W�4����D����d��wjA�8�8�,F����������;3�X/���A����}᫰��F�t]�g�h��i@�0x ���嘉�4��?��Rn��_Im�{�P](r����5��;�>9����We�Q|��K�'�d~����@��+�}�,(4Gx��#ڱ��ؼ�v˻�5-ԟT����a��q�:�e��rI��B��׻Em
�U�D6Q�*$Д�����0�S���K!g�j��T��'�
Vm���� P��̕륆�l�����ϚQ
��cA��x��¨+W���(��}��ɯeP.��0�
5�墶1�tz��n�L�n+��-~�d���)�A�FBr�顦<�g���.D��U���V)_�V<�_�坠>5:vڹ��6� a��>�l���`�DaL���c��g����q+���2�����8���^^9�5���:a�Z���^�����A��5\�]�0'���>Z�'Z��ΨyU���թE��Ppu�}e���%�Ϡw��d�r�µ��7�$�
��~��.�PXj�zw�ýi]O������r�ny_���C9�������A7i�s^�8�xD�W�vP)�����I�
K~�a�{��EhH5��F�*��WKT�TH==d���#I; �S��GLȀ�i�ÏZ߸�%��Uu7,@oW)t�<�f`i1�4�86�OV�!J��0.{�I!���f�Z,p�a��JU���˞��iYR"P&��ٟ�4XQ��8�F��q�,<�P>9�NTB�h�O�|7��o��L��Bѵ����֗�-��|ޯ�6XY5W�>I[';�?�������[�]	O/F�i���=��t��	��#���K�+ƶ�,��5��	����@՚`�Juۙ��R3��[*q����X�[��.X1C�u�oQ�� ���{c�0ȧ��.Q+� ��D�)�.��s��s+�����{��5��Ǖ����X)�\��UOy�逈G����?�&/�������?�6�dGC#�X�|,�QQ�O�(QV�OhF=��+W�A�rML����N횄T_&����N«��fmB-x��Q� c���y�*J����Q�F��s�L����d	̻m?�,,��|�o���svD�'s���S^��~	
�:/[�5:.�;��<z���I"
6��sa�8��⒠�$�Y4�6ȐuZ[��S@��o�r>N�������A��IJv��"o��x��ۤ/0���!ǰ�P��4�Z�!���5HMt:�9�j��4<[P����A1�.����]�9�	GzE�~Uh)�V�]����^}�ӕ��	�k�����V��>�bF���q{S���ƱGu"5��L<�q,B�^b�38��Fе�Y�R�枿ëQvP�&���Q�2T]�F>��GO�U�m5q����p�\V�G�A�;{>%s��lۻ�}u�<O �8��&=Q�@
��`��>��>d��l��~�۸�s!��?VE,ͯ��5\���sA��������e�4�,&?�ΏW�_ãTNAz���G��Z�˯���`%��Q�����>��9���#�;az )Uk��݆S���9�y!m����6�-J��C-#�	��R�E��'�v�e�]i�K�rr����`�� �Ɉ6���5���n	5��2g�}aY|�	�[Ȑs�ï��z3�X͘I�aM:���	�����I(��a����[����*����W��R�5+\�^�2����3�h�j�&�lc����U���-^�>T�V�c�ʼ}��Y����R6~	�����c�b��o��,f�j��:��6u@t��S� R����O}w�6���t��ec�ʹ��r��%Z	����x֐��}};���h�D߶���"v�	w��,4A7�+n�]9$9���h?GK�(R�ǫ"'�0]��W�H0L�@#N�\@`�8�3�Y���X��Pj�!y*�p�O�Z~ S{Db�<4s�'J/:m��YM-nQ�+k�t/QOn�����M��m壻�@�����{`埘�*���gzŸ+��oLG�U�ΐ><�{&B�"N
l�2����L-�`�Z���4PRvEr�Df�Oc0��"�ބ
.�Q�]�W��y��|�[-�����
W���x��_&��x�Ѯ��h�1e����y1�90#���,�}�w�i������y<���o�D����u��=b ěJ�x&��b4}r���\_�ml 6��yFD���c�~��{|\`ճ�p�5�����.�{sm��O?������W�	̟���;��u>�@��v2�9��A,h2����l����(�3m��ܲ��Г���ؘ�%[�ZX�� ���bN��B�̋l�8������3g6[���Vn�����BdU�	E�ɢ@�<(1-�^O��V���&�>Ë{=��ߒ�j���0�_0�b�j��J�,��+��ّ�Ӓ9�Ѐ�'r���М*���<���U���E�)}��tbW�P9�Ƿl�BA���&*�@EܗyWK��Ε�Y��v^+jL�A����d�vP��	���EWĤ|��Af��������-eb:ty���(p�m
[�4���Dq�~��;ƨ�e*�ؿ�Q�������#�x	���������qպ��S6��I��2���G���e���1M|~c���z~jx�|%����C�50b�`�o���%�m=��1��J�2	/�~U&�)�j�}j;I�J/5�h����A��I�i�T����3�k����x���G���ژ	Ƹǈ�#�h��f�"F�T@p�7�j��U�X�B`�(\%J.5�N_��|���dr"�C9��L��
��� �B�;_.�.�%N��+��RQ�����'C�W.k�O�~��U!�e�0�rHn+��gU�l&�9����=�l������9���[���gKĠ�Y����-m�9(`:�� � 0�S�H������.��#�p�M?�T]�aƉ�g�}:�et��ʥ��3ǗK(Y���L��ƃT~��˩�h�wн���b�!��87<h�ݮ j����U�LNN3m-P��`��Ǒ�O���^�%�^�?�u<�p�TU�|�Q2P��D�AuS뗉`���ehz$����	���������g��D��Q�ϲ�RǼ]��uLIHU�������GZ�K��S��OF�pX&�F�.��E�y]jTD��dϜ�#�P��c�ڒ��H�R� ܝ���_��{}l��b��Z�������;����-T�y0��]cN
SP�[3^Ƙy�0&�e��ό\�H"T����b/LxԵa��$��o��yě��r{�e6�\͔j4�_�zr-߯�,w�]�ҕ؁;�_Cr�)w�0��*�H˖�5"b� yQڶ;�@�^�U2_����C��i�?��C�,���l\�	�Z�0F�vÇ@Yx�[#^���0��5��A� �������!,=���C�ɜ���I���Qj�7�Y�id�	ni�u}�RA�����Vң��{�G���S�t�D��R���N���1?0�n���#�|�HY&�'��Q���F��
^�Fu�`I"�t�w䊠�i � ���O\��h���gYf����-gS��ޘ�.�:%�����_2^[�i���� 4�kŊ���Ǝ�݆��ӊs7�o5�zLI��żz'k~j�F1Ϲ��ɝ�?�����Ȏn��0��0lJJJM`�~�m�x]��g��`9�L�yn -'�v�g��?�6j��E�w�~M���Y����I$d-?��k�a-!�/<����	~v�H�EsJ3[bb�x4�i��Y�GXfm��C�Z�Dc�i��zb�Z�p�tq|�c�X�h�ȹ��6��:�-`'p�m�!���
�����\�5�s�c���H�V@
���b� gt�`��8�@f��#.�?��,O���qg�H�j�~�)t�!	%�R���)�o$q�/��'��Fۇ���;��xr��z�" ]p;�mu��p�*X��F)y`]�N�����X��P�8���*H��hC�(�#M}@�Yn�}����P r \ ���i�gȆO���Y4��L�O)�4������r���u'0�;���4��q%ҥQ�9�(�P��Ĩ�g��	�Y��fN�e���Nia�f= �:�=t�	�i�W�Y=���b�%�1"�7��^Xl�]|sﶈq�
����T,+tN�+�o�m+
�4HV/�y��^Fl�kq}.��ߧ�q6�t`���B@�e�ۤ�mO��4�@&х��5��o�7�ܬlGK�
������,z��OńQ��Ď�)�;�B<r��8RV�m�BE�`��J�Ju0�)7:����pkR����oB�������a$Sᐍ$�(_Z'��6��׹��a��VYw��j��vw:�*)s�?��0X6�O��~K�t}��1� s$�#&^I7�$��f�3pno䞧�Tj�o�>�ʰA��T�]a�|�Z��g9p�]�&%�Q�2�Y���rS�v?�빝���mX�����8����6i��}��4v�ȡ�wI���|,-0��v�PJ&�2T�/��b._���ዡj{C8����F���0�f�ź�N�����S�88Pb^��^�8�F����c�n9&�!gQ���&!��%딾�%�G����#��<b�e� -�A�jl�B�3R�ev��@iq�d���Ԧ��tG�#/ujȲ�R +�S�6M��_vc��ۺ�X@|È�C�顜0��2��P��9o�[�@^tU�nBs�)d�����a2�a65ZCTW~�<e�6�<7�M0���]3h�7+�d^ej���1�;��ʳ:l�Gu�C�� ~��}�Iӛ��Q��?��8�f��s��[�z?f�bÔ�k�:ڂl�1�P9�2Vzޠ���E,�ڵ��;��2|��]���%�����,C���dR�@�r�(�9��xUJw.(2��Fde��-C^Ȋ�>��P;���Z��+J0��	�4� �R�J"�}��M��tŏ]�`C��<cA!:��=F�,͐��vjˁ��I� ���ٜ�]MX��C�e�٧����\m*���>Pc��v?y���=,^�D���>���ٲ.����o,IvM� ᔋ\DG�@J�E�/�0�z�:����R����n�KVs������R�ȭ8�%P��=�Fd����Q: L���h�XP�� {�!���VY�d!]�o�{�Q�ܫ�A@+��K�c�p<y�����s":�bT���Oh�̀�S�Z�G�H{����1�0���`���*� ~r��X��W������i���ܚ�An;c�7�C�d�MI1���k�G�����s���;­�`�u׾�3���x<t��:��\�64���"����Џ�ʤ/bHI�֐�mFyg�`�0�1e�4��w���U�l*p��G�2��1x��K����ɍd����xO�FϺ���̾�4�b��-X�8W'Ph���Quǒ�_�z*e�86��zf���I�G��CB�6�!�NR]�c*�*�4y��޲����ߟ���)��#��fq��f�sO�Gb��0��?����~Tc����ZR����ˤQ�e�G}�1d�����.��,�K��&*w<lAXf��.�W��3c�Nƈ�p�/f�8��u#��Mb/q�!{�4�����ۗ��"/�*� �4�n����{s>�czD�~��:R��ɠ���|���+��[���l�}�+��8�qq�kn�B���2A'I�Y����Zz��|�(�ۗ`�Y��J�g�(�bt�v�Î��.}���r:K�
K���� |v��YdrpeZZ�ʬ;�)~1�ڑ��8��߭?T��5qE���D���n������ rk��,�/L6��CH��-XL΢<>�biSWcV<z���=}�͂��Z}�]wyv�_U&@�F��X�����B�A*�o���n?0-�K�i������RL-TW�D	��Μ;�Es�?!���*�gj���q�"&+!Է�٢�GN�	 �M��D�]WAp�/<S�����\g�e���tG���ev�U{k����HK��o��fIA(�d�Y���Ԙ�05cO!�yi]�-ԋ��+;�)���^k�n�R]�.�����Q�?e�ش�̿
������J�A~��k���č�{Ӏ�����c{1[�f�_ʃ�nÑ���K&��(��g�S8_S�#�}2�`�EӨ$Vl�(h}�����D+��xFCt�����#pE�h�:#5k���C��^��}����_��,h[�rYhV63{��0��e��t��G=l2��]�7�i�4֍ʠ�����Q�[]哈%�:�`ɖ�����x�a�ݾ&z�#<�G�w�|�q�'�3?�*��V2�ө��և>-|�w/g��V�g���42-�Ei[�Z>�7��)A�5����>������"qV�*.�⪳~F�U\9�x��+�
;��a�H H�����ýN[���)jݠ�|@��ء*�in�/�����ur�����[�pj�V&�2�K�����S��B�[7���/ύ4I��M�{b��u��s�+�3x
��~�.!�n;�[��*�'�~��.0�{N�.R�j�he����"���w����9���3����qnp����R���ܳj���k��H~��G��/��s�7QbG�juV�L���<~�&�N��y�(ؗ��o�Lԥ(�����#���)��t�
�w{qq��'೾+`N��$��r�й�dw�6�4��/K���
h�[C�r׃T3�݋˘�1o�xs 4����L���
#�Ξ����=-��[��Ҡ�m��Xv�78@�JiA%<�;�I"Pш�V؇��<�%�s���j$)R�CDV�Q@��.��^Z�1�L�O!�a�:T�۟K��\�}u�{���	7-L�22ӛb����� Z,�������Ƈj8)s$� ��h#�#���q��J�gs蟎�'���h�;��:�L��@`/<�R1ĬKIA����:��r�2�"6E[}��2q��!ӣ�Ȧ;�CI7�^uw��q�m�&?#�� �*�bg�Ut�uW/�C��BF[�rdw9Q�8\���Uh�����Ɉ7<!�@�fe���G�������C�kl&�.�	D��e%��v�"2��������#;;�ך���M��}��|j�!᧧��V.�ԓ��"D��[Uk���u#&�^�8g����@���1�Y�5-n��+;s`�/2��:�M��T�!G�^���.��8��+�c��}��=���=��=��r>X��BX���D.�,ߝ���Dؒx��&��9,� h�Շ.����\CڵN�����&Mv����*��a �K,Xн�d-�OFն =IX�\F����������x0
.wh�.sPGjyh	;���+�ݗVJ�����Է��z(T�2#呖���8?���6m�s	�b*����$��!�]��m3"���KQC�������_��ï����
�E嫁b�E����F8�K)h�hL���@��Q�	��| Ռ��E�F?�����ދ�*A�[3�r$�Ƽ��\0PU�[DQ�>��cP���ȴ@{3a�v���=r]�g/��X���L��Y�O�$�R��<=��Y�z���]�vj�3S������03��+�Y@z���z��j#s���A̖.�;��"@Fd�W8m�&�A�υu���l,� ON�(�����j��o�X@�W��|����\7���ܞ��i�{��a���D���,�
L�p8w�S��_d�0�9�Q���yiŇj|Y���C[py��ֿ�|ڼ��A�� �І���J�J�4�hx�J�E�Y#0K�j��e$�	;�q�t1ͥү�y>�W��R�p5�2+��V�e�&RFhsV=��j�F��N�s$5	A�-0���7:�R^��q
�[��osu�v��j���Y�+���<��i��?J�E��q��t�[#���������0 ���(G�h��B�V�W 2*��3�<��ͬ��lxW��j�XD��6=%�5�a����ӅŰ~�N!]_ѳ5S��|��K�X<]����':��Pg�����g@�'��$P�彗T3$���j2ؠ=f���?���l~6��d�Ś��o���ƽo�	b$E�5B�»�`.����$�5�V�WX��'�r�?���R���6��"�Z{�_)�u���1E,��(��;�-��ħ��k���d;��~p`�l�(Ħ�cMțeEAh��j�Z#d��.ֻ�ݗZR�u\��Ѫr0�n�,��o�r3�@�eǭv����ٶBZ�@5-q���|N�d��ل尺	�Jn�	���>e%>M�N�m4N�j2�����K{�ٓ9��Xn��_��荹Kj�ȴn��G��I��7t����EjQxf�8iꪆ�o:��x�TЉC6��!l��:������$l��C[{8��������YƮ�b�v�#[�dϣV|�/�rD	nZ�Ӽ���p�Gq��S��w�`u��d��(O�	
Fl�T�s����C������eHL�規���A;d��p�.P�o�w��oQ����ؚ�v�O)N��������e%ʏİ�����1�%Qb��'�c��Ʃ����]H�Z����_�􆯟-fG��y�
�j���g���;��~ٞ,f��Lj���9I#�}:���;��=a�h���,O3y�y�=֕����#\��-x��K� n��oX�,�]�GE��A�Lm��*1�\����� S	�2v�k�q�R����}�oQ�s��ԺI%�U�E��eOT���x��2��(���������^<F���!�24�^�m����mE��Mqj��C�ww�I|!�$��i�
��W���8�!��!�:Xl��E#�)O�F��y�A�t��p�c�(�8ǽK����g�H�=D.����][�v��.d�e�5A�". ����6J)���&'eW<�}0H��/�٬����o,BG�C��xN����
��E}��|E�I��a�����+6��y6�a��@z�U��T��<�{:�"�b'����۲��Gu���ܝ��o�B2�5 y����_�m�0p�~Ew�t��U�/�^�[�W�cV�:!
Ï�Z"u�8G�M�cx�;i�Lk�Q}N��ArжM��xK�������&|z���A���_A��r���"�Pc�K���Bh&�HaL^�&.���A��4�k�5�؇_�%��������^���v�R��K#ɾ��A@Qq��۳�t��y�Y^%�_���9�+i��U"��h8�J"�O�\Nt����~2���36�M&aY&����U�>�
{�۲@���׻�"J����\��%>`���1��� ��ƅ���z�8�I����P��G�+�~���|�s�/�S+��Vr+�ԕ8�<2}�uFO'eޝ�i�Ѐ��"�=>�?�$�m_��}?������0{Ͻ��)���k3Y���{����J��\K�����=��`3�0�N�XD��>gr�S��D�wgΡl�,�T��W�l;Kl��h5W�r@NhQ�ofI�S"=�����B+C0��yz�xg��˝	0߹ָTu>��aA=�M�i3x�!s:3nKF=����h��|y�8c��L����J�~�
j-2у�uvK	�Z�S?I� >$�=3�Y�������>��B�ۘ��R���V����7����8z�w�5L�8{��IYMq�bE3��L;�+)�J�,8�����7��*�ӺHm��:8_㠆��Lj�Cy�Usĕ�WD}��]����p��R�ރ����!�r\�8bk��.�*�͆O�"���l맟�G�ZX�b��@:��\�ZZ��V�%�*�kőzo����e���M09h1��B��4)�T�/B;��L��nO�+Le!��p�|�c	����������/���Yf��}�6�`���ܻվp������vW������ҧx�R����ٌ�I��4�͡�%NƊ��ǐd+��G�V�ӿ
H �r��g�XtIr����d=�=�|h�	�
�K��ʸs �vT��Vo�7�Y�Z�X���I:t{�+P�{���iR%'�0�;�T�'ۆ���u�6M�%��m
Ï�)��\u4ڶ�[P�IA̟���+�g�5��[�ց�լ����A1�7�9�x��: �R�m<�	�[��@����:&�����+�cm�� L �Y��*F~�6�0ڕ�S�s��'a���+sq��b�%�&���������O�A��a�Д!����#O�h�/'I9��Q�Qp�4�H�qMUag	�Yu�q��{
���/|������"9p(�@�j�Τ{�Kj�����K?03�U����C[�Q]e't�/�
v��\$B2>���AeB+U�)�Mk3�咆I�)	������F�;W8u�L�خ[�Q���.Ȑ��Mm�����"���ԯ����x�CgB�D������i�l���5��F��x8F�V=f(&�����#�h)UF]�k���G�8!����2!�E�J�%�<��g���~2���}�&0*.ڃ����¶������Lߛr�����-70��v����7���:��;�m��M&��p7��y�ܻs6���a�|��M�2���Oֈ���l������ܹ�GDe��+Qw��+��'�{���dދ泬�7����@%��p�@�0M_���s"u��}�!q�� -	�M�[r�g��W��h�=3�q���죆��[Mٷ����ј�؇=̣qh��+�>�������)F�E���w������j��h�E�(%�����0kptE�=��&^�@m�>�&���ƜD\ܞ��1b,s[�`Y^o�U�^�mV�����b�������`�=ws��,���m]�l�ȼt��W�'v�U�a	uc�ɮ�Q�^*���"F��՞:�H�rK<�,Jd��(��x��=���r>L��Ma�W�3�q�ϟv�+tG��R��A�����>C��4�̎L�
��vmqJ֔�=B˽!��_����'�2V<�Bx��ND�'���>�������>��_M��MxT8UK<S> .�~UoN�1�Ai��Ϗ��L�=D�II����V�w+�XCU6�!��)|e����Ֆ[��3&i���,Оt�n)X����nk���"8�5%�o;�'��������=
tzV�+���H�7� Z;�����k�@
l�K��pG�
]�vՅ�UKo��z�9b3tz�mʁ,x\H��鸔��h�'�/*M��M��*&�w�WC��.?Ǳ���&��Q�vFy�Z�a��ē$�H%ۄt����|,�";�U.M��B�E6���Id��i�8�@�c^tF�V�0��B�n����9&ɩ��	�V޵a/�2�jMO�8I2�,N�e'��D��\�� ����8
�~�[Z��㶽��R����83�L�[mRڞw�е��&A�$ٍ�/�u�n��������'���)���/ӏ�S����+����&�EW���gv-!�EџR1Yr��Jd�H ���	�EЫ��P;�g��N�����
P	���k�dOJ>N��^�xΕ}��)�l#��Jy��>��:���c𑽣�'=`b��o/l�y�T�o��r"~�C�h���9�:P�O�3�~��łZVk~�K�M�����9�55��=�g���e��27Ve�2������쵊B��}��W�_��	R1E�9~��C�����r:�=�`[�o�NZg��:�Ơ�Ç�W�LW� �+�&�}s�����V��1����UT�%/����U]��&�M<$A%A�l�Np�]�P�;��R-���>�հ�~�_��v�(�I�z�N�:��9����p*F�[l�RJ�a� Y�'�ix"˱ŗ�GX?�U�dґS��;h�U�DGH)}>���By�����=��_I���+��-��l�@��đꀻ]�u7X���Y����l�<p����I�����Ê�U�6&�1@Xt��hA�۩ʑRfX� %Zf����՚�
��}�شl���~	�xM���1�YL`������̗��xk��^&�;P=V�� $��
-�J!�	�5h�5q��j��/��U�}2�ij��1����s�Qkp�Kp������};߈Q��3j�8�f�ê{6l�e�㍹�����sd�\
`$������e4�	:���_HA��%��L4�G
g��z�hQ�3���ۇ9F�{wU��.!�Pz�5���>D~�z�ןD�-��8�]���X`����O�~�-���*)���S=!/Ms����(A�7UMQWh�t'o�y�0F�^(v��uO����$�y_���6%�m�F�7�S�M(����xn���c��O;���^�>�=�&z넝µd�i�	�y(H.���b��Ԭ�:���2BH��s�C
�0mK5.,��Yx����.n��䉺�d��
?2�> �l��h�hKU�/�|��hս|E�ɔ0V?��v�#̼1M-{�o�!t��
Hֲւ�YƵ�Ϋ�	K
���T������̦������o�R4�@�ުW��/��>V����	3��f������Դ������G���i��5p$o��.����@.#��������Z����ag&fʫ��vt�?y���GF/�R�}�V��tK�GTmGŻ"(�T:�5��r��.��2�h�_h������������s��i�ұn}�����*� �p̢:�������S��\���@�ʩ+J�Y?��u��`1tw���s�6|,Fn�[/��A�ɏ���� ���>�%���oH��ORR
���O��U\���gW�����F����%�p2>�e�$DP�4����z�X�b[��FR"}ֶ����Y�W��?)n'�Q^����-�.�r��ݤ��2�ڧQD��D��͛��LѾ%8d����Q/@@d���=�7�P\�*��z o�'�ZcsE�ȓ�:={P��]�f�n��q�|�� ���j�<k:!�v]�$ߡ�~ؒ^����7����`X����M� RP��ؖm^�N�A��Tt!G嫸��X濕TvP���
bښ��NZ�A���o�I;}H'����N&B9Ų��:RP���G�	h6�&]�m7iw h04�!����M���n�a�'���U��N`5�UvT�ng��T�P�K>�<�t�R�\UU�����f�m�Tp��9Vt�X���T{h���ym�?��� yF����T�-H�#��W��)�A�H{���G�Y��d.\g�|������smD�R���(����p�2��Z���{R#vЏ���v�,����W��uϲ���=��GǶ}a+ע�r���O.��yͮ�y�%;@�ix�at���/�[F�W6���6	�41�5j�i�����7M�~{�q@�yPS�rP2\T�98ߩ)eIwuK�6��^�*��8��el<p��Ӥ���JQp��:��UX�:'���V��.�Zm��h��mP#�/Q���>n��0=1���V2f���+3مva8~�7�����fJc�{喥���lb�`�<"��G�~$J�k�∾���^��ũԜ���[��Ū��t�v9�yC�Έ���w�p��Ֆ;��9��W*y��*h �	Blx�����TI'��TϞ��������n��B�*�m��#7X���ן[�q7���~p�1?���
l2C���>/}�rB���酉?���+7���'݂jh�\�\jWa5u���'ƍUl��S�Fu!?�
���ka�1�E�V(��Rv�%Px$��̓7/� }����!�����7!�$��7a�OY��+��a������5*SR���_���ˌ���;iCh�vq>�˙Ȋ:-s����q���=uh���s�%���L�aN��"�r���Y�P*t��O���4a���r[
�"=���>�"��K�R*���ͤ���<�4�z�`q[�<ُ�#���a'��@;��=�l7�:�C�J�̩)���u�d�z��_K&�aI?����cdJ���л+_�M����V�z�Nۥaφ��'�i&��YO4�[�M3�\Ƀ�K�x3/f�<C��������t�$�W,��Og)9,)j���d�,m4��Ӗ��!�
vO�2��\<�P�����'G�k������'����36���w�����t����8�8�{��@ۗ�B���]/Z��jΩ�`��'K�����V��:NI��Ä��7H6��eIڲl�#+���`�)�r*��ܦw&�:0uO�����y�g�v��La�2&n$+��w,2�O��(�aa�)\�7��D#��7`u����`0F�i=�g��%Y� �2I�N' ��6���[��@�z��2�����H�w5%�]�Mb3:zf/�(
�����~�'����R�>��?q�e_=��J!'����#X5��{�HRv|ZŐ{�*&n!w��a�C�Ȭ�	�[۬gU�C}m:I�顃��B,dK���+����7���� ��������45\��� yo%�g�G+�t�S�тkcv�5--���������]�
NNQ�M��S�jd'fƕ�}@]��������/�3�]�2��iD��'eQkS��%
�ذ�)�4��N�U*��Pr�T���e��)'�#"����$(@y�x)zm8�'?%]��D�~�<�xG����32�cy�қ\}KȟTݧ�c�|�E������י���y�e
^_����*��g�x�|���iZ=� n�>��ѝ�l�)���)�q��6��E����sB�gK��Wj��@�f�"t���RN�mع bUq����aq��H��g�:UF27�:Ն��K��\�,�iQ8תG4o���T����� ����8�Mo���t�����F���%Q��Ђ*p���Orfdk1@(�������	\s��d�e�OԏunWp劌b3f��(Ww�O���c{�T���c0����Y�V��;����<|��k���5�d3R�a����	�
C�u3�6�c��>d�}��ٗs20�u�;ބ��No�����8��X9v�
h���q�/� �G�f���qa��X>�*���|�|nۭz��SL���EТ���uί;�b;5(�M��U��!ǭ�cd��.ͽ�n]��z9R*÷����f�7,6�hi��X��� �VcliW��w�X a�����hAx�������n�r��LTC,6^�q	��غkS����?TB��y�]��~S�[/���>�F�,���w������{r��䬺��r���=,�}���R�O�!h�Q9?�KH�"N��{�C/_b��NH��g�����)ˁ�-��j9�Sw�WLd.:BP��,?g��һ\�)]Oxk�@�z��Z?��s�S�Ve �9σ�G
K!j�V�W��Je1�G�r�'�IU���=��1�����1���f��O�m���	İ�c��/�]��J\��S���8U`#t����{�E~���#�۹Ϛ�"�:7W����q����q�~)�:��u�FqZ
ɇ���v��>��~&jF������W�u ��/�\�Z &�C�tO>��yj�j2A��Q�Z�ʏ2����T7P( ���&�Y&���6k\�y���*L�:��j��Fz���p7�U��h��N~�Ί6�	��okC<x\aVSq�w�?v��ƌu8�:&��E�_��Db�R�������`K���:@�1�9�B�b�i�8����9%�� ^4H��Kh���_�۱`\��g�4��_O���hO�h2�������|ƥ>���H*�u�}�H�&��h��?W1욑��/K< �\�"E�Y57�d�w����x�޴g�4��4+&6����rj��Ղԑ�z��yOFH����ʂ`k%�\��^��#7�c)�:��l����^	��.ّq���F�E2��[�5�5�/��@��s�K�.�zp��ӱ���S���zi����d���N,�-�F�7�:�F���(0 �x���!��C���t4�$'V����x2�{���<�Ig����.t��ܜ�G���4>��¶��"@*�xK�C�p½�ri�����G�D�3����%J�*r���Ĳ�Y��F��� �DZ3��Т�-傕�F6����4 ���>�\�3��X�8�&rY�7?	����$(m���)�.�X�rIC�*���gL��3��b���g�|Vn���3U�lsJvৼ�}	�� j?���v�S.��` ]��i��4�g>�r� #v�=bYA۴�F�\�cD!�Q�M��4�f��u�����CNȚ��b��R؏=)���w�:U��(?�6�,~��"��նe}`��t�G���ݦF��JGyP�N�X�!T��U&��}�fߠc���KgeC�(���D���0�L��`¼7�;�ݓHN�:��s~�kmK$/��+$�ىN�i��Qb=SkTJZ�'�5)���TѲ���
�ok~���HӉ��I���J��_+*|��ǽ�7���4���(�>bQZݳ_��T����O�!^�ɀa�P�ZQ���i��g�}گ�s���6����5C���4�~� �k�+�	��䞥�i���l;ީ�����hq&�k�?�}��^�^G4�E�mp���3�d����2��~M��`��U��wMMݐ�9z}�.�ڴ��0ߢ:z���WC�B�X��.]oƉ,{#$�9��oF�C1PNd�JTAV�\�w��/9�(>|��	H
_��s�Ik���l�: ����"+��}P���;�Fs�^��c)�j��Y�	�1�L�lFu���x�/2��ʉhS��������=aut(�q�p�q�W�����)}
���k��$4,?�ُ�5s���z�ڝ���lȧI�1^,w.~�a[P�dh�l�5	A��D��g3a�����jI?� �툱j��Hq�S`N&�|M�b͎X���؜)�%9�>�杁u�� hy��.���eVF��G3�e{��>ƾ����Dsj�Ѫ��o)��ȟ%	F &��ۯ	�i���`e����u-�HDMF�U��垚�z�鐠��̌,�W%F��a-��e��+Т�]"���(���etV�	)c��bC?@4���)
�ʚ�i!�[Ȥ�M�Ԋ��!{ �6i����<H7�m�3�#��Y0��!�;N՟a���|L��:���|�j�Cu`35���#
Yޱ���]�(۝���z�ؓݐ-��A*�1Uz�YWæ`�+dv��l��ݭ�uS��!e�yd8�HA��ɄYc,U�I����BGeֺR���_�I��jU���¨_�qY�i�s3ҫ��{ ��m��E�����ޣ�X��K(HNt���X�"j�����i��\~�J� �]����t(t�Ll:���>>���i�t���hd�'f�cw�W-r������<o�a�;�
i��?{F�P
�����K��>ߓ���(Wt2�6��X�?�Ra*SKk	V�3�fU�-wE�zCѭeg�`WM�F�8�*l �W���	P�4�"r�fVc�苩⺳��/:Wq�
�w�R�s�:۩�/��9����j�-��p��F��-~�&y���7�p<i�����3����b3O�q޿�OXi������+�Y4�H_aj����*d���=9e6��z+W�r�7����}��:������3�q��&��|�ib����̃^c��u�=�8w��N;��]v��>]����� F� �O�ױ�����������
3��˩��%��[��Ō���ͷp��؟I2����M$Q�w�#2�C׊���4�_0>l(d �S(�r'VLڝ�粟¯�Ґ!v�����9�����-a�V8�&���wsZ���spx�9�V|�54M�.fw�+zQ��1�ŧ
���k�(:�׏�\h�:�\�T�O��#���|�i�9S|�V� �j��Lo���Mo�!ϕ�Πo�����ߞҠ���#�t�\s�'�0 �%T�>N��z�UxH��;�}�4 l�+hf��cA}A�*�ڝ�R��_�$m��p2�^ᬈݻ���t`�p�B>�)��n�rb̡�������áK]'�$I��k�Nv���{=��n�"�[ZA�͝.��5��r����ڵ�C���Q�ɨV���g��?�R�KH� ��P(h���Lng���Z}p	)G�oS�V�@A�G�p�e(�\�%�N��7����(o�����&9�����q�h3	�=��h�A𭫍\�Ћ�`���������ݪ��{��7���E�9�T!������?;�d2��Kl{#a�7M0���u�@����fQ�㜻GW�2��:m���?�h�;P��)f�� �8���<����zΌ�;��r݀��b�q�SE� kt�FP-�i'j�*�AU���"ɣ�(T	�a�[�	�1_�u���Wut��sڤ�B�Q�ط�N�R+�8��cb}�4��������0���{������1${�z�]mhE켡�Ǣ��R�%��0y����1s����ʵ�G+F�-��U�����N�x�!hI��rX197��" ��T	̥{��$&Y�Z��Au��1����h�ٚO_���!�~��hD�xºT"�F[w��M�;�ˈ��N�rj�D�,�`�j��.���g��[%҂×���^N+�#�vO|�b�>��*<�7W�"�`�\��,"�_�\�������ե��cm�oZ�wt�L�$0��'�,�O�5恇$�^� No썘?����A�к����KxxZ����1p��2���%��=0x�j��S�$ؔt�PEY����wn[��J�/�.��z2G~���7x����s̖��ڡPY⃹�֒Л�.�~1�A���>$~j�����ȸ5�������"6O+�:�,ψ�\�������W���yV��KXl3jp��f���0��%Dj�):�a^�H�}��R����HS+W�J@�[���N|wZ&����]��^���!��b�fn�������	3V���M��Fڽ�����Fٯo|��Y��ZI���ь�Jb��B����	D���q	~G'��i�� T��0n�v�3�V�Uů����
�R�+D1�],PZ�61����^/qw�5�fO[�)��2@,CJ/R�B4�ۋGL/I�̈́�d��oz�=[P۴{�U�?�lzs����u�?[A���'�l\�T�2��Soy̫e�����B"ذ,!�n���IH��;b�4�t����$�v�$۲�,�>�P���AWT�������F��h��6/���|����T4�1�C�:��[¼���x ���-�R_���Y4H�X1�z�n���;��R#.����Yǖ�HZ�'O�m�\���[�W[7hv
ƴ���h�SƠ8j9�������%M�7{�dFƌ�r�}[����#B��\�R�?nJ���-������ h�1��Rc"�h��@vh36vۙ��5H�9ݢ��QIa2�$8� i]���@��7>�G�2�`��;�H펠7OX**w{Cv��h��p1z�P��6�˪�����$1������Խ��@��Y����p�������L���T-����B^Sw��|����[�[�CJ��e����@��lI�D;�.��4�%Gع�$zPt)i�͐j�;+)m�M�Πt���bL�Bj�S\�%�.9sK�yi��dH��hqWLn^�ܺ=H�ȏ5����2��@.B�)�߅��vř�Σlt~?����3	& �]�ê�g�|ѧ�e% >���т�wY�az{��H�9��	LBjq$��P"�hY����fYj�~(��~����%a��I��-`��A�SqD��੕r��J�*�c��ڼƔ]�h�����g.���T8�FSr��;d�b^k���_�Y3x���e��q2���r��!K4���n�p
��f�B��=�����-��p� bz��[[�$�������6Ȱ�݋u�-f_�M��e��;�1�:��OM�Rޅ�~��'�s�)Ϟ�Q*B��&I�ǫ�c�{���lc,��6Ѷ��e�Gh_�����4v��k�`}��<�Ʈ&��Lsk��&1��5iԿ�oH�+�u�~;�"��l�����z��q��"����C�%R�NA�y�n�&�R�������.�i(�!X+Q�1�CE���ŉ�{m��j�^s��@-{b���H�.A��'#�!��}̦�C��{#.:Y��'W^�'��z�^a���D|�Dt�3�yJ���Kg��mٸ�ֽ�3�Ϡ���Q�	�J#�#��Pz�v��c褻߶6RM8<{i>���!Z�r��`:�xu��	�{0a��>pI	�!]L�|�ĜW�A9��a�T7
`���=
'�}�x$��u%z�i��_�K��^È(#�(ʤ%�Lj����୿ힺ!��VX��Jz���E��$��?*�����[0��;�{�0�x`���V8�̉��m޾֗�,���ϝGͳ�qw>��ʠe�k�g�~�cg�e��Չ�"-��N�n`���	|���*|� ,�;C�L�b�⦷j��Ń�{q���W&��T�
���d���}�V�b�N����P -���D���pl�vg�
��̪��>"{<��q�9/�FHUR�T��!����n{�vg�]<J�.��uW�1���-ХQx�����O�#�����p=�u�[�,$���d5��i��j����cB�,DQ��U��6gW��r��~JV�t;�ئOrܶ�̷�ʀ��uh�d�4���G�/êB	M!�1X�Ҩ�]ѡ�9�<��Y�n>!g���+k�?��! �]��o!��M���o~k�&Rȅ��WW+�:u�[K����K.v|jgN<1��5��$15{uT�A���v� BX�͞E(��q��@�{��`�]��п�7ԅ���H6���LO�Ĝ�(�\&
���6
�=82jl����9�-�����4^U�D�"E}��V>���#�������\Q��[�%Nx�I�t��bċ�`�i�%+ٴ�t�<���~dX�%89kk�S��T]rk�O���d>��[�E��j������B-��N���&@���w�u��xo:B�%e���Js������s���t��QJ�y������:T�$�}��Z
��w���[�h���*��A�-��j|�}򏠀�]��<��_���t���V빎hH��k`�B@T��F~īK��$O#@�zsD�vA.�
Ydվ�w��h��:U�VXK��f��ڡ��'�|-HY*�6H"�`6�W����K9���EǄJmf������+(�(�	��SŜX��F@��,i,���Ñ�֛���������"O%��Dm�Zt�;��'�i&y�n���-��M�In�S���zo�%�O �7VzU[��%�G^3e߰E�8�w"��.rIiC�L�JRSphF��9�jU��v$/E�+��MM��T�9��^�W��ŋ`��}ʄ�PodWÂ��` �ܔ��A�Է�ځ	+�)l�����D�0��{�GrN�
��w]�(H���_j�r�"!�z>��4(�qӽ��r�s-��eȿ�~Gy_�`Gp�p�+�t뫚�+88��t����1E����8t[h!m���>�q���x�U�����Z�E	��w=��bq�M8�K����т<��^	�_��y)���ؽᗬ��)���Q�;fƇ��e������lL�Н���7����O� �̏Pd�%�;&��F?�-�8�93�@4��D��$ϐuj���֮y�Z�s���-�3�ALV���F�5����ݭN��l���E��d�0Oϝ0ǝl�KjYr���$�����*uv\�^R�)i%+>�{M$ŗ�l���V��4~L�ޑ�A�,���\�'�"_F~�CPL@���(o����6} iK�+�x뒻u+�c�������%�ȳ��ew-A�9�d?��2�QFJ�耦lqa�{���2�<R�GC��;�v>b3$���K��I�V����1b6��?nx�O/ӿ�i�l\F_o���%��#.%�ν��,��<{���޾�oK����r�i�����72�=c'�OT� �3[��H��nh^�=��������$_�-�y����UQ��\�b/���P_�_�����������$�f��� ��uL�K	p�?�����m� �8 �*mt����)Lb�v"7G]�|R"�;�����' ���>;%S�r��=RH����Ҩ�S��ƺF��n��,bژs��3�&���u�_e�8t�����f�����C�Kظ5D$�u����o-�]�U]M� �H�����SI���<+;��7��7~������:/��*�,gF��M�=����W�KP�.iB���ͧ竩�e�����!p�G�B8����	�h�A��h�ot�NA��@�ןG�o� �xe�j� ;|~C|u�������-��Z{�IM�)���M�(+�8ji�Ŧ�b��K4��^$5����U���ɆJ�V���ޯ-�J/���5/�[��O�?����1��U�J h�6Oاψc�LȲ֓�!��Y����D� �U�tGP$�r�p\Ba��g��e�Zy5�x�4��,�����<#@��sfʢ$�]�?Rh,)���
�^_R���{S�H�Uٕ0�.�5��O��)|�i@��;���nއ�_����M.C$]LgŒ��-*̃6a+�0w�zF�a�C�n�2�� ���F��o|B��೰<���R0��қ�\���2|�}�6��ب�Ҏ�V<.T?!�����u^�q����HaWX>b�v�y�'U v���o��]�|�k��uB���w��_��c�*��E���"'��K���
.��3$,ڮ��͜���:�;���:��1]�40�b��@�<�r��k?h0��bg�1h�±N2�s��S�x�^:g�|�����,�6��G���E D��B�K��3�Z��	/Ck���GF�I���tl&X�}Й���B�Z�&��7OfB�e2�Z�2K���[nq�B"���W�5H�Ӥ�Ϛ�'��i6����8��/�W�6�a�]�����Z����G�9�>ξ=p�S�`��N��^�~��_}���� J�w���ל��ڌ!!:]��`������+�Q`��Kxd۔�f	^��7K�z5)#�W]��s��@)���B�U������R-R�4��dk.`���ۋ�^]TI�NCG?c|pLA������0;I�~ ��I#l����~x�3�����1����%	��d����$>R��{��=�֯u9	���E��i�dV9�ـ6� Z�9`�[r#�C���e��4���{x���M���m甹���{��)r�a[�P_��;j��81|�I�%Q����ྨ�p��߀��q}�[1��p>&� �]-Z{3G��&�����FJA7-�������������)��Ej�7�d�niF:��`
SC�a��k].���I���1`�5ba����Ӯf���k�&^�`D�[���P&�8 T}�QB�q?k,�SҞ�"��Q��e�d֒��$A�B�S�Z�+~���V��|��RȢ豺�#�u�����=�{9�H("�?h���$qF{J�{����˿rqܽ�/��M� ����v�ŋ�&���{�I�ٴ�	|⿙\K�gWP�������U����/���7K/�"�wQ��>�CpAEk٧��E�j1��^��ⴺh�Y���/R�ņ��
O�@2s{V�9�@�?���7 K�F�Q�E��d�"�<B���[� ��jn� �󥈳L}�;Z����lpE�
��(x^�[	�*-FFR�s`�o�ˏ"�F���\̥��gP�/����?C�y�G:��ͺ���t�R�b+*#!l ��jNl~Y�hǲ{�V6�D�K^�v��ic�N��U�b
oGtv������?H. ��W>�v�t��֓���V��uƗVR���,�Xh�x/��E�vwxo4<��cq���z�g�#��J���UO�&Хw|U1֫Jt���B�4"������	�N��[����|��R2\}�k_lM{]$� ,�	��z�*���B�e8����ug���3�d��={j(3��7�M�r`�n�N�A��-�U���s�D�^��a��D��!��ofѯ�U�bM!d��oh������_�����\�UʣBX����6o'�b��Nf�<���>aò��Ք�*��ܦ��-'Lo�\ź�|N=H �r�[;X�6��X��;�%�Peb�ƂU��`��ށ��b�IC����m4�5%#�{���. �E�F�g1/ң<�r�9�tV�Rk����"����I��VR#��� �Za+q���E$�����g$��lu�U���T���آq� IZ��͸�j�hgKչ��@�(y�9co��ɕ��;� ��F~�&�ԋ�#�u�k��
�����1��^��_�UU4/�#����i��v���=vB}��؀�k������?�|ts?h�d��/2hE��ْ�]_��IY��D�b5#���N��+����v�󅩾�O�Rc�;��뎤��è�?.͉�%�e���8\�Rc{O��wT8'~ٲ�5�,�Z�.���w!�R9����Y��W�=�����,�a�Q1��T�g��s�k��%h0O�+	o��I��fh�K��A2H_4�Lt�w�7:~�s�^&�m��"
$k��;���*8	^b�݌d���D #؋����a���3�DG�mк�S49?�rtHxcZ��<w����@��Ә$�?��)��w�E�>�#�pJ��+���o|�S�1�Ɇ6p"����|� _ hu$�5�ԃ�p~u(ߠ�;W�LQtю�Uc=2�P0$#�mO���!!�W�ho��K<;$'�ߗ�B�Ԍ�P�o��Q����*�$���\m���7DM^�ee�(4��E�?_�F�
Ϛ�U����}
,c�[�u��:��٢j U�0T*}Ѽ�8��V8{U����3�d2n�U*�Ya�?|�?b��<��g�e�vd�����֧�m��8}�@f+�
?�	=����VtgzB]�#���ڢd��D�n�?�i�t���q���#���"!9�p������]��؆Mi);~^�}�V(g�Ɓ��'�߽��hB�"�3�. ���4�C�����Yޗ�zϰ�t0֜�-m�y��KIzR�<�I�{ך�����u�A�êu�oB' J���Z"U��x/܁�}h7 m{w%a[�	�rv5��5#-�0��ʛD�$0����6�<��?*}�����n���4�=|���s��'�vS6��8a��	�t��_�r��b$x87���/��S`	�VX.E �n��.e�S��\nm 7D�9N#6��I3�鷎�ޮ5ش��h���B��Z�%Z�W1�\m���e֩��& ���{Vh"�ۢ�W�2��x{MwI���'�Q�D���E܈����T�%6��2+�N����Uiw>���G�8�i�i��4����}��m���VpF"�
ؚ	̄��3����M�@#����Ha�ɧ4V-'�����c���0��I(�xP��UV�dI�c<v `*x��q�J���R��T��)Ɋ_��^ڶ��G�l�/(���K���ԶY)�{�'��?�j�JC�Ԏ`
��@x���qc�iq�&�=5�=2l�b��{;-���Z�ƚ��ŭ�Fyow���@/_�G�ulP�77a̾���+(�R��g=�H{��?���+�Ğ$�Zxs��5@r�
����]�5�oN��#�~�)t�u#5�$ކ=O���(O��7�o���r(���97��{��-j]�� h2!�r�!K�E��N�I��E�o0��n�E��ANAm��U���l�o�7~5��(�!�F�dW��Y�z<=��N���_�*���4��J�P�q�}���?�����.��7۸��
#z��AMUOR����,vR��mCu&V���e l�s��Mi��2q�ؘ4�BW�#獕Y��
j�]��>N�����*V����/'�pP�4�Rn�&f�/�W�C�~�^I5����v��2��t��ŋgߖ���A��?s
�A��b��� ����"�:H��>��Z�;��Ӄ�!̈́=��Ww�hơo�#������o��Q-^˽$jb�J��LB��)3Wm�o��"f`��=�%�(�l�tz���Z���u(4k�&���6g� ��P*z���/�ІE\�/�������u�v�F�y�@�F��Xd��BPl��8/Ch�C�Ә�G�D ����ǆ~�x��w�����-��@�GS\j��?�d�X�vj^����r�F�$L�oh|�O#��l?X�=|>N�!��o�-E���vI�ݱ������+��$>P�h�ؐݪ���Y�z��7x?���6�cD�*~kR%Ώ���g�[�[��l3��GF���3�۝67��UuO�\�����Wj��U�@��c����?�Qģ��T݉��ea��\&��w<��\��|�c����P#<P3=���o`�7*h��m��X$�U!,F��?Ǜ�ڹ�F1�3eSol��d��bZ�vZ���1jY����>�L2Σ�0����p�L��Y��p��x�g#���,�фP7������21��ܤ�n����j|��M��|�g�OW;���Gs؁�
u���*�g�`=��|�Cؤ��)��;���Yc�ߝqNrѽ3E9�����o�+���[��b
���	 �.^c`>�ڶ*.�]��I"�*����epV&��C���Y˷
�1)F�,�i>�d�7%��yc����Z��a��)�'%��dYC�,�!	��$��Mcs��Z�>]���Ը�VnW	03A�Y$�qP,�Pq���P�O�f�(jB�)���<�]X���M�A���N�2V��>9�s5��A7��V ��-knj�N��v�_�m�Wa�[����Z^���'M2�~�ىgL�.��3����4a� �q��NU&�?-!,ƍ�NLx%�'8U�Z�&��y=�У�נ�s��'�i��'��/�Q�p����/mV�̐w�׏�Q� �f}S�õ�턆q/��MR!ҽ7G*�ߩι�J\k�̓�$��~r#-�,	�#y?��d�;xR��f���S;S0�'B�g��@��Ԝ��M�8���kCp�{���B�����P��^y��π�ĵ��/��7�s#���<Y��ݒw�3�.ڻ�̆�M�}//�0[�`A���&�G�)�R���Tm��T�aD.)�Cϙ��b�W1A��]*]��"zV2����gVTQ���!�&���L�|��2����O':��Ι�IȈ��=��.�+	�v�OО��@ٻ�5�{��M��.�����_W8x�M���]A��F���-��t}AQ��~T���;��_Y�Q9䌙�Hw'[�4�X/U�l��%� [i�m��˓İ�+K���L梽��(FO��㐣��+,4{�WS^�%�*��5KQ>,I��M��d���Sy@fع�}����4�g]��Y<x�[~�Xxs���rP�/O˅	�b��U��?�V�B��*bA����s��SIHX���A����R�2����ç.�'ih�G���v�ŰsF�����'fܨ\�{�6mD���P�X9�\��b~�$ɚ�lQ��q ߿�6ǝ5*x��ƕc��F�3���?�G<���A8�gD�'ڣ�Y>��I�Ơ�����8��H>s�d&�]jx.�U�Q=��.���o�
g�uu�'>�����Պ�~\�ǩ�}ͻsj���G�P��}��Wib ���}?�4���� K!��p�₟|���gS���V�y�f�N��2�I�y���F����>ܢ}?�VW�&��J��*(�7m&<�ՎWʖ��#\�4�Gs�[�S��ѓ�:�k�ͧ�����vx�T�f���B�n��z�U�0��}�WN��'pz�.X��u˃l��FM��^ʝΦ�M �p/��֡1�������K��I�OX+�����`	������Y��'WJ��0��?�}h��>��b1�غC��;`�U[i�`<���������[<e%d+:��2ZM�,b�R�LɎ�P���˭c"��Q�D۟1����,E p�Э9Å�SZ��Zݭ�[o�C��x�E�!6��%a���F��.�">J���~���Ӡ����<>�C�ud��t�m=�@2l��y�EH�@�rv�O�T#�g�������dњ@�+i�9�?ZZB�G�w�����1�u��lq>��!9��Ɠ�I�;?�E��K�DV�i5���WQ �.H:2G 4�k{�����Ǳ���Ï~{��s[Ѳx��Of� 7�p!;��ġ����e*�^���>93��&;��2�!���ś����0��A��!����-F])�cS�n:�m�!�,���Ƣw�� �Z�F�/DNkb�eǽAu}���|�1�4e�_���5���م_͎.�~<Iv�2�N��,ǋ��@'��B�ғ�~>�4�@�����j�QT�>�
��)����g�K�ĊV�!��z�A�Z�螝-�~����zx�{�
 ύN{M��K�t�L�0�[#)P]y&����El�\����$K��`� �T�W�p"d �r{Ԩw�U����:�G��v.%���[�}ƹh��ӗ��PԄ�����.��X
��a]�ƻ��Tn�*��N`�N������9�e
�μ�ln�BjKq8u��6�yB�po$!��@ބ�~��b��j��醴L¹@�T��}{���D�D	��٫L�������jT��\��{�9Gw`9}q�f�[����
׌�P��y[t!۾P�n�3H�C�4���ԏ?�{IZ�-�q/UD?A{�;M?N��H�ms�� X�i���Q���T��$�9�������WdU�P�D��V>����n��uF�j��4���s�S��ix�)֘$(aɀU�	��y,|Y���k~~���g|�O��f���h�k}IV+��{��	���i�A��Ƒ���eTaG������)�M�������u�CtN�����m���??�%V��BS�fc�w!n�?F��qUqE�<��i��m��;XA1�qX�Aދ�ս��c?�H�
��N��,�@2�we}ɫÃ��0�X4��r��7��=�}V�����k#�V���E}B�*�����|���L�R�	Z�U�[�!��U�,�~�EmJ��|��A�����%�QI�Q�)����8BAR}�L�[�;|�~Ry�Q�X%E��v�Y�^�w�s���Z���j����7�$���36f6(�~O`M[ �f�8�����v�q��"H�w��#���U��_u�� =��& ��,�$�B|w���egh߈/���#�5'�d�6Ԅdl�����.5���$l���fY� ����6��^���G�-�k[_�c��b]촺}1/&�F� �� =`2cuٌ�Nq:a��9g�un��լw4�r���'G���ͿA}�'�%�~H�)��8�c1�F�@R]�A��fk�" ��1�1&m�g��16�`CX�O��/"۫��G[�X,TX3B��p��.��b5�Cϣ'i(�e�M�@�l9��S�ڂ�j�<��g����W��m�̌�,O�'�邌1���b稂 ��H�͢�Pf��s���Q��\E���-����+x��Ug��_�`��^�uw�;Vs��V��ޡe����d���?j vTa\��Z�wo{�Ur�`*���	�'����[S$��V�����>���v��S�����
B��x�S�)�eX�`�ߢѓ��s��Qg0of�1��5��o��E�xF�s�d�`vq�_R����YDL�T��.�%2Hzむ�i�r���e~}!�x�l}�$�P%�0ٖ�P�9���]E�Z���V�6wí%�@;�����	�����-aA�S_$��h<�æ^���K��n�㭾���I��`޼C�\&4a�؂K�	������+=ћ�p�@�ت��d�����2��0��5�`�z��![�
M��1%��:����KqkK�~��Gp���g�N��)/� )5?��[�MC�A�>6��Lٜ*�H@.t���M���>��&��bI��M2��Ϭ��:���d��w�qvie���Q	���Jn~����kBCY��
�	���G�5ۊ����E�Z�[������A�	����笓X�z��{���ϾI�?j�2)���R
x�`�=�Y�l	]�{��[F�OzUBQ�L+��GtC`�{�Y�6z��^��(�%~m�����ku��|>�`�r��Âd�(�5q$	�6��;�mZ]a��M�L*$0�3�[��2_]H��X�WF�8ˏx$y���;�zp�DT��	��5�]Ɏ9 jf�O���9A
6�m�xv����`��Ӂ���=�t��s�����o��ä����pZ��
�jE�-�@�G�.�k�c��&�<z��Zd��g��Ȋi�Z�(������[B�#}zؕ��
b}w�[\����%6tᮟ�����AIU�?im�(d����w�;��)u����`v"'l}ߍ4	��7;��w�Mx߮<�&�6�
��#Hɳqx:XC{�w���78_�*�I#U�W�����D�,��im-��q/���t��?5Z��;-y�6�I:�S/o�K�z[�MA7Q�P �\��uP�w��V��'�k�<���#n�e�V�j
wUg�cW̙3/��x�#Ң�]�S~�$6�
t1�=Y��`��W~�%F� �gl�)����������<���&�\��Y�q�c�T���?�4r[+�W@�$� ���	7&+�v-;)�R���=�<|y?I�1c��VtbTfB:��U6�,�,�I�����S�WE�s���!X���Q_�A��}+XI!���D�o�p�V[$i�����ι쳌�����w3۶[~�\�qe�b���\�kgPGLdNd��]s�J,8@�7�C&���&��0[zmi����W�+?��C�	?��'�&9�"�H�L�B�T$�Z-���d�1%�_J�q�Mg��P�Ȑ��W��K�|�gk�w�*� ���M"�:��{���$���1��b�d�U�M�w��iO�-��b��j���W�,'�A����\
uV��A�U�$S?����Ûh���[X��8�	\�Tk�=�05�ed�DyN&d����N�,��#����:����۬���}4
��2@m�c�S	�_3*P 9��=+PP�f)U׺�� C��%>�aFi���+��O���_�nG��~U��Sk���@t��k'� �X��.b��|m0�2�a;�'f�Qgc�K�|!��6��^��q���p�>�/�"��]�1c�:;f�5EbiyP>�c�*�M�3�=ma������Je�8P���5��ɦ.�P9��.24���eV��jʤT�F�g&�w��1eD����3�uqc��C��4,��52z߽7 	�~��s�Ji�/��b@���D(T}J�R����Z���??���}����d*}��I�+�O*��{�"���0�[G��F�n+��	��y'w2HD���FbRC��MK�E-!��5��✺4�@�X�)G���=�{��� ��7���b�S��q:e�h^2V \��'U��l�@s�0���ڢt�N����ؔ�(Lq�1�+�iq6�f}T�.�FT��G*"�ٱ�6�wuP�����_��J�/JI/��0�8o7Ǻx��� ����Y3��NKU�7LHv�)d����P��l�B���`��Y�J�OC3 @c�|�lzpE@W����ϸv�����ԋ�%��<|�iM�@�a�_n������՞I��yѽ����DC-�����e`�-��4Ē�=N?g�]s.��p��53i,FC�R�Hi#�j�T	�O�&��7Ѫ��Ϙ���9���0d�p�����1��C�����vƎ�\=��T��6ͨ*>D5��E��N�Q�i&�*N�� ��ì��r^���+F/5u�"�2qn2�	`�<����}�c�g\Ri�Ad��l�h[}3U�� R:���}�و~~��<�QJ����\��q���BBUR�I����
B��2D���u)���*i4���U��s��Z��K�F|xl�In9փ�6�x���4Gȴ�5&�}�ZK��[kM�9{��(����H��f�
�4��	B����3�X,�d��yC��IǶ�C�ܩ4
��J�n� z`����G:F�i=T�ث�;3�
������o����|�V�W����Ё�܋l�Q7���(G|:���x���<\hh;�����7>�iiQ�V�z�R������c�K�+�["�xG�syפ���8��[b���'p��ɬ�	az��i���[	2�b�$��}�ڠ}�u��2hj��/�iZwY
��0W=]�*b��G�&DYT˒�iߩJ�H�خ�S2l��Bk%��F�'�@_g�Tbh48���G<�o�קQ�K�,ԓ�7j~\�`G,�3ڄ��D���#�Y�z+((hl8.T����Xz�2�TP�0��g�����h��J�f��V?l��2�s���*Z493�d��<e%�����hi��63+Չɀ�Cto�U�������;�Uc�<���y��1��u?�Iv����v7��C�G�bhC55�rm��(k2���cU�0�X9��( �����!AVw!(� ����;��t=�X�@o-�+,�G̪ⶺZE鿤q3R �]Dҩ�k��)A&�&|E=<)�D��ByE�Ċ i�	0l��bvjV5>p��!������ܨ=��Zcl�SWJ�T9B$jp(\x���W� �JEH%���8��W�ˢ�`����w���e��P$��:L3���}5�Jclb�%j�I���_�ל���9�'�*5��
H#���Z�(ݒ�/��{�s��OI摲]��b�����l�A�wG��Â沋��p�5�#?C�$u+"�������h���O�� �::�1 !�����gp��q�n����e��� �z�좼�@'��J�ҭ�ȧ�p-�:����a'��0oq޾�A?���y�B�~�;:��9ŢI�.�*���u���&�B0�'�j�#��g�jǤ�	!e$ :C�b��$�q��{8x�\�[9��FVߵe�Bxp���1ǜ�T�#ZHM\:#�0?�_��w�?���V��c�ҝ}� �0�	�+�E� s��;v_��g��to�C
��y=d��>��!1	����a���ޚ��qQ|^#��$=�!07��r��������w��cU��@)V��G7f��������@�{�nn|:�f�i�u���Y~�e�U;=�-�g��o�@`1��4F�dS�(��=�n��G�>�Y6-�aZ<��v�+
�CL�ʪվ�.�Ѽx�ب/��J�^'J�Q�?�O�}�}�(��Xi��n.P���qP�.<�x���FFP��^涏}'Xh�D��Ƌ���Ϡ��o�O����Q���H���`���6gs��>fe;������s�o�N!\Y�rW��Q�C$C	;�̙�^;A���ܾ~������4(/^���R>��Hf��iL�X�����S�+�W�	=���?��H\�àហ�;G]���P��`�]����b����	d�{�+�3>�ndJ�o|8����M�����˽��j��k�p$��_���\�?����(�DA�&ӝ
��-
G[Tp�$b{=_y�gx��m��z�$4���U�\��4��N��@��\.-'�`?�*oy�22}v<8"�������j�����*=����9pRq�7���M��W�0�p�o�{ޕ�,�c�+�R��(���QH��X��#d����"���mж�].U��*6l~'$�k����Z�GPѨ���'��V�s��j�H�!�hh��kXy	ߌ��fh�I3}�ء���񾲰RӸ΅z�i�1�Q,��}�X9�"0������T�������`{ge�.�!���&H�j���E�"|�<�Sa]ūZ�n�#y0�'��Λ�f����	�;�Dr)D�m�p[��M4�Ѧ�,�(�0lt$�� %�"6���b�;�������B��n�`'�$p��x�=}����;�p�Ke�]o�F_M&}xTY�˓]����vO$��5솼_J�~��J֘х�G�G(AZD/�j��h��jلg;��?�LR�ng��IEE�$��9~��V��U�'��-��JK���̩1g6��TG�7S�BЕ��5�INFp��X��_�p�����ۨʰv�L��Wd�f��<��ϑ�]g��Qi�bc?�~>�X/�;�0�Շ�jw ��3׳knV���a�*�$�E�:�GN�ř�{�,�g�0^#2	Af٢���K��A�L�z���?�A"F��ÇE����0k��XC�\,ey.�;��\�����9R>����Ջ7�t����$�k'rJ��e�����w�W@�і��Z5���}f8`2�JI��'��F��9� ����&�Aܷ�9���{L���V����
�Ǩ]��i�,� q�+�X:�T�H'�H��c�3|��~' Ò�w-��
9���\��}��E;�����kw�G�Ǌ�޼�lSu�iV�g���AR�14g���'�Ÿ��!�]#-�?�	|�6
��8���͓a�=�	���߅m��`^�97����-2L�蓐>���9�����p��b�NZZS��Xw�P-��k&�ث��~�t� o(��S�a$].ة}�q{\����b^Í@FEO��5~2�f4W@��#Ql��wɮ�Sݢ6��y��v@R��\��@E%��Lb�ß�:�:�f�_�����xC�:S�(�*�0���鴦6�N��;0�#x���7\i�Db�M+ ��ܐ ���]A�?\e
ku&��0h$<�&W����eK�%�IN�~R-x��5Z6�s���:$$��'��`/S�"��b���?*�.�<S	o�Y0�����)�I��B��gP��q��5yk�����Q�ܠ@��U�����W��|B,�DY^���2��%	F�KA��XF,���1�a���� �}�`C����a��XH3��{��`���'<�D��J�b5"z�"��so�ȹ��[��ݯ�*�d���b6A�]]لkV;��Qߐ:�H�g�x.�d��sA2ɪ����R��ữHY?�3��͉�����/T*B��w5��
g���"D�Y��� ŦU���'>BN����u�鰤��u"�@�C�~7$�J�|��=�?������e�Y����P(|<��E��Oa����;�^���$X��^$�C�g1�@�B?�d��l�*H.�g�0Ȣ�Po�4���[M8��q��~ia
��F؟1Ġ�\G���ѿ�v�Ӳ(�"��Oh��2��7w=�w�U�0��o-?,x���Ŕ�K=� ,3,�������u
�A ��n+)3ˉ �r�?��x}y9�@T���~��� �h���B�H�"��g���=y\�*~���F�l�Y4�t.|S�1qy\̩l�Eԥ=w�c|�O1�F������l����;|�r�[�Rt5�P!X��� ���⺘���~�����M��<=Х���P�n�b67�Wv��7eį�{���-�g�I%X�DO��{�L�:M�sΫY��T����bƼ�C�ﮑ��O�?�:C[I&���(g�ъ�%Qtԛ빟�ْ/�Ԯ̝�C�x$�d�i�9�$?�����9�77��|�`pzY���*�ɒ杧!֊��g�)�k��u"�ҋ���{0�|�=�����H�VwǛl�*\�Z�;�cf�M~>�o�O����/)^㨚��x8�MZ��N�)��BG��_Zwu���x���و���W6��:��+|��a�`��S�2���X�����[
�S���XM�.o+H���d������v�o�����,]����oKNȌ���e�����c���ut]
�B/3�B�����"�.B$���<Z$/5!�}?$ЋjP����X�#��l�=qx+e�݊5�,?s�1�\}�� C��n	P[��!�px�5��]LG] ������rި-�S� �r�ݾ���ۯn~o�6���Qݳ�)y�|#7�*�,��}׉�����^\,,�p�QY'W컮K=�iE�b�:��ywKT<��jZ|A�
�Sr~ܓ.�G>E�6R�#F�\g����|7��m��Ρ�+�C�{����T�,�`[*�~@t��e9a���p�":L�Q��A3.��_�����Bu�߱�����)���]U*1�#�7�Q�M��" ��K~��(�G��HmM©�7�iG��ȩd��F�n��4z���VeEnz���(ph;b]�ĄY���	l7�m�׌�LB�ho��t뒛IC����z���ST��g/Ώ�m�i {l3ⰥK�ֈ�w��(hh��/%c7fگ!�D'�ߎ�, _	�_��ji���]�,���}��x�M sn��ϡQ�����h��O�� �	Y�-*����y�pϔ?��p��Z�'���Lζ�k�7$c�zG�/�H�s�(퇧\��l70�=8��#�Hj���/�@Z~e�F��<UL�<='{�d1{<ā�����0��@��8����\1ʍ,�����W���I�Vo��:%�a��<-� �>��"7⓻�xg�ݵ����
�-�,��u���T�۵O&�EW$3_Nb�]-�Yt�D���lAR��9y�V��\�1���o��s��7���$,c����~A�g|��Kp4C��i~��h��e ֜}��������*J��[�������q'�N5�*���?�X�g��O<��v�K|p7>%Z��L�nH���G*0�X�Cؼ4Y�C�����I�r�}FK 3tաO���F���3�i����?�㩄�+�M���"b���S�JQ�宁�9�c&!� %mG`m����F�Z�)��VΙ������/dUH�������I ̆�8!�Ā�2�P�Y�:#p�A��X�>��xO[e�E�����,D���-�yUς�s� ����csf���6���VB%��ڄԠ�d���Q+�]��]���6AQ6�3���&�{ԍd�۸\@���(����0���݌k	��Q�ۯ�'��	�-��B�����;E�_�%T����(�����d{Y�i��!1�4�����,t�A ��W�!�ȟ<�? ���m-;D�)-���[���F��Ჭ���J�s�C�5��Օ�	�̌�[�L�/UDx V�f��/Y�����e�BKA;���n�������Ьr�GZӇA7�H��1$Sd�H֣LT/:���0��0�t�@!������ ,{R)l%�_���]�ܢf#�7�e�w{�O�-3���?R�k��R~	G�5���0�_�+�b�@�p����uM�NOf�z|0�_��
�^4W����ϸ$��C M��t��yC�>P�����G�0�x?幟<��Z���q�T�{�0��uuf��ȭ�H�x8�B[
��)E�ܢ�~h�Ԏv/B�-��!_,W����x�|��$�j��fc���'=��Gq��k�]_/eSC��p�0��k�D�2���>�歚L���H�G	ξ��z�*�)wT�(�N\Y�TE�{� ��V��2[M)�e��0�� @ɉ�C�$���Bj<nW�j��F�A����N1+VG]Uo>D�n4�/��u!dq��s�"�-��>}F>:	X젞A���]��M �+�[�^=����W�iP?�G�ʧ��=n�0>��)�Wa��D�w���<�c����{��z�����
SuԼH�yN�"�j
<_��CLN���}�|a��6���@C��m�b�c�M������"��=`�����-���D*m!�U��j�k�nk_���*��Mă�N�7�d g��Oާ+}&�jD���[|�X�HMV�g, ��5H�|B)^r�����T=�U:�*(�U�rG*�<����Dc�^c�f��|k�1;�fDl���J8.���PC���LVC��}�(��(Qg|}�j���x��,yc�G/G
&iM�e�Wj�3R�\V�3����З�P�5����gYQ���2��*��c�bI����%�em0ji9v�o/�l���1���>�gs�fi`%�L�Ӯ��Vʾn7+DE>5�*J�Qr���Q�l�!�P�����@wGۈt�~c ��E�����/oέ�Ҍ�h!���<H�i:g���2%�>��'�ν�A:��,d>�8� �N�����~�H댃%s/|_�Z�"��,x v-�:�j�g}SM[�b3�^��[��f�,�1�ПG$\0��+��S��t���|��Q���W#���0����F��^��gTo�~Ad �C��9��7������P�|[B� 6�̺�) �{ ���@e�C�j}�u�� �#�ۅ$O���%6���a��qj�Q��@y��Q�58bG�qG�iz��C�b�w	��٨m�\�J�$��0<_���X���e��>R�fl��I���,������ο�I�/�N�q�8����k">�eK��,��%ף��e�}� g��?�}�W�����H�.���y��Y����aq7���"#�&�u�W���"\��{�'��0o���r�ŧ��(b&�M:H񱐥Y���T�ԁ#�=�~�\NY	�~4�8�FHK��{���@�ږ����f�x �O�O6qy
��| ��22O��x�k%|Ӏ��.@�+f� '-@��f�W�BO\�Ca]UJR�K�S��;�&"��|r�5B�W�ǿj����	�w<I1ܥ:�֧@>O��o��ɣ1��d��k}�����Es��Ԟ(�n۱:��H$�^_���y.S��J3<,Wj~�v�Pۖ{h�
�s.C� ��b��?J;�a]7�-+B�U�=(x	J�<x��.�tDP�88a+qh�X��%Ӣ@���s�+E�q�^��k�q���	]W�l��-l��IQ�n�Os�6�ڻ<�@���þ�s�u�lڞ��`�=r�>��R�ҟ������[b�$zT�����u C
Lǆ�?v�
����ӄs�����<=N'.U��
A��Y�{["����8�t��z�1!�V���q�ĵ�U)3�r�s���x����m�g�$�FU����R��T�����8��-��fs;я�3%a��vL��
�GJ�4���))�>pL���@D�)}�I�՟�d}��' ���|- p�d������ʈ14m�Qh]u�5cx���e�E�^4����7"){��5_�'!ȳ1o�H8/��%�e�
 �s!h�=��?�bJԱ'��ˬ�����qH���(E�=��,��&jSߡ��H�$�D��˸����,�4���%��6"Yy�SP�ˬ�,k�&��"�΍�P�t{K>1rnY\LI��P;mA]s㟃�@���J�C���m'B���ʂ�����U}"Ƒ.��b��@�AU�?�$銈f�/��T�o��!P���e0x✯阁���[�l��zt�s�zg$k�UET���6�ǘ�Y������ij���B�_���9H4��K��������E�_#�����о!#'F����������o)�<a�3^�����k@'-dH�o{~�6�u2�"��Q[L��GVSw��V`�w�#W�`�q�Hwq����Ϩ��EL�9-6�5B���vb0��U�.13�]��4�f�G�4���Fߺd�`W�$绻�_��ug��腤*�-��\��O�����(I,zSb���&�)7�XQF�S<P�*�����Q��`��B�_���-&�}��[K_�@�=������Er)?��/��< ���\0�=��0dt���wA�A�3���[��RQ�)D
�6�I|~�ZV�L#��5m�9��7:�\Ӂ�]朋�LW M���G���3%���}�;����0�K����Z�Ո5w5)mP�=�4�<��Wf�N�� .>s�@Дnq����ߚ5YI�L��>�x_��E ]+[PM)�4l�3T.&��K�yg�#.⎘��b���3�w�֌�	�!xT�-�X��|�Kcj72�OL��^�%qVv�X���6㕇�@��l���'���7�'�\� ,j��3z:�4�1dR�ێ�-�sԫwꯡک��
�3?O��[���l#��	]~_J����
'!g2����q04C�Q�����量Ǝ�$�2�����b���گ_�ꋌ�$(l�E^���(��shm�s�T����� 9ϟ�m�\p����w�@��!ZPE2�8!�|���nvK�e��<UH�ՅB��_�R��^z�K���h�����F�٠���	��$���0�=�M�Y!N
��"Ŷ�+v��GJ:R.R��ƣ���[%2�	�'zk�P֚eg����h����=Xl3��:�7�v�R�؎��".�7�[#qB[2�j��@"\)��5���6C�P�<�ta�❪�ءڳq��4<�׭��<��$i��9��CZ�n�_� 7��B}n�^������L�/�M=�9�q�F�P�ܹ���}��q�\d�G��`Z����o�Ֆ��g�2b�M�Ɨ��ɮ�t��~�/�_=��K������b�d�-� J�%��$�������R�����>V��h����x(���e]�:ۋBPpkxmrd"��V���*g��]���_�����5]n��m����+�#���@ތ�1"�I�Ց�L���`vj��P!�sf�j q��2�P%���@3 �I�#����"tq�/ևU���]U��N�(����|)���.SG�k2:�®��ň���(�5.��E�F���l-ϯZ�qq'�I��ʦ�R|;瓯�����B���&���b��U(��NJ-��V�~�9�÷r{�h�8ߜ�M/]X��V���,�q$�@ޫC�9��.�'o4�4|���Tx�J����S}r�R��~j�����O���ܣ��c$��-��0��l�~�3Xk��V��1��E�o��4����L[J�^{-�5��yj��G�E,���Qk*�,��,�i>���&u��ݦ[��	�����ጠ�_b6ȇ�{�}O�뻮J0�AJa�_���l�5�+'�#h��@�䇐Ek�Ia$�+���c!�3
�z5�_־i�̧év�&���xpǝ�?��:;p�^
Â��Ao-������ӊ��iȫ]���?\���fHC�'�b%2�Wnw7K�����,�]�����r�1�셍P�}>#e�H�%l��vx���SVͽ��:�7H=�l]��Ci��N6�A��0�w/��cRsf�7qU{��(�C�k���R��uBm���0���铩Ogg֠��'Ԥ܄���I���kҵ֠�h�9$������Y��,��$JW���IeN�U�}7���"�n&W�d�v��;f/�0_���M�-�9c�{VۢG {_���ᨲwK�%&� 6�a���]T��:#?3��Dbbq�q|ҧ�^�
�f|c`��1z��- �JI��x'���(��M+�]�a��K]"SGǍ|��m���U�c��U�����F�@@Y�89sd�).Jp+ǆ1ڼ�~
U��Z-_#�|�F���ڙ��a�.$,G�u�r����pl(P�`��)\׺/�?���+4�(J�{���`�]x��7��
=�P���J��@d1@3we^�6o�U��_Rw�)�𐱘ٻT�ڥm���
�\JpBծ�[����=&*4�H+�cD�_�S���֫	������}S�Lw�5�ˤ�Pc5�L��,�ڿ������w��F�iؐ����i��q#jr�/,�)�W4�+��xl���=�g���`�����`�>~Q.��c0Ũ��S�	�gT!z?Z���?��a��݇H�<�<�hb��������"��7e�)��@�F+� N1��Dô���l�8���#dϴ�g`�����.�K|���k8b�b�����q��8���ٲ�
?������k&����;�p� �S��?���@�nq���nUNL�rf���,x�d��Z�2�C(�j18��v�bNyANS�?Zh���z���{NH�sT��m����f7���OeD�*f!����+�n�Ǳ������o�F��U��#���qM*�rHQ_����LӲ_�b��\���\��xcp�$X�18�A� {�6��{����!J����:�جS(��B�-$��8���>�����8d�b*s�@wn��F���c0�iDL2J��;��ϰ�`PR�;��$XIv~Thq�-���됊{�kuA]0�,ۦc+\�g����L�9NI'�U��"[�K���%6���r!���P�����G���T��ʋe�N.*���<[1:؉�͘��t�X<��ҽ�d�W�KOQQ`�`���+�b= qm�$�9R��o:�=("��<�e=��4������i8I�&!���[��6g��2>�G��[`�蕴9��Q��*Dg:J^ ?��(y$�>ι�,ݘ��s��D����0���$��P�s���BPiLwG�������*��paPO�ۭ�/��%}���o5�����s\@5�����d��yF}D�5E�"/'�2V��T�0Ě�JA�ю:+Pm�RN�$*�� ��Qb0�G��g	�ޥH��>�Vg-j�4~n�I�.�L��fͧ�����o�4(������v�c�����gTd�cHUP��+�9_�/l���֥�b�eM� 㐖��h���FT��I����AoH}��F�z� B�`1���Z��`�b5�
�}D��6�x�V��<0iE���p�
��}T��w�������ŅKr�}>�0����d0V����0�oML#U����ݡ�����-��C)�j|���b���,G�N(� i*џ�4+�Q/�,#5���~p���%B�w~��C���Cɮ��o
���J]((LT39?4�W#�%�^}- Q�k���x�a4���^�[�v�~�J�i�{�~���.��V�UH�䴘K���Jk�	�6��e�(J������;_W�<*�i!��K�*"��7�Z�T���>��h�teM�}��*
���&�8���ڂ>��xQ5�k�k��� L�=�*RACM�:<~�n�d�i���G�^��_�}h�#���:'pK�f{z���9��{��	c�Rh��t��)m����=N�{�J;�=��������P�~���b{�}���Ui�O�|��Q�Omv��l&�)�a��E����8�c(��)�s�\�fz��W�LhJnؐ(Z��0o�#��v�8I�pP��D����[��펠ڬ��y���4���T��Ӗ��Z�ED+�#��I�����O�8�o+�Q`0u4 ���� �p��
��aq��G	&����k\ѝ���I�v�>���I�����q�C���^F��S�Є���7�R�]2:���P����z+r�N<��Ǐ�3fi�W7d�h�-�΃��6:��Zz�U�7�[wP��g�.�����Ɏ��@g�='���a5dO��;�/"� 1�&͆��zTO��A�	{d����Kh�Q��
B�KlܠMk�W��׷��*�&������n8U��%��pavpz92�yC0V�T���693j�l�z������=�LW-��)�]L4���to��!��e�7(R�u�����ԎA�I$�Jn�q�i�[�O�Pg@�ܬ$��9��!L�R{\�X���&,�Ƙ|��������8�ji��)'A�k	_����8;-��1�̷28ҡ
�-W�/�B����=j&QJ���=�M�#�'G����e!���Z?WC%��QRǸ���{�m"c��Q�a)K�0����a,�8�	�dN��:@:@�n��B�[�7��$����Пݕ��z����0m|9:"U�u�����*0����(�A��hT�o4�~LXxf���LUD[hz�n���Fd��FpX���Ѳ��'�I�����k�	Ϗ�'>m�bܸ��;a)�b=���w�NBї'�,XJ�k��snkZ4�� ����,��=�6

4��g��r�d��������ɳH��1i�j��}&e���o/�oԳ&
��Bb��/H�ȍY��2:孿ϑ47Ŗ#=�_ �U)��c|���x���6o�ۂ�9P��i����7Q<%e-���aVJ`�K{����V)�@9�+���:軀`�Wl�WӨ���dB�x$�V;���7p��fRh%��Z0'��9���Y�o0"o���Ҵ�6�i~�@����+�P._��m�%ͬ�W͚8�u�lܫ�fq�����̳*?�{&,Ђ�U��5�-�X#��Ú7@�ȓTR1tqT�ի;�`PXH�"��?�r�Ө�[�����h���S�c���1�&�丢Ky��<l;��;»ygV�k���r�
�P�C^iC���;�ϩ�Y�϶G�^�B�e!�Z��)�g���V�e	m�a�m7�l����w��*�iB���	p��1�w��m�����XDIi����k*.�u� =�ÇM�R�ʷ8		5ti\5!~̇��W�˺y��e_�h������o�k���5p�G�2JX#�#�$g��eٙ͟��=u��#Tá���8���$�ӯg<V��7x�$���	�}У��	�l���*���~�ЋK�����i�;	�M�/;8��\�L���.��ڪ���P��Uŵ���صt3*?@�`G)���=��;�ۜ�6��/���o"��w��x߼����Hi�V}�5`�Yd���[�\2�[Ee�@{���!�꣎��X!���� �*�x��>|�Oi�����Q��/�F�h��
��x��vpI{�;k�*���`Q0�=2U��E�לđ���J�~5.��j/ˊ��z/V���c5�X�T~�CUF�4���b�:^K)\���n#��M����o��?����!��׸�H���iَ���״��d�FK�N��Q�O�Z; &��J�Q�K��k�\S]���]D��+��G��DH~�����!��_���H�?����pM��Ǔs\6�н�"��&=u��6��&k⏯�����֧��)���XA��y� ��X�ks�R�$1����-��( y��/��ۜ
Im{N%�RY��uyة;����P����QmNz�XW��:���v�c(�j���s܋���ƞaT�Gm� x�h�1`k#m�
%�io�\ὄR.%��������d�5<�!��R{c��'i���]�}�̩J���÷{��<�j�=B*���s��f��	�P�<��{|	IFg.!��M��/�V0c�'W
��#�ڗ���2 ���dD�V��_�ۯ�K"l���?�4��bYS���j�����>4ߍt���X��9�Z0��j��>I,�VR�|]��#x\�W��G��� L��������o��@N�W-^����<���b΃�l�񙨼��=_�XH��1Y!��~�ڔ{��G����0�g�D�%8&P�^�����Eg�A����&����C�j�.k��p-8�x��*ˋ��8��[Nɢ���ba|'��b�=�}2q��3٘�H�|w!�R1�+���,�ΥL�
 ��ܞ��D-��:�ͦ���V�B�����gG�]���3�R�����[�)Hќ.2C'�7�j�ʊ����;�	7Ƨ�-��r?Jy���t�Uߚ�]��Z4�b�1\����
8^?4Vu\���x�k�9�A/�(�4~Bi��c�q����A��er�_�|N��ܧ�)����AS��S�ݬCt���r���Q�8��p.��}������Q۬��~�^�t&S��0WnJ������5s�:���J�}��������jW��w��x�$�!%5ż��Ͷ)d�i]?.OHAX$K�{�L����,Ǹ��`Au"�8`�9+��;_a���sbfՉT_�r�X<�4���O�>����^�A@&�+��7�#'�J��^x����豒-}Eh�HX�$
�L�Pa�VT��U߻�uGdҊ���d��=�%ЉTǥ�pbds]W[��*��/�["�;7��T(����&<_�Đ�M�+��\'�����u�^�}�& Q��;�S%��v��[ʑ���٣'T�c��J<:��F)�g�BB��������!��/+��-
V�Q%�Z@q�DϠ�L�E�t`~u��cI�٪���[gf|#M����/�e��JDqQ�vH'��>B�E<�2 �Kg럵P��0�n�"d&��GR��9%Y������) 	0qx�o8� �&!�K�Y���+�?��"�LJ@�RϏ�#�~��b���&>tLI5���XW$�����Ⱥ�`��9�������^�b�$�
���DwΨ����������{k�Jj�?�؊Hh3��	f�`-��"�TK�f;+�s��ns���沐�q���������e��I�KFmw��bJq���3F�%�S|�,��1�r=$`�2>�E4��%=��w/�N{�;����0e�&�#@4Tk��� ������~{-$Δ�ڇ1����{��G����Y�W���y��`H��M���S>T��	?H�� "���\%��/t���� ������Aݤ����{��\3iG�����F�4�K�A�a�'����k!���<=ϖ@�vG1���+|&J�7�'Z�\F��ż����4g\��T�^6�G�PT��]���"��Ы/�~F��Q
���M�`��@�Y�;r�Oӛs�x��.!@���؊|��H��FY�{OQ���[�~��dɮ؇�̢R�j�`�� z{�����WG���K�Y�5��,��B��<�:"����u?�i�y6�V�K"q�XDYT�������z���~��Q�Y�)k�����A�D}]�#�4+&`�Ud#��*e(p�����Y�Կ�Z8��S�n��q�m����ݘu�P�#zluK&b�೵)��C������c�x� ���`0XX���S��}���ڴۈ\�jd��h�CԤ������[MuAx]�+���2���x��S���������X)�12Ω���o\��+�ދ�kgo3�[��Ār���P������B%�%z��Ӓ�@�2�s�:��ק�XǑ�?�4���јí}N?$�K���v���EoD)�9��ҧVn�g�p5������Ͷ!���,���U�;ʄ8`����RfQ��~�s���
�ШC�N�����ٌs=d0I�<nL�23o@�ɰ�u���h=<�렖	|oI=R�amrE&�� V�<If9a�����%�8�k[��h�]���z1hK|n��z�
����U*���Wa�V�H#oA��k�k�2���Mi�r'�MIѕ�M�y���pj�r�`x��^�L�$������~�HD�?PN��5z�� u�e�)�9��bj�ʹ*j�N����o�$�cث��n���'} ����Ҭ>ҳ��o��q#G���/s��0=Ĩ�$�$�Ñ�o��e�#�f�����? �bǇ�"�t���JkV6��>̐���0��D$�SLfb�-W�,�X���4]�|��R��&��XO�YR�Gщ��ܭ��n
�s�=��Yۓ]��/�����ȯA��Z�R�����sRg�k��hu�h��2ɒ⨴�=�P|#�x� � �BP��0�y9v��sz�?t]��e��7cҵb]��Zt�&�d-7�T�n��Z�������#>�M��x��3N�$�&�9�� �^�pa}���U�̚��n��l�0� P��>��a"'Q8٪_�YqnyyV<�XM�t+�kk�/�U�B��!q��B�!�JP�໺����H��N�8
d�<ڰ�e%V��!՚�u`r���@���V7��:_6E|=���~I�bZK������d8��,�Nӆr��#U��.�1�Cl�%U��QH��݌u�xr�(2E�Bgx�uV���9�~�\O��Q-�`_�r��S��*�P��P: Ԉh~J$�����Va��(Nkʉ��K��î	6;�(��	/����+ph��aqn�?W��P*�B���Zt���`�C�{]a?F����Q�1>k�n&��m�;���4�����a��+%�TJ�!�T��,����sⴅlÀ�6�D�����2xn���lK�W��ӑu�v4�r�0F�&���-�Ov���/74�=g�F@����!�|�Λc��g�:�d)��Ɩ�V�]��"��X�a��]�u^��x�I&��.��U��n��������<������R<�
'�Р}��;Ejٕ��$Lw>%���ӣC��)|4��D�oq;�䚶��b�l\������B A]v�k>��dv���v�`"�msQf��a>�ͱ�U0"�P���*���W��RB`�qD��_���\�� _�R�r�.5�Q�dẙ���C�O���9�� {w�"�s��e+�1Ŭ2y���4�r�r��?�����#�"�%l����MH[.߻9����Vg{����b���c��QX��"�b�p3�ًn��@��q�Ta,m޺�뛖B"�(�o[`j�mw�%kg��E�SW��z1S	��|��W^h��ov��<�M8��k1�Z o�Cce�4÷A�y�5 z>/��OF�J��Jm±{������U�Uv�kx��b�}A:���¬C����F���/�Z�ᚯO����p����IEM9g=9\�R5�_l��DN�Hl�}Y�bL���]�jedV^&��O���|wA��C��YzP
�����L;b�%�_Oo��2�;Ř+J S{10`�οײ�XIf�x���X�C	��O��y�J�ַ
a X?�P=�B�nմ2����k���x2�T�6���y)����^q:T2�5�R��~��"XEi,���9ǣJ��詢�ysج�j���k����M|�"��mr��^�|F�^Oi�=�"�o��s�5IJ����I��L�X2˸��y�BK�`f9�u���`��D�L�a�@�14��)�4y8�m  J�809t�fB���}���l������Mb�?]rEOVK5�~����S���ES��4z�_�.ʊ�c'Mє,��Fc��8u�=L:�,�r�'e	�P���L>/��%��t'.N8���kZ���f<t�Z1R6hJ0d㋽�
��	9���PѨ8�)��Gy��d�?@wO��+9�.C� ��#��^�7c��D.7�i���t��k�)qL��	�^^��"�ݚ��戼��|L��1}�op��ׯ>#�A1�o�Ɔ]Q�H��t,�b N݄ߧ�r�W���	���2�T�WT�3��l�h��K]��iP�:%򁸝��J d�����a��^�x9^�r�(o<E��S�G閊���e��0�q��]!:������|���v�� >�heh��&��=5��(�գ��B�YJxV�r��VU��O�j��Y,D����}Xw��@��d�F�k�&��`m��sgBz�ye�奬���~��~3��#ɽ��]��8ls�t�=��X�:E����x�v��.�/��q18��A�"pÇ�rh���(J�_�����{�C(������c���Rj���h�"v=���W�J���i�r���'E��*�8��.qO�&�4�d��#���q�:,Y���,{zxk��딄p.ѽ�����4R#���&9b��'b�MJ�]���\�H��R�@�?6�=��u���w�Ԇ�S�x�k��)h�s�g7�vu��|�~%IM���5��s$O�w�+�ޥ0�.OT09���PXO��
H����܎N�r��9���].�TT�G��,ƴ���h��u�K�F���n���<�I^\~�U�ᵣ`�CC�%`S.�α�0E�ϥ}3��HLtu���5|�YH�x	X�M¬���T�eo�y�]���m:h@�vn�R�`�l��n�;�C�&�t���.9	�EGQ�仔:���bB�&ZX�s+g�8���U��l�,�N��ӫ1D_#��Eͭ`�@�ᕔd�q���.��X�k��K
����z�R��\y�I��_xf���������i��D��m'���
����ފ�}	m�♔O��b�*+p��j!?��ר�϶�#|�>Pa�iWc���4��,��X�Z��)][��cYc�$��ƣ���f��d�[��V��Q��y��2�Z����H���7e?-�}�1M
Y^��~���V�Tʸ�l_��T�[mw�']�����%�+�w��\pv�O��o�b~��1m�.g��0S�:!�}d�6 H,2��CNT��q����I�Pka��ĉѩ8��>41��<�D�W�^�:�CD�Ìk��P�E�)N��P�����X�A��xi��@TE5Ѭ��z��-�k�3r3=E(�����EM;�h�eN��)��8��l�@��4�xa�t)��$�������R��k��Z�s�9
)����)ɍ&��e����� :_Q���H���ƅ���E�u�G�T0U��w_�� ����T�;�1�fFނo�)3�3��,���A�z)`�����x�.��`|rPz�������żC����7��te� ���D'G@���y��	Pdg��)�K��^a.��R3��ӳ����Y;�@�-����a�Q�,��2��w4%���O�H�<����][�+���.iE�*�SY2����e�QQ�=����&Jߥ�-F���YLg?J���.�y�[��2p�M�+d ;(s��E{\-�z,溡�&ݤ��Mvq0�nþ�NHm�~�QS�E~D��V�M"���DF��AQ˽_��2$�+&�;Q|�2�LPqŀ(J58�`q7��՞Y`2�B�����C�C�1� �	�ga���2���.0�.x�H	]���t��F�m��3����<	�g.9�Nw�yà���EAl�P{soѩZ��.?FXJ��Y�;Rn)�眚l�z����3�I�(N�?.�P����w�;��c]����*a
�%��0��67�E�h��&�Q�9���>�x@�v�g"�6 aD���wX���55�^�({���a���)
;�y	/��!c�J����[��.� ����OK�l�n�qL�|�}N"�$!7'�v���q�qE�:\�'�J�Q#�9��Y�kw8��$�Rב7�-E�QQj��~|6�Q#(Jٟ�w�0�HN��^^e�	#bY3�k�g{Y��u%�����H������F-ȗ���e"�,ն�v>2j������v�E��ѹ ��0���+g��o���Yg3t;��I,��+u)_�ߝVZ6����2�)�v��(��7�"b�Ms[QW}��1{�~����y�lZ���t�#q�X�
������eᱼ7ʐ�x�*�j3���#��|ր����.'	�/���Ax���c޽!�1�b��e)�m�ζ�/�Q{C�CE��ֶ��yp9o6�7G���mQ��F������k{�2(!��hj�
�hS魎���F����܄`@eP���dR#��8:!`'��i�JŴպ�z�Ɓk))�����.x�*9��'l���y��.��/|ʖ����v�\9j-A��L��+U�_��-�NI;F��S=?UcW%�D�� P��
�$5�=-Ɛ�طڐB��KM��4�N�H�H�\�rj\�/"�"�:��V�Y����x�ӻ�,oa�4�@�-�4�J���A]q��@�@���{�u�&ʔpN�� l84�۩�&�t�~�b�S_���c����xT�=3𰜠j��7r���e��G����;���iLb��d�(@dU7Q<�GW6YXj���mA&g�w�B|)1�^�d���l��4<w�m�c��?9���\F��RxV�j�ZWq���͑ˡ�5W��)q��� 5P�-���;מ�A7@/˱��B�6ÕJ��S1�@xZB2���bh�
��̀Z1�����P��) }�1$�h�}W(������P���y��b)s������^�!�Lxy�oBO6�"��T���.L$�z��ɢ�ļ��!�$Yt �SˎӉ�z	�O�DFm���^|?�C��Qz�:��6'd�q$���K�B�űirE(Mg>��z9���]��8	,O���G�ZۓB���G��e�is)'�<Ԉ�E��j�Ԯ��ĲC ~�J���Q��ߧM�$H��TZD@�k' ��8��-bRm�Kw�3B0z��p�#�{��8��j��`�ާ�kB�=@�A�=f ��ʽǑ������������_p�Y�D�C%P�������ĸ�K�O�!�{�� �>�������Q��������"�W�OW���,6�M/��v4���!��R�a�l��7�s��/�g�;{̜��C�_V����8�)��KS:N��U���l�G�z8r^�H
�ң����/RD�xb�O�^�2�W��B���Y�ڠ7"�Q"n��%��~�\�Qf�)��Y��I�������I606���A��Q��������t��H�}�p�qڤuQG��mB��.��.���\�+��ￒ?|���;�y���m��$wW�z0�_{Pձ�[R�N����J�a)Y�KM`��X|�H��:+��U��?/ȆȈLL�I�!/0!f��g�^��:_����i��H������w�
z٭s���~kW�c~�oڎ����R���	�:��\�Ԅ�����-W�!g��[�S��M~�>#�2���Z��̍��IϨ�C"8��8�G	�ssK�V� M���H;	ZtP%W�iͦd;�б �)2�Q�ν��7�ñ2�V�X&6a�T�� sVd��'O�V�\FZ*��G��d���}.gJ���OV輕�F��>�8�*�5�a>5;�>�U�,PW��<ˣ��)Z��ѣWF�kTp�6�������������{n����K���8U��fZW*��fdR��l�#d�uQt�+f���9at�l��aox`�9�Q$�*.r��ȡfq`G��y���a�g�u�X;e��<>ވ��c-��)t�5N�[ѻ�BI׉zퟆ)W�=cAb��������8ߚ�mUɟy�7��?3\���9�#6����Z��*M� j{�]t.���*�l�n����yP�M
��� �#T��=�u�&,��&r����ʵ�(�p�@�8eΖu�Pt��Y�ʮҙ����:$���[\�EI��PT�U��EW!qͅ�ޘ`���V��VE�N�$:5L,*)G�!%[F�21¹=���85�G7�XMT��";|�g_3����Q����L�i�R�7\��*�(h�"�+�֘��K�w��Lv(A��������Cx��{jE��/ڄ��W~��p�Ro�
���g��p���: SB��4Ys��q��V!P���'�/�{��֬f�K��/e,�KB9�����c�d����lگ&�yGs��5+Ԝ�Ӽ�X��8���#�(����Rc};?�&X�jD[PC�M$�
����@O�J���B��s=��NɧK 8�(��+���V�>���t�j{'B�%%��,_�����A�@%���N&
XC)<��#/o����B1q�'���?��Ō#�f�>b�M"�ъL-����X#6/?ʸץ���d��&Y�Y����n8�D�!x�Q�?2iq�	���qzL��r��r}�F�c*(yu`mK�Mq5෱���_�6�������v��Xp��k")Szqz"&<Z5�F�?������Y���������;.��z����i)�J��̆| ��df��I0&�u0�!�����Z�e>@<>�ɋ��<=�TQ�O�lEH���G����S�L�̪��t�C����c*��v�͸xLHo��_������1Ԙ��&�Ri��Q�ǎ����ћ�������D��=i�b�  3 P@ݍ���Us'�� ,N"L�_�+�S�;�w~������}���>'�_�?��Y�|D�U��24��No"��xt�S����(���g��30��������Ͻ{cѹm�-pȊ��-�5/e:{D�<�z��ۡ��Yv]Tn�i�zBF�v�r�_���8�Iz�00 ����+���5'L��Q)RZP:�\W��`�N���m�������(iЍ����]��/��� ����B�f����ɇ�-�`���;�&NRh�U�A�Y"4���l���@�G۰�m�3F>���8��?'�
:2^�}���)
gc�H�ѕbP""](:n{��;�X�{��iP]�˷^J�C6�m�͡��^2W_����2�J�<)������۱F��P0��fe��&�R��(T�/͗�2fj�L��	:��KLCÂ��r	��m�OZ�s�M���������}���=��YI�:L����@zY��;�����a�9��O*C����`�!ˀ_ԡx^�*~�
l>��/�����@U��b�\S����s�P��PS6JC;6�=�L��w�ɠnrQR�0 +��1�e�o栶��M��Kys0bѫ��sI���S�W/�"T�Յ�a_w�Wjza(�"�z��5���e5��/R��\`}��	�D���o�ŋNݟu�hڹYoÜ����( �4���)2�3����Eׁ���r��B)}���ך�Y�^}���� �U�6Xjw��je�v�����������������m/\?�%�˸�y�׽��Lה��=���X.��oB���r���u�̦��vϜ�W7�ZZ��f,(�.��׎�1����R�X�2��W�üĆ�\h������=��¬�{)��d_�X�C��Ǟq��M���'}�6v�H9?.�h���*�q*h�|����ׁdP���9lN�t?8�vUѫ���z�&<�������|�'b�gD�"�����o&��k�j���Zbߑv��n���>�GG5Ɗ�h��*��������I�q��<��z���$���P������Z;E����eD"PBޠ^b�%�d�]D����0� ��3&!���䥉;]�a�u5�"ZW-Q��5���n�\�������_d._6�g�O�m���0#Q�N�|�����q2���*�p�#�Y�q�C7�g{���궖M&;�xL���"�;��-�B�Ӹ&0�ɫ�%�;-KL���4�J)�/hw���1�B�CZt�$��F>9|���љ�U)�݇pc�:�>w��Z�)���N�g�ْ�dˢ���U�*�א�	~@��1"p��4}6���`)�oeZG������/e��׈�g�&��!�8?4��6�$l[�җ{����PL����l�~��+��:)���]�,P�w�����f�~�r��H~m��xrJ��D~˲��A`ъdH��U��'=k�қ���<�r�f�،�LPu��fq��	�٧߲�*�	ac|n.xt��td[�;���X ���X$MV%%�c�����£ې��6p�,������ˁ�N\����.
��x�������ѾI��V�H'od����+���檸�>]�	�fY!��H��7k;(�'�AFH���/mb� �2*7�~���u`#M��*C�Q���ݧ·&�kТ�e�"ܜ�����_`���PP|!f��/*h� Q\g�Szd���N�����uQ�Jץ�$�!�1kH����W��v�'�t��V��tz>�Q��/q��\*ч��T!��H5���G�Xx {�t�(${���������Kq�S�h)�`w>teg+��,KL3��*��a/���F㹯�〥тU���8���A��ݩ���$����5o��Q�ۿ;���i(K1]��n{\-NjPN=�'	Pj���-�)��*��Q�"�̿���,���x#t�|�+���E�Z!�����o8���JPC���
	\�\
����<��7��Zq�:�8I��e"�0w
^$����y���e�+�mr3���}AR��|yX��v�(�qm���X�L�Y����8���r��%*�A�͌��Μvf�� s*�}��~�B�^���z<|*��Q��5�.��E��f�a��d������ȓ��ʿ�B�H{�t�DZ.-�ba��~Α��U����ʳ_Evj>Ұ@6,�巗̢���m�����G��5�\�v�}��.��,��5���ϣr�v\�?�ڐ�%��\=��ֵ�g���ϻz�:��ZF�uLv�W��)��ǁ���u����+c(��8V�>f�̌���,�[��;�p|I��X��gV��;w��E���ѭ[������3a!8��b�l9���@N�����,�q ���|����$�[��K� ��H����U��#����ox�ʤ����3�c��3�����
~{O�h�װ�������#��Ɂ�$;�~��4L$���ZD}o'�=�v�|��xkQ5�`#��w�73Nr��D$��!p����&�*R"!��6%���8G�w��?Jiv�3g�iPz"`.��}����#��|2��%13�*�����Bg��f0��׈��lz�J��͡Ȕ�#��P�!�K��y��g/	�'�Z�u����O7�7��B����ޡ�â���%=�I��Gl5��%��Pg5V,5d��]��F��~e��x5�	��NZ8�w$�>�bG	j H���@[%WbZ�����Wp@�q�`�&v-�y����,� �w��H6�y2�VeřD���7���ʞ�n�Xu!�32\\p�|"��L��d*�c�\g.N�L��� �(��vtT�N)[�<XAQ���C��I�����~��)fS��<��N��K��ha%��aW,��Eˮ�DݸW�E|�[�3��Q1�J�;�j���8ղ���()zet	C�~�@/�ɴ�(zA�"�0�����6n@T�^��:E#E��g�~��3tVG��K�n�+wf=�y�[x�H� ڑ�R%*�+�\�������l������|w�_�b+Bp��\y�]C7��BbM,i��	7�j-(?O��+��3ep�v;��,pG�����5�8�tcz��Ei~n�١E�
�=�()�]�}���T�2k�0��F�;��.*�ci5�7/#���%���6��kc�Š�o�7�2֫pV��<��<^����(8y;֫��?�#s(�INt��
�.����0���
ʾS	:UsI��@��G��6!n������~�Jd�ٶ�CY~��+�a���J8V�
�o�a�!� �@FSA�rj����$��t�{�:�Ӳ�E��Ģ�N����n<1'�Yj��!'6M��D�Cp��g`@0o97f�-)W�tگp/����G#�m&W�z[ѶH��F�Ҙ�kJ��ԫv�r�����;r�Fhla�/Zҡ� :jR@|�c�0�%po�vkFt���O<�������2�����B�9���=��p���N��mm���@SZ����:*��(:$��x9�B���K.ǀ�+�7�0�r�����BVH�ܸ婢�S�3��}"��1G���	FC�I'��vOG�4rߑmR��:�ɹp�]��c[\�0�e�떂���h�"I6��
�k�g�	�,-e�8�8��������㳐�-��I1eSď������H�I�|cW5��ş�8�YǊ�q�q�e"�������G/��n��l �sr��yS{Ĥ�O�^}��Q�jV��,p�q�Of�U��OS�!lp�X�������9��k;N��8�1 l�M���m0G	�P����7�)k1֓�;��"��d��tp9�P���"C�wK�j��fU���֢	�̶!ZG��*��T�[o�23���C�Ա�p�qC�	��5�o�
��8Ռ#_~��n�!X��o������d���k���`�s)��}�������7Q���9>���~�R/%�Ȍ~ڸ��$�Wkl�$������w^����jʅg�d�er����p��S{��z���C��l�}�%v�O��W�G5���1���W������՚B	�T���p���^�F�=�J�:zFip��۳�	�$iPQL�m[�_�i��E:"�b&��P�ߪM"IH27��9P��� ��+s��xՖ4x:��+������oȬ�{�bFc�{��B7A�V��	��{���Þk��"n��E�EFM��sw�����}_����'e��R�'��(�ˉ�K�c�#�U�;�]c�T��􌌀��^���c
	����:��F�
��h�FXŃ�n���B��KTK�>~<��a���;>��K������4犙x&ْ�(�{PĮ����-$�țA�+V������u��!W�\��*�݈�n��j�Mx�MaC���yqN�NRDy5�Mf*��x́A˥y�/k���}�8�/ogd�65Z���VM|�7Lp����O&�E�j��~)I���C�-� ߡ�|V(l�l�����A`�~xq��~�z۵z'ǯY�¿p�~p"Y0pG��|W��۸0�0śj>���do���&'��������v\�zG��j*a�,�e���
R-�r���G��Н�H�i�:��6҅m�P�����7t>��Q>�Sپ+�:��U��m�Q�oeg��V��KvHFj_��:�~@F��N�B���J�}��T���6�1��b��)�;��++����C�!�]��'V��G%��5^�����<�ys�o�,�aI)"�n����	���P¢&H5�JQЮ���w��7W�&�V1���Z�ֺީ�<�'.�����&�"k�� ��H�1���
��X�{�Qm�%_�Q�Rn�)��C,
�J"�O��A.w{(tN}�+/�>�r�|�H�*��Ey|�*��W��Z�3ɚj��6}!�v˜F�ԏ�6y�6co���|��ܷ,]��:4o��9ǉ�.��e�����#s�wٲ��ӣ�艋�ג?d/�?s �P��d��i7걦�!�p'�^=�'�ի�y4 �a�=��Ŝ�<��1r��q�w�Oʉ�ѭ�EF��rhG�toZ�6�:�("�E��s��r����h���8c�R�W�~��gloFbz�sU�렾��_�ߌ�{b�ωͽJ%sЅ���0�H��#SMzOH��j�LD4��e�Kn���O��/���>glV��.8���0�e`c��n��hV\�����P���9D����(���>�r!�P��y�.~Uhw��C�R�^Š�)0��.�IU���}> .0q�>�*�&l1�a9�%=�2���d����7K�aW���z^��1@�
�Jh�$Ύ:�|���b�,A�U�ٹ���+�	q*߉/�c�2���l��0����t���XW��nx���� �vN]PC\P#tu8
�R��N����T��&��^H�t?�qW�?%Rvdtj<�MNϸ�M����_͏əB0��`����%��Z��=�ަ	��Q��~��"�Ve�I��������3���1I�v�T���톘�ni��5�_�ȁ�(Id�0-a�h�+f��C�C�D�:���O�/�P�������s��{w8�Xqo���62!f��)a]��[�9ʥVTE5�u">�DN��`Α%�`1��w��� �P>k�-O6b �gRM���>闲5��y��V�X��[����Q݋wPJ�� !��Qq�y9.P*�˒���0��tZ5�T�0)���7�n�0�A��/������| ��m�E��f*Uҧ�$~g��ۉ�����-��t�c84�'O�L�I�q��)�=�Vr���C`��t�G_E�I��[�f-t%g0�M�����/�[�r�xn^�kdK
$��[��E&.ʇ��d)C{��PC����� ɣj�gԍa���Y���Nw+��<y���Nm���0��VNґ�S�;A��8�C���P�_��1�Ϥ��*u��b�^�b))�셎v�d[�c��QXI�{w��h\�'�\��M#�6�e�;Z�B�!�H�ri7js����|J`�V�]���d�,=g�f0�JB7��U���V��+������>�r\7As����ڽ1`�+�l���Iߗ̤Z{�7cŨ@�!�����@K�;��J6_��n���2P(�o��N�9;�!|<Ԋ$1������YL��o�0} d�H�VE��&u�<W��Yʺ�2�aq��h��R��j�3+sZ)��؎wYT�������E&,C[�D3<F>'��|��;��ʸ���*���k���ad��~��:�4�+���W���o-H��xi�XCq$P-����c������`�2OR!
��g�������A�+\�� xϮ�y�h�C�i���բD�N�(P `�󖔥��ï �־�h� ��RѩNrXb��r)�f�8�+1�Zȝ��b�S�%�%����]b�ۼ�y���C��m*����%��8�"��M��}�&�Z�8�2��)��P�Gk�=UB�"!\�M�)����?��%C�a$�o}3���pC
d{E�(ﭥ���Id���TϠҦ4 '�F�wz��"�J�&F:N��Xw�u�]�8�N0f_�7@aA�9ꧠ)˭����Uk:H���tϑj+,�<A[5i_�����)�>Z�!_��K2#Y��@,i%kk��]�uxo�(�N��Ɔ�"��8��Awey}#t�ea�mX�!�!$K�	�
��������������ʃOWQ�%�q��#h�8A�h���]QY�M�:��H�՞��u�Y���UQ�������h�q�s��e`Z��c̪�W�շل����!�g#���'_5"u�xF��2+��pr�N�	��K�֎-@h�k��b��\N\x��׮�2����p��4U���t�y7~��9��֭
7V�L��D�>wQV��b�%o�$�;Ug�2A��0b�ՑPX���n�����kP����X}�c�nD�����n������z�G��l�o���*��ܒ���y�z?(di(?�8$��;'3�ʹ�)ym�
[$��Й|��}��^QW�y2�X�Bɡ�gYR����&>c�qxJ3%��û���uB5#&���i��<�0��k9���Gs؝E,�G+0���O�$�Q�O%���.Z��ۍ�m�W}�m�V>��I<%E���!`ŬAx��:q֤��4�޹�yo+�����A0����r1�3�x�6�^<|�ܐ�xFu�j�$s�̆����'e�VĲ� �)4��	Iw���Fzf$S��aMID,�֋_���Cq$�S��g~�ʞV s�˲�V�<�%
��z?�������e�~IqA��)�*�M�U�w~�]�ywIPm�1&��F�"xG��0�oÑ8�§w�pDq%�9/0���ꎁUr/�~Թ�8�� �_հ� ø�����	�������`��B?�U�N�=��������2X� �P@M�&�����C4�(÷~�DϜ.s�h���a_��sH+[���z{d�eO�)h�o�!h�����~R��X�jh�&���yrwɿ�Z��~	y]�y���ђ[��*s*}�a\��!0�5P.���fy��\�I����M��D�n��E�et��L�BCٻ���%}lm ɉ3^��BP:m]bSKBv h��[{�4�<��9���;��:�V%M��E�L#�e��)2�'^#���V-\S�=�M%��7���I6�1@�����c6�$�"�1Ccj-�	C���A�?){h�v#VG���h�j`�c'E��c:]�A��M�@w*m9����D6GO���z�
��P�r��2R':Ń�u`Β� /��g���y�Dw�,L<��ppP��vS��۾[>��@�&���3��.7�X�uJ�/E��<?�qțD�~����V��:UϽ���[� ~c�ԙ���ޓp�z����Y�����f2ڊ&r�z�4s=�g��R�m$2�C��)sWՑ��f����@=�
��r[���ݡ$4�b�Cb�岫d\�����y����{=n�Dp:�w����D�ޢޚ�0��bz�q����N�;��["�׫hŊ����$�˴*�Fь@���Ց��*�$y��=1��5:1 �����R��O�.�}�x>�6kQ����Bp��)�@h���#��vѭIi��y�e���j<ʟ+�j�Wic}��Ҍ�{'��E@�u5���o(��Y�����I��cUp���]�WE-���$�~h�
z���5�\�������x�ۭ&:5�ǀ:+�����p�����j�.۬'i៺7_��w���ő���HZ�����L�gm�F��\	��w�_u�p��&nB{\�|ğbj�T)$�E��T9�,�s�3%�f|��s^tػ���K��ri���H�(Td�}��E2���n���� "i��R��4�߶�W��zu2��e��E�������m��q�f���W6���/a����:�ٰ�[�=/��������JC��3|����''��&���:�"obݖ����֬��͖!� $���Fv-D�v~Ъ>��h�27BXh���^����E����V�xQ��@�BL�uxs* 1;H�9�g��/���je�/�S�?%������g�ņG Bj���8k�Ckh3#�z'�5T.�5��Ts�����;9� Mm)!�3��&|d�,�k��ILK���@9���%�4ד)?�B��!W~"���t~���?@���o�b5U2rӈ���/ �����9��=�u03)��1�����(Z��	��>���| �ڌ���-�4�����}n�H,y~�~$q��������ƞ��Y"�0[��`�S^IŊX���/�k���E�[.��3/^�-�h���S�X/�|5;��pm��6�+��h�E���$��"�X5�I��1H�l�a�`)qc��^���9��pBl�D���}ڦ�w"��c�Kٖ���y���	��/��Ā&�m�k�>WxW����ʲ�{�z�nK;��'g�x��T�=�w7�.0Č����� q$�q>O0����ǫ��,�Y.��@����{�e!
"JD��Ό�S;j�'�Z�X�oP�;W׻�A�B�Ϊ��rI�r�����?�L����k܄�N蹮i%D\H�ґ��j�����K��u-S���R�#�Vp%?Qۅ͡e���=�~�����Rp�Z��~�V��ꇹp}�"6��bI��D^]xȨ�-P����Л�$��M�7/Ŏͪ{W�!4�HX=W�ځөj��,��k��;-�Rf�# B���8k�Ʋ8��b?M�$�a�򆌢��N��V��f�"����[SL�M�(��F�or��@%�A�_��d��R4��(����`Ŕ|l�I=���4�bwz�~�ЃP��tڗ$[/�~ k����iJ�A