��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d���麍�Ks�%$����+d7��/��������ߔ,���<�E�]��&��z>��>�X�����k�0
��F��p�J,:�D|$�'T*6��v,ֳ`�7J e$���Rv��QL���M'm�l���e��d%����U���Fh�2yRp�.}`˩HD�c
j`͔Dr��6�;F�c����:������xصV����2MGބ2��/7i�RV�	4�[�-- p��Q栳��U��Bm��}=t;�cL�Y��e��s;�)�u�5`b�mN���A�ڻ�R�[
 ;��VK2�"|�S,�b�Q�U����:�*8`��~���F�c�@I�{]�~�����w���uFg�<�Zk�a~\��c�ͺL��)#��JpJ��a�tO�b�2�U1ў�Õ�9��SΗ�M�~�u)�n��%]�9��z�E%c���_���]�C���*��h��.���}��5�7,&��`�iQ�E:5���
1E�@*s�z�` Pr�>��NEl�{�%Oz�{���G_��+ǒ=�V�\?�7�Z��<A�]4��cg.�"��EVk�*X�H��w���S�H�վ�M׭W6�RSCT0��+�eJ�{ny��")����.Ps;�DEJ]͠����e�\��@�k�Ki/��n�;��A�`����xa�c���g���,����d�!�߁,����͇����֖U�pC��@�K��v�g��+��dCS�^�(�qLے���6́����cSɹ�|���B�Omy��98zj{�&栰k!���Q�Bɷeǣ���ի:��9b�!dO� �$*	��\����,�7�IQ&�T��v���R)�a��5��ݬ�?��~}iS͎`C�O�Ǭ�>��	���s{Q�}��8j��#�=aBѲ���ՇB.g�@J9Tᅾ��PZ5�:�t�y��:~��$ �)�P4 !�N�C�j{+	�c�x��͌`�{f�"�|L�D�k�Ԝ$���A�)D�L�y�� b��Ɩ	�r����:O�ӑ�[�b��L���Yh�5��z�8����b����Ƭ�Z��T����`뵺#�ƍ��Z���]m�ʞ���+���ߍ=�º�X�����ˣoR9�<qMt�Hf�|���rꝽ~�usꋀ~���z0��a�'# c`.�C�_9����bi�t�yӥ5�K�R�zV-�|���\�V|c�*�hw�̘fnwxI���C�����7��~i��N��Pd2��c��x�{��+������7i+�L��󤼠�&�G��U�.�E��9:ˊ��ۼF������d�|\̢�l���������y�N���T��L�+坟Q>�`'�@�2��j���^=P�����N����tlMn�����.���[��F���:x 81Z}1F�%�;��3hIE�C8dԳ�=��5 ų��Tʊ��F����#V��"��'��(ˢ�����E�Y��&������}X:��qǾw�}��d1��ɱ.����釾Py����U�Z�0U�1�Ӕty�>�I;
¯����(�}cM?l���bx�� .ڮ
�a�x7d;��+���.�f��
�7��k�|��my�^��[iǻ&���2��2�C��.73s2�{W{�K�h�����pl�o�$�QR���޶�D_ؽǄ�_���4L?���"�R+��G]+�Bf�{o�F��*�L�˨��<�7�'.��+"�vφ��ʵ� ��A��PF�v��b�-.��%]��摹��%$e�B.ޓp�{�	����vM1ya��V8�{�hy�0U�h��|kk/i�V����ڌXJ�7���$�F�5�"5m��V~�3(>�o/Q+dM�������`L�n�9�����L�����s�T怛5�#����-��t��3D��S�kvh)�MA�S�Y�BR���$��È�&�`w�&�c��B���6���7[K���+@@4�d�M4�{H}�����pumG�ۍ�O�5D;���W�@�b��:i��]8^J�Ɓe�H��,���}���zp�����q�Kf��x�����8Wx?^?��X�b��Տe;��	 �S����O�R�v�"�%)�Y 2��Gc\�i�����R��cs{X��B4�#q�z�JC����;��/��A�Mv��csJꏥ����m�,�Ό�P\z:W���7O�U�Y���<��#mB�S!�Y7�o�S3_�H50{��0x߸���$!L�>^ �X��%ti��=s��x����������7���?��,DCM��r!��B9w�$�23QQ;�W�'-c���ji��,i`�)��\� ���"��~�����3������:�>X�����.�Wg+�HzL
��ʮy4�P���4�b�n�nĚ�d�-K���g�q\[@�AW*�rKJfw�7�_���jsA����	ގD�꽣䮥�~������M^�T%�����A	���$����R����Q�
c��?N�۪_ 0����7�/��=����S��*����%���(w��k\�w�\� #{G��Jl8R���r��S\˞4ܕ(��E��Ll�ьXV}Y J˘4��P@|?:�!�����L�ȍ*�k�VQ�+j��@��B��;G�"D��!o�FҠ=��(���f�叜C����_�=U�?V+O����u��ѧ��Ӵv��+�-L^�6κ+�<I�`�>7l���Y�|��ϟ#K&2�u\-[@�忭�� HӍ^-�61�	�M���$Ec�=O��_ӥYb'��o�ڕtO�uuę�y%����lG#�e7���ԇ=rC2�=8g9G+u;�<�)�?����po�XEA#z��vA;D3Cp��|Rԫ��]<S�nA�:��46����jh�B�Ơ Ѷ;���#�o��t�����'{�Z�A^a�9���"�#w3��^�D$Y�?x��j-'�ֶ�5X݆�}x�l\�G1��IR("��O��pW�c6X@�e%�cR,%������hL�)G=�zS3�ʨ���#�Wef2��w������	"q 0v/pnE�M, �9K��Wh�KAR/��s�sG�ų&q�Nh֙l��b�|��1���\�4��T�u�s���Y,{�,�0�G�иs�xD�R�����D�.h�D�F�$��+7�N���3n�l�:�]G�9.x����=E�n�ǿ3��U�A0Sd����=��J4��'��I���Ϊˆ`o�� 5ņ�I&�[�����`�z����M� n*��x��]a�6�x� ��>ڼ�'@{R�c�5N���{�q�{ST�K��z��<:ԕ:ݻ�#z�i1;��{6�u�S�Dc�
a��$�N�����_um '+���uW(�3l�)Yfȹ$M�w'cS�U��g�qXד�r.�>J���y2�c+��ByC�,|���=*��,�,�HF�#*2d�z�N��<~Α����0!��dĘ��[}X2��[�쩕�ԩ�9�N�g�A���a�q]��1.�FEy��|�A����jsت�	�a���Ma���aL���M�5&{�+c��=4D�c\P��083N� Lwt�K���C�E��eoZr|�����	��qF�JHa�Е�R|�}W�0�/���A�g6�u��t+U��Amuo{}��i��Xc�jxL�% ^s4��L�L��9ȿ)�ς��mݝ4�RP[���V��ƫ��+x�%��L��2e��U��gӁ.4������.A�Y�FCD?�v���ii�;R�����ak�{Æ��|| ;N|o�S��g7O��h1N��(�Ԫ<��luĹ�{�MQ�IϚ��E���#�OD3̼k=����N��!f�76��e�8�%܄��)32k�e �)�/W���td�:6F��'�H,����k��5KA�'X�SX��&��b�,7WK=sj2.� ) ԉ���(�֒�X��o�MY�L�
��}x|?IRh�-M�?���O�+��B.,���{�
AN�YY�;���a�2ۤ(5�O7�S�����wV	���*�	k_�����$�^�8+C�D�2���<���0�����-�=,z!(�L,b#�%��d�ڨM.1!W}��O�C�^K�X��Ӫ^�����!�c�J3�ۨ����8��'n������d�{O�{W�'�,��X�2�3��i�C�$
wЄz���i���{�j�p��ǜ�tW�!��܆�o�Z��K@i�'e1���@0I▞(��	i¹��Mג �:� ]i*r-��Q�&�+��ܼ�WX���sU��Q�͋<��\lF�p�[��17� r��]_�3DD��?�7\E.45�n��5���߮*��K�J�f�^ �5rl��(q$#!�\�v?m�U��is��sɶ��-�+�|���3�%Gi�����I[�"��"k�\���f�s��F�p�Y�����K���[���JX�HwX�<	��)��Y��U��5i�! �@y�KɜxN\[Ozq�.;�(�Y�#vP��@M�6�U�%��N��+�`���8��Rko�3��3����X�Z���E�Qӝi�j�G�_���j���X����7��H���_p,�)�,�UE�Ux�$Ax|�4	 ��s�� ���ɪ��&R�λ��敼�����x�����F�w~$����(�����K��[��v�w[2s�m�OR��@�����U,؅����NX���xU�9��`ʐ�a><���猝7����q�P�
��.l�F��m$B^ů=�����L]�	ú2'{�>�nH}���$�O$�F�R�M!!�U����·�z�����2����wQ��f/]gj�m�K�"�em�C{��:���-���j�K!����@i;��ބ�k�<�KV����$s7l�����t
^y������N �e�ї��*V]�_*��lI:T�p
Ĥ��"����i��RT��֏�C��L��y̎v��o�Fy)�(�Hp��Z]�ړS�{wim�A�j��$\M���nկF �1/�"4?�t{��G��]��?L��pJ�U4&�|Uh(�F��dD��7�8�]�>��{����1[v�.���1-#5e�.�1K���
�+D'�ڞHߧ/�Xdw���\�7X���!��Z� �������/w4��<s��փ|�ʳ?�A}���f��-p�g&J
7�9U�c��9�1�'G��9-�!XK7�w'��F�FxoB�B����"�Oa�BR)8�pe}���hBq[��f	Lǩ�N$W	��&��P��v�<�?�TdK�|�s���;��;J�ή�&��*>�J�����I��._�Y��D��e��DD`.�6,	b�6Ǹ�bW��i��Ҋ$�Sq>�Ц,kۣ{�hOi�;����
�HG:;�H�\���[�+R�����9;�"�w>��/��1���h�]e�8ݎ=T'2��+w��c��ő)�D�l1����Y�L��/Lⴻ78@o�I�y����&@I�AMY���GO����Q�6g��~̭,�I���)�%Hҁ������	Q~΍շ��]-<����&�D{C;��cI�|	�m�<o��n{B99��}���6��-�U�J������l{]�� P��@�=��	 �W�9?��f�]Tu�52�ãov,��Yj�Bq@4C�\��8���e1o�i�b����2Ri�-�]���(���ޮ"/ ;�����ː��w�m�:kx2��.�b�a�[��  � jg�b���m�F���W@�'�5%���ij��!U��yg�7��r��&�������:�4�r�tO�Ǯ�|��x
�B�����NX).$N�r�V�h��.7:f��0��p8����r���3b|��\�zX�a2�SV��Q��a�F�V��\л����q����eJ����s�Ga��d$�G�`2��D��~���=����ҘVA^0錷Ս|Q�Ҩ�ݟ��G���\#��*��݅�ɾaIP,-��ô���%E
�g�qB-� ����������j#邩ؿ=6~USY�/��gc�������+!ĞxO�:a)oOv�Ƕ"]ʢ�B��Uh�q��=�d�r��i��@�N͉E�9U}"q���9;��"��3+�X�����v�v��⨺%���"##0x�@噒��."cB��qT�Da�01����a����N*���A��P���l��y��rԴb�J�5��xȵMa{=�"��T�)����o`4�>�����8A�m:uEU�Yy��ѱ�K.dx�Y�34��w]�/b�l��,@��?�Xl[�?q=�y����������!�����,K�09�M���y �>��/X[�y.��P݉$j=�����/|w�vq#r�I�5�T���p����3�ut��Z��lD|������m���xB�g�!&W)�� �>���҇�S�FNK�����"�,]�k����!���9@�v��hە��-���o�2��I]>]xY�U�e�*��iҍ�Q�$ܭ��!C�E�ƈ�jwC��I����b��@�
��w�g���`.촩A��癫��(o���91?��JJ��*���(X�#���i�Vߊ|u�m��1�{6B�)+-I\et�v�U�dQ`�3��_X�Ky|���4�W�;��ß5�M�k0wn�rB��,ď��3�lD�7u����16��z��Ɲ+o�[��'m��rMVW��8��%x��ֵ%W�%�/V��h�74�`�qo��g����Vr�ղ��y�BC���G�	]k^k���6�j�0	���M%���U�l���mn]@�hK6I\�]1e��P;�]�O��*~�(I��uz�¢�%�!��m���@��rA��>sQg�A���:f�|�g�	o��i��3X{�tE\F����������ٻ��;�B|K�5l�"�[34��D}�;d��:+X!�@S��zh�ڿ��_3�;�Vu��5�*�?�o�/��+3�Pt
���)\���/Ї(@'�4)�n:*g6��ۧ��qR]�Լ�[9NӥR���S����^�J�؊��	j��h>��u��;���c����	5o�7����.�a������y�]Vb���a�?.��2S�'|���|{���4�İ�V"����E�G�0��aܢ"s������ �:�9,<������^�qP$�oёf�S3�~����`��ǘzZ��0��<�K��9��)� ���T�Q�tNu������^
�"g>��2�ǎ@	H`��#]�b�$�q��fE����`�1<��T�)K��W[�� �e��%(F��x��hb$*��6�I0Z$�����P&�y�q���9��ode^�G8�I_��/V�<+B��j�Jfs��+��b�z�Ev��h��J�uH^���%KA����tV��I�c�q����g��P����l��/۹:�-pY^���L�J^*0�b�|�T�ʵ�ԙ�2���^��_4 ��?�'>W�.i��5l³���Ly|��0���B0j��%��#{��H��Kf�c��%*��:��K���Ѓ]$�=Y[�=Q�ʓ��������vz*�G`q��<���H�qc)��G4��o�M�'*�zC2�"�>�h�ؾ��w�&G?�ַO}�f×�d�݇��i�ZZ�&s�v|q	����F���[g֏0���Sռ�?�8�*�R@�hW���]��	3�|�p�̨�.����$^�`LX�+Y��35�)�P�?i]vҨn���_��,iJч%��8f���e	}��a(9`�<rm<M�.t�x#h��p�ol���]��\�\���>��d��^������8�úi�[TC1�O�e
�1.�#rױ+<�)�ER�)nr�^�l�6Q�=��&n,�8�wV�@eect*>ծ�"!NO/�EDщ��Ĩ�����5Oxs�(�o���[^zY#S���r�;Z��R!��Q�e(���~�$xD�}�b{f�%\E�يa�Ϣ��Q'���6Xi�c��G�|�rR%'�O"HT��ᇐ�N�@ 'TNE����r~����eӊ������T��h��FA��V��70�]�w���"�C������K���7���o�_|t�e
�`��s$2ܐ2��nm���;�AȂ���a��|�&�eX4ź6c�U]~��:�	>��� �e��~��s��{o�����\���S�x0��%(7�d��Qx�;�^pk��}�̚�6@�m���_k���.�
ڑ�o�Ƚ�7F�ή�@2�G����o9�j�=��ܑ��3����oq3s*&ҧ�ah�u�lq,��|>J:y!H5CG^��}oRԷȱ�ɢ�v���t!/e`��z�b�D���^��O&A�olc�7�mJO��-��X���V����<S�S���[�$��� ׾,�**�����.������ zV�����[����3�Z0Һ���nZ���x>�Ԟ ؽL�|�3� ����z7���f�����ɧ��=@��7�V ק�E���ÚJ/�(��(��|CX�M���PW�w7:P5����Ϙ"�J���o��_J5�{���q�а5���ν����n(�=�w`�O�/�%�LS1�Q�Y�q�n%��W�pG�*�����M��}�Q��qԏ��B\�`���3SO�g$�tN��%?�R���Y�	���bbҩ_�>�R��:�� �n��za�R��<��'7��{��i����W�,օH��XU؊�1�~z\ƙ7٥8a�s���kw�VtBy	a-�e=Sb��;�����=�����͓~�E���@a�y�D
M��2���&ߕ����pI�|$c�@��_�fg�~�n�i+s��)��r����W��}�N�~�A��e�_��9m�����4������^�A�W��y�{�����q$r����s�J.4�B��<��0ՙɍ���X4:?�&�+���Z_����G��Y�c�&P���?TU��|a��Y����Q�MA����]�]5�]��~(<�"V��td�PRq8V'�� u����e��i`�p	eV�\�=tN���}"�3���]lӆ�4CQaZ�Aj�Y4��:���F�ͧ�|6������d�9.ټ�C[���F�<'�C	I3�o���bg��PZ�C}KW�(�@�@��h���s�x��FV]��43�]��?}+�+��Y��kQ�^�ܔ�{�BfϮm��;�ܫK���NA�x�������a�:�z���v<��e�u�R�{H���md;���k��/�$it�[�M�x�|IOz%����jģS��g�Ѭ���{�!^n���X�0hLZ��d;W����J��^r3wtf�Q�p�H	Z�*���5� �ۭy�PBM�L�R^�s�%lT��c�7#n���h�E2��������ST���,U����8��q'����'r*W�E��D4���(Mcj5E����~$���a����ߒ�@�n��2����n��}�p�R�_����1'p2Є���x�����EP�顕�q��j2X�Νf�hN�����n��1�(+a�`K�VRĿ�i�g!��
��GR�q��F�؇(��xc�@��k��˕A�yI�끷��+SE��������n��R����"�OV�t��(�%�}W'݇"�WB�fG�8��a�;Tg-[��L����s���AnD�rh�[v��ͅG��(��&�0�(X��t�b�����>=�)�+��1VL�Z�R����^�!�v�Q��E��?�'6&�`���cI%��]���ꜰw�+ۏ4>]��T��؉WW�O�;Eu���O�mp��O���p�bS�N�k/VPp���|cz��io�߼�^���1/b
���b{R�_̳���p��}�Z`�r�p��hfvpYr*��t8!�1=;�!	�oo��
fo\D"M�!>����#��>�����j7D��0c5xV֫5x�6aE���D2n�3����[^E����)� �w��Sf#��C^�YN� �j�laP1(Ck����.f��G��놄3J�L@긣�;;�����(VN����7M���m�"���9�i[��ɹ��c���( �K|ѶMj&�;��������Q�
1�nZ����[t9>)6����8�_ye5&�9|�s�����.
Q������+��Z�o�ͫ�d�,boO�䫆��P�Cw�ڿ'H��ɇ�P����x-�Y[�󐌊�'y�*�[���r��T�|3�ⓥ��-��2sӲ�����(`Z��$N+�O��B�@+?�i��m$�0J�:�Qag56hS� ;��R�9),����+R;�`ap}��~���y�x;=2��߹�2$T�\i�_��E������~����n��D~�7��Ko�$H.��Vq�L�F�Zz�H�Ӫkot�9"W�ɫ����޽������Qk����� ����?��1Z̅%Z�겜%��Դ-{�y{�1%�Y7[y�^k����^�;�$�Q�����W���&Fa��#��B��{M�N3���zV�&�;*�h��%���;h�4�%׎K)Pj��v'��z��+,��3�B�u�t}@i�)} �.eR�;u2��6�}c�q�?�����=�$���{N̯��%
É*�}T���\sӓ��׵!~���\����/o �����%'	��K5�fC�d���ު��%Y:���prz��FL�$#�o�O�����=!�FΫ)O��^�΍�w��zmu�0�vc�|,�q�P�[���5SZ�����J��h0��|$�yD9�@;�������!,v����ih%��~�2jC])	�P��Q{��'Bہ�Y�ӈ�ʈ����u��j6K�j���+%�#2�3q�ɔ6�<A���T
 +��]���eǏLz,��
����g0�@�[!d��li6�S�y�OF�"�X�&�ٔjF\A��N ���=�����)ҷ\Ν��w�m]3cl>Zb̠��4)Z�'pL��BI�=[���}�Y�~�K1N��_%^K� �O�4�(F���t�(3ߠ4��[�E�/k����Ғ��PVV+�5v�Wk�<k��Fi�䗎˅t|���(�8������*���i�Uq��E�B��<�$�e��%�-7�s+H<}ILV��y�㶯ԾyH��!S�U�@�Gc\�3/��;x�S]�?�nS�}K��M	\!d�g,���PX?+��'ՓW�⨵;��)�����H���z!�@pJ(3Y`8�37���l��oG���-&�
���*�7)��\"S��A�� �,��� b���W-�YSJ*�{�����X�b���&��>���4E]2�	�U��y�ZU7�yz���'{d~���ơ��#�;�I��52ER�´�aNohĲ�&���t�8�.y�����٘�<)�VW���#y
��� ;���\��iџ�X��?G@ZG%/��Tq�:{g�)�PYJ|���"��ޣ.7P��>l�+��`g��֋�~׹�Ǿv��^��t��|�)"�gV�x�rX��N���kX����Ɛ�S���/�v ��բ(t���Y �w[d��2LY��S�Xiw�f�����a���fU����W�|\!P?���}X��[�;_a7��������&��9�Z\;r�G�7��ɾ��x/�j�C �F�-Awd{��2a-�7�p^1Ƽ��m�2|�=B�S�|ೢ���*�Ȋ��Ә?��w�6cNM�4�	�h�0�C7͉��P�	ґy{~�֋2�(?J�O�vl0��,���p��<W�
�I��e:_H��/�ꓵ�%%; B����0�+��\���R����@C%��Cbc��a憗�Q�f��������]����FC/��S����L{ܿS%�UP[��=�:BFe^*�q���!p�;U1� ��ɾ��V� w��T�F��|� 	G^��0�&�܎	k��NGT��$�\A��`�ʊ�-g���A�?���5�}���)�Ƿ�vz���׺FΑ� �.��K$�',rUb���y��s4�R�"B��ko�1�I5�Q�م(7Ғnԯ�s(�a��)�d���c|_r�:w�Ɋ�|����`����6S�&-�H��z���0`+�U�q�}�%����%��2h��y*S,��8Bw_�"]h��Aea��H�D��\�/|������l�����573�D��2��x�Ce�*�(NV������gE�`ܒ߇2�`/+�ٗ�f������Q��t��)б ���R���b��c' �E�<�۪:��|Y�����Z�xOy�p<�!3�S%G�4P���V�d�[+��0��Gkq����<Tm�|s�dF���Q���+��:&ӹZI5Rj�Qu���6ޝL|Ǖ~��N�qlU���Lo�o =-�u`���������������j��e� �����6gzi�qX��ږ��5����o�C-V�rB�����qi| Q_Y/��L�.�A�Ip��'��A�NR^�	W�A'W��PЏ�����f��o �������� p]�$��剩�b�g+�ǆ'�Qe73a����r����_dÏΆ��S{��4
B��%Bk�n��]C̬-�_o*\Lk�m��a;��v:��"8�d��a�`��ճG�U�#Yr`U���2JB��nβ����<˪w.Z`�F
���+� re�w�$�0I��@K�"ٜ��`�7K��F�֘���hq��g����D�y��,���7���4)d0W˹�����D�x��t�����͹Ft�
�7�H�%=��YV[���������Q�YC7���(e�@� �>���L�{ Fդ�X�bH����r�g�r�*b����⫖B�����y�s����Y���T$�H�2�R��S5�����@3S�� =qZ�R�1o7��&��,�!A�NJ\���jZ0���G�W���FIO����/q�l��C������ �M%��bqQg*��Ng	&�������$0O��u���2\IJiɶ\Y^n�K�ƾ�Q��Ӕ�7RwI��D�#г��?R)R�L�E�ꑳ�z{^���zc� �s�xX5���`��C��<w�!H�%���:���gW��Cs�Y�}�?;���l�ld�_)�.��#Isn��j�`s�>њ^L�b�t���y)�����Ȏ��{�ч���%����EM:�����n��) ٘�h�V��8c����r)�|����!����1\���ҁ��<}�8
CX�q�F	�-�yn�rEȄ�$A�@o'$�M�΋!;�{�ij��v���э�b�s��й�\���x�Pƺ�,s���XԽ��^
�e�Sģ@�vX[o�߅CG����^����A��%]�?���K��U�Mvm:)x�n]��n�4�P�D��<��q�{׸�{��Z �8Z��e��cfS�������Q���Vt����fY��9:X��N��z����LQ?�R�?�9�f�F�z����q��O����<�XM��L�H�t�����������"e��>a�R��-�sf���1�.%� �-���V�-��D�'x����w��O_a|��M�^z�򵑲r��ҏ ��,3������vX��z�8F���\V�J��Z��^����~|�k��� l
�_���r�5i����!��W7`�%���)b��S��z�C�7$qUB A0_�<TX�٠B����o� lw:��{���_'�Z<�M: ��$"@����R��oOB� H�D�`��FD�41sͳ�+g�O�Tق	��A�3�a��fM�0�!���㤬����o5����1�z���l����:Ba�,_t~Xд�%_��4�ۜ����]!��+�%�A�`'�1��"��Z���Q�[^Z՗���L�i��+%E��L���J��-� *����Y5�bn�>�b�8�V�Vܰ������ ��i@�ʯ�O��C�D�+�&�hp���j������˗1K��á�+D"S�3X��a��5{�I���̟��%矼`�ˇ�Nq����_��w�K��X��6�p��^�su����Ƣw,�P;.oqz�E����}:���3/A �b���VڑNT��SPb�E9��G���UT��|L:�d��u��!���ꎑ���n��5��� ���2��9Q �u��#c&/c��ƪ���0+����o�.u����}�w�o�Y�X_��qd ���R`��T��j�׺H���&�+�R�Α�s�����
,��˭���H�b�u��2W����u�+qV}�dE!�y���["E[�ޫ8�h�ez7]!q&�4çd�oj�^���X�K<��zmRc�U�͗B�l:���GO*w�,쪐��)́��qC  ���V���Wf���(�Q�"��UXq,��}D��	Ç��&}=���p���h����/��P��z@a����� �0�UW}����[3D��a$��������v��W�Gיr��@;�q��P��.�f���~�P���������I'k�=�T7"��&h�7�N��A����n	i��l����.x�>g^^&��Z��pђ ��3�tH���Y\���KN�b/������������MHWj	���G-4�e@�XS�!�����Z�;;�|��
+sg ��^:� �u�Ì��8�=��غJr�֥$�OnE��ܩ�di�d@E�E��M��T⯈��q%8��S�40�_!�\u���`���xU������$6�{��'h$ު}��y�l��1%��Z�ڠD���3��<6��)C5�m.��?u�s�K�N�2�^z�.8ɧ��~�#](�@K�"�vB4��e���z��.L��	������M7U�����P�G����[�s���o�L�oj=H=u��tr��d3v�0����Hfh�.j4��b�6p��Ä]�D��>t��SV�ڈj����3<�"*��s�)�V�|��;�[�) �� ��_|�Nv���n�ެ+K�T��D*�j�?�YuS��67�jF|�K����:j�6��!�'��H�Mk�vgK�����\-��J��*�5:�99=<�G��Ϭ��)���B@�-$T�D�o�%���
I�|=�d�{��VCGA�g V���?�n�w��$ޛ���ڦ�_.K��!QǷ�j�N�m�����?�z�nYN����-毳���"�|i��fᮧc�+��	�]&���_�PH\�h/O���H ky��w;q�u�'�3�����w�#�����4b�T��	�?����]v�Sz��(.)�mz\�ҳw�.��5J`_��Ĵ�y+r�R:p'���A��WonHh]��i��t�!C�ŭxj�6	u"����NV�[|�������2PM\���q��O}J1V�/;1D-oN��Vu�}̒��"m�����Y�5�И�˺oa�4�]�ֳc�; �{�L��5F}�a���Y|m��*�cL@w�ܒ����|s���M{#��a!�H5�g^�\��w��?x�1��yC�Ze��cm�q��M���#�.�%����bZط@����Ij;S��|ѿ� ��K�����$�tģ^,k�Xa����ѐ�O��?\|#;�6�H�<,��&�Y2�� ��j�Τu}k����B>& _�뤹s���Ó��z�u42�?�l+���-��� �	ZI�-���L(6B���o��PQx�T� B6�� ���ev��!{]s܇)�dn�8P��9�'���ֱ�d�� �i��K`5>$�=ؑ�F�^�m�mZ8?��<�K�x���5Fk�#��R���I,��YM�<B���47�<@�>��)�YYw��[�Jk�ן�7�@�s���4,@��U��oMl�u}X��V�&��g��[��Gh�.�z�I����A�A�4"7b>Q�`L��-��d��w+���-��gce���e��:#�z��F�Q�{���54`����t��6Om�ۖА�
1��z{"�t�	���]��7��P�����U��?�0�W�G��)����=$�|.ή2�~�g��W��/y����Z�'�$m�K�B�۵�.�2�r��!����iv�Fc5	��?��*����+��ԅ�~��_����@�:�A���,z
dH����53���G���v��Ec,��j�Rn�"\�xhF�8p<&��Á�|���4�Q+��_�a�&{��˱�^�
���
����j-.�B�	�i�j<w*��u�u}|��<x�X�n�~D�Q�T���:Z�Y��-qH6Vݬ_8a�5�c�Wެ�#�
W�����^����W�S�["� ӂ�2jE�O����n�H,���^\�]Q쓧�{a��`Y��$�4�Dw)[���� t���b�q���zs<�i�_�!%eՃP��$�}"d��\�O��5B�q��N�L����&4��k��I?��J���w3H�}��j�P"��cN�����7%������}��}Ɍ�;����k�o,��A -�<��Ԅt��`Y�Km���&���O>�L9\H��L�����Nt�H�������p�<~�ӱA:7y���9���k��o��Ζ,N5&�Txz�`��ߐ4�/; ���f�� �(u�D�T�>�5��2�CK��"@�T�{pI	�q��IT��d�Gt���1y�x'�w�{�~��H��'��L�Q��{r���Un����*0�@)h��qkҀ�WRw�ψ�~U&�R�K��q ����~�/3�GP�/�!��e=5Jʖ1XQ�r�%^�g�!�;DP�@�[Q�HH�	Ǡ�T���@_�ó
��c��'�a��fƖL�:��%`+Ӱ�:�� ��G�(���l�B'&NKx �΃T�����K�	�52��J�rp'�ZrFs՜���]g�އ�WSz^ Nc����g�����xeꊯ�j����s�_ό�f��9��[D�1�cX~��X�x�v��(��B���@�>��Q��q���1�(h�U�JPˤ�(�g%�J�����pY��禮ǣ�E��t'o>��~��H�b�F��^R�����m�~�葺���AH��|�4�{�w°PT�}��媿A�^�}}���m5�;��`H+�=����Z�~&(���c'��='�^�u�UV5��qOޞm�pu�1X�¸7osd�)i�r��Re�|��S���
r�Y͕5c�-Կv��ch�X�G��|-!��#���o���x�Oj�׵vt��:��rh����j����o �3u'�^�]���10�7&�X�N#���D��f�t��QlޒN�;fo.���o�7Lߎ�3�9��o�oJo_a����v]�֪�B��̓2���
'��14��jy���䜜$X���别��DC���	ט}��O؞t�?�F�~�������,%4����� Y��s���k1>Ij�G���|�գ���w�Z�(���z;�����4���І�B:}�Fp,�LEs�-�Sb��;cfLGvr_���v"o�Ei�PU����3GV���������0�7�����s��2�O@�5���Z���ӠϙU�ѫZc����"�8z�W��ſf��
�v�����ЛC�=��9�L�5mD!��:�Q5+�@$�D�1ҍV�8�I�V�bW^bigj6�(�c���$\L�դ��ETJ*l� �vXfM�;�����#Ge�
G������V�离d�xC���,a^s:��w��e�0���w�Z�_�&�f����^�u�N��O�3�x�MV�������Y?��Xh_��)B���x/B~?�U�d�
��{���T?��o!-�gKf_axFq7�҈7�>�8g�����-��� pN�o[_ب加�dM[{�P�(:;_2�$�d3�Y�o�+]U���0E�[e*���[3б�j�vV_��Ěc�n�����ud�޿�.�!|���WO�$��U�`��@_������ ז(E��#���l+�Od��ɫ)��- �Ԓ��e}�X�z͎�"WNr�^ܵ������@�޿�3Z�%�j q�*Fs�]�E�1�����6v,H���4Jx�<ۗ����J]C��hϸ#�aE:���To�&{~��)v�����_��nN�92l�u>���;�v���5\s�y��f��ƛ[�֝�����M0�VWk���q���?���\�����
�e���ߔyɃ�n*.%�㐄����J5�.G3�}��([hj=��wh���I��!e�{"̻��4&E�x��i��F�ϱZ��u˔��wh_>S<�(���x'�Z����G��iyӽZ���ם�eϺs (	�2ec+k�����xEb�v�,4�~"HWd�Ҙk�T5K#̾�Z7���zo	G�G��^�_����� 69I�Fӏ��:�J�[1 y|DMU��R&k;S��c��>*[�g�s���8�0֮h�JIp1U����u�N%	W?�&�O��H�E����C�8v���'����ۖ�Km�m-͕�=�xL`�=��	+�����$q]0���&������.
�W����U�F�541�ŗ|e��_�)�6�)<���8<"CB����N���-�[���S4�pa�[L���жNA��̚�O���ˬ�C�Q9�P�]���qx��`N��E5���й$������jó�V��~]צ��TՓ[��ao�$'�|0���؉���*e� �.�v��"�CT� P 2���k폳����x'�3/I�9�5�:�݂���g��4�X$FyU���E�U��6�Yz�i#Z��^��\�u�D'�V��d�6�/�)R<�~^1�ox��	D�~���Ϣ�E���U��"�!'9u�$p�� )n�|U�';Ǖ� �b�o�[t��^��չڟx
=Hb`�%���i����6Q*����Y�2j�ѕ?��
>��߲�_ddq�?)��\��|��� ;�.oh'Q� }�Xw�(�?�|�ݗ��S�����;Y�$��Hg�˝h��m ����	��엎_��C��o�}���x�qA��jdr���hVX�`m��X���op�c�2
�*�A�-����>@�ȼS.<'�:j��~_��<���S������,0K�_ӝ W�����&�09#�7}��n�)�xu���x�vy�(�+���4�l#oFβ�#�`��ܽ���jl�,]b��KE���cz��r�vtK��
��r	��ԗ��\+����Q'�o9Zy?�YO�@;��|m>��$��KO�:�.� ��L�~��L��ܯV1p=�6�Ş`rm�o��2D���"���
Ԝ�wݵ��#2M]���c٘MC���]�� FP,t �\���HF���L	(��a�V�W^2���N���7`�PYE��WSw��v׳�s�i�֯p�(}c�{�Y�r���Z����jڋ��߬��0e�D2G�@�O��B���Y}�;��MU�}@"!ET(F[�v|aud�[�, ��ʏ�^搣z\�F��iwg`��҃�K :~�\e��ڷi<x��b�	;�9���A�j��H�aK6�R�Eh%̞WtH�>kp7�;4�S>��پ���w��8ݻ�.G!
��H<��ɺ;����I�*�ԇ|�1�{US3��J�|� ]G���b��9Ͷq#����^~�-�@<�GЏ�*���	���wӯ�E�e����Aƿ�8��},t��(�-���3��W��a� F<��D�y�'�p;�g^�	,E�.��F��Sf�qY����S���v�:5-�OU�Ȩ�=]vE�C��ړ������W]��Ơgn�+�{E�6�XB�;�gqO��gn}#ƅ����M?`��zO��k�n:�#X4�����M3�ռ�ս�[2(��|G��\�[�
��5!2H\X��=�ЈkG�*δD�����JS<{ﲽ�%��a����:�J*,]�7����#�$�#N�!�.v�L�%���Q8����F?_^��l���pF�R��]�t����YE�S����@g0F~��S�E�>���FK�^N�ɏ����#��͕��9���y}յ���T-w�⻝ߗ�:׳�������\��*]��§߯�n�i#�� �7��cH��X�0!_B��Î�8-je�"!��X��>׉�W�p*{*Gߩ�b�z�`){�6���N\u�Ms��v�9+ը����j�?�6B��#�]文FN��3�i�����W���B��d_� ���@�7� �v̚0S����7r��o�-�Lip�]y�_m[�ʼF����D��C�y�*�2Z��1�`XԨ�n)���<�w�H�1�j��0����+�0{�a��E�ϭ�\�ym��Q����ch�`�C�n�����I�w��Xx?���^��4>w#LI�;�\�ot�u�?"�PR����ɮ8ƼW�Uj2�+�;>�߾�z�CPP���80	��[l1T���.�j���ٿӄ�$\�X�6��!����Z<���	�Z����`jQ�o&���p����Ϯ�K�a�M�]1�t&Z4|��Q��[��L^&SyB2�*\S��"�,�Kh��Rnq�}�$-?ӆ�܄#ͨ�\2�{X�M�5�?�D��6հ�V�zif(����iy�����04LP��qZ�v>k��`W���<��^�!����"��=T�6y??Zo��A-�d
'��.�;]+�(����B>�vM�fd�h�m�#�=�����Ю�[��?d���j�i$g�d>Q'�<�H�$-�a� ��9ȣS��'rga=��]�8S;��)��"T*>��֏��s^�:
�R8���e��$Q.�l�0}4oD�D�@ʛFy1.��B��3w���գ�z�r"��(%ǩ�G�
���?��$LcV4~�?�R�Pe�L�������B�T�cy4C������UC劯�νV�.��n�������k^ ��~�VD�XY1�{Z��F�e,�����	�k�qn��w�|�sh�l���_��ʴW�X� 5�feE�Gԙ�K���f�L|`�m�䍪v!����;�2�Y?�r� ��<��'qJ�iR��z_�X#�-U�kf����0gUa�)߃�?�l��r���]�&��8��g���9�%�2A�S��~~���/��`Ś�*�����3���J��Qr��$���u|�C"����M�6��r�T�9@2ʅ'���"�tK��vc��Dɻz���3�������ء����\���n~��}�mH<r�wu��0;(oq+�coN�yژ+�4c��6*�ט�ڛ=��u!n�rd�N$S�vٜ�"��X#��>f�6j�ı���>���Ŭ�.�*�j]�3t-�6�z�bpO�H��xIlT�8������}*��� {����S�rD����˄���Zed�o�(�|#�4�n�ٔ��G����5$�n��k������J��A�)�q؉�)���Z�����Ԗ� ��>���5(q�9r�e���E���5u�����H����0��7-�RCr�`� j	�mP�<B1j�
v�����/O����A��&�n��G���,��;?��u�_}��&2�����-Y�|��rYED��Gu�&�3;��DE's%���g��J�b٩zȏ��A{����{f�k.��D�}��eU��N�y�}�=AFG)O��̝�|<B�Â6��O���,_���+U��yPV��9a^��'�O61u> ��N��~�c%�v�hJ��; ė����Q�VO~��	��'�e��#l 3�a�ytCK�DOu�,��s���� ����^vV���y��fa�Ի�xmwi�(��mSw���(B[��(���g%�y��{��`���^&
^%�yb�q|k����.T���<)����0~0O��{�%&���{� �N� �C��آ�{�d\[�-B��F�2���䈧�F�ɮ��T���1M���q`��v���d�	Fj�$�0��`���3fL+��F|�C�;���O�<܎,�B��8��Y�-Ⲝ>�.�eCB4A\��K�җ�/Xt�%�e�fD�m� ��sr
�]H����9��HV2�ZJH��e�9�ƌ��Y���h�U��\��"ux���oOZ4!o2r~�5|���1nǛ�R'� ,Ѩ0^����X�Ȁ�m��.C[�Ah�9l<�KXK��%�0.�Q��'93�^OP��HQ��	
{��4G���7;e+�71�&�]�w��1Sʾ�_�n��X�1�&����DVC5�)���g����F_�H<����j�ls�г��/VC���&��.Y��l�BVT&�YO��vFR�q�v�<p���a&m�p�않�Mr���OM���L���/˝�'iF	Xg�F`�c��G�@���	y��!y��Pu���C��Xo{��Ea�4.�p�9�J	�6a�����#�	�FM8 �㾋��L��ۻ �J�o\o���R��r/
�ؤ�0HD��ʎݟ:��p�tpPMxt�\h�][2�֣�P׎�O��6*�FDox	���gg5�f��ff`@*	b�o5{��&Mݬa��e�'��4�M����z ��C�r3��ڡ>��}��@]���[Bč�ۂd2!����q�����b�@	.���ѽ�Y�8���S��g0�!h��զ~�8d��<)Y5�5�w�2/uH8x亮W���v�>_z������x��(�1H��y�<���(�����v"K��6]�D�����]��(pi��� �E<7aGVB��,|�g����.Mӳ�hv�#�NgP��'?� ���)Fd����L�n�	l�G�)����ά\nU��Q��5��^YdE�|I֙�n##�K����C��%��H�����#�^T���,��n�r79k��3�<�l�g�E��� �=�+a�J�*Ȃњ��1TEE(j�I���bfGI�s��!�5/��>&��8�o9�b��%�0#��C%�ukSr�X�X�(��s�64���6!��Q�^�`	!;�>b���T|=���	�Gk��^�e%]i}���W|���ħo�5��7魛̝ߥ�#��1[�=l1��
�����a�����Z��4�H���Y���$��>�Ky	>]��,+� i�_�#���"2JO�7&�X�ݸ�{Α�zsA�I�h�s���~к���Y�~�'��ʋŬ����!eX�*��vIZF/�N����w��J_��yn�/=;"V�Ĥg�#֣�=���0�7<fXՙlX^�k�b�=�z�yC%���Xlt��$ċ���> �@��Av�q��cű�n�!v���&x�@k��8��y`���jB���A�@LrB���P���R�3ZB�tϰ���bͨ��R�X��+�,yB���h�A�Z�.�x�m=�f�ޑ��4ӕaf��P7l.!���7�_�Ͻ�_te�8�����H6~#�����fR��<�\��% ?��y����2B|Cm��f"�{����J�����F���|E6��x#��f_�^^Z�!#��Zw4�`��Ύ�vz_�!�R:g�b��=¾Ȅw���Y�w-ӽ���[���L�)���Y@���BF�V.���	����8F� p�g9=�[2s�Q�Z�
�\��wV�S��E����W$4{)I�o��2�g�	;ɒ�F�|���ယ��/�7���pn��1�&}�D�:�ӵr6z��'JB�@�y"�G)�;�}iW��'���sX�p�.sE�l�P�I{Rx�RB����Cլ
���J�cg�u:I;�Է��oľ�z�\QJ�N�*&:����������Z4�;�n̟���k��a�m~͌]� �t��r⢻%���[������i�|o�#�,)�<530�ZӴ���I::ƔI���Y�84hu�ʇ�]��O�1�H#�#�9w$�����
 �y'
x�`jZ9 ��,U���w!*���lZZ3S���	�ŭ���#���1��JJWBg	�P��WzZ���7)6J��}�~{Ɩ�0����f��b[�W�	5�:���3�V�nOׅ�Z�/1��t�bl�~Y*d殱Ց:�	���xnD��~�!W2 �mPв�����!.�l։��yM%�CNp���5���ea\�������Қ����!��R0��Y	��0	��)�G((ta�4C�c20%H4�+��k�+Zn��>�3Lۮ#�W$O�X��v�f����[��l�'L��� �&n�+kZ_�j�ļ�=�7(U`ա��PLJ��;:�^|�1I�r� ������j�H���K^M���#��Wx`�i�}����h�N{�>@��iĦ��y�e��������1�G���f����F>c��o�SX���!�<Μ�ɵS<I�O�ݿn��g���0 �-⤘A%)*�W����5{h�AZ�0$q���*L!�����>e��H
/my0���t��5�T���?��էT��bq$�^�%�hޟ�Y���$� ��a��ړU���+���%�Opm�����J<2�u��@SGG��3ϵ�����[���v�Nނ>\�z6z�����3d��]�5�Pؚ"����MWR��$C���<9O�8��ۆsJ-�J�����o87�gC<)��౶�Bo��ҥ�ݹf����ʯ��"	�o̦.��Y��BH̴,0�h䙖]�ջ]7����;�o��!�ǋ���F��=n��v�q�S(@����e���2�~, ס�t9g_�i�g�x�p:�)�Vkf���M��:��)_~z���ͳŮ�솠8W�FO?�etA��]Ȫ�Q��.L�9���BZ��Z�	���N�?�g�$d��������^RIth��.���t�NX _g��]���,C��v�-���>�K�Wq>�u���Gv�~��C�я伝1�*4P����<����Ju�~��	����� D�XM�ͨ�~]E� �����KJgOVPQٴ�_�kt-�*�׎iQ��E��iMP�^�",zb���[v�Yf)AcE.n��2�ڙ8'����&�b˃@���K˃���1��<��W_Q�㋔09�&#Dh��
����"�����6����$�=��hc�FR~5��|eԉ��J��Ŵ�:�~	�aA�̂��w�j{\µr�f�^�5�'ǎ�����
�Y����w�C@���i�>�{���c�s��=OѰZ8./o]�`\��lo�9Pc�K���.��C�y�O�M��}�t$<6���ρ�q�{cf2)W�����9*�����S�� �J��	F�z� m��5�ӳL�9��6�~��G�3Ө>��k�L%,�O/	Tn�5�bka�����o%zS1�`��q��x]�
n:�G��fIW����c�����j��*n��X�._��"Լ�Z���MI-`U>5����Jbh�A��i�Z�#F���e3p��8-�f�`�\|̩&�K��f�J(o.�$��|wϚvu�CDҽ\��5i���Io!ĺ�83`qT�C?�,��aO�v����9n��^~S������qH;Ul�X�S��4���pZx��4vga�E4�G�
7�dh'%��/ވ��(ٓ�/�AUL��E�\��O)�������"J�D�8�T�ۚè������pp�;Y'F*d�'dv<��v''�p=��#�R�����#�������~DLz�"��6%���6�U)���8۪�2	����	��j(p�$w����9lz�2���+�����B�"7�a6�R���(�D؊d�X$7˨�:��}����a,/���H� �ݛ����l!���s��z�ӧ�z������Eh�`Nq���R���t��_*xhjt:��<�{����<��5^/���jY#~u,~�g�؅ZG�l:���UIT\�H3�����F���������ٍ�q_��B�Z �L��nYA��}0Hhy�mwS����~����ג�ӍJzg�%d=�Q��)��
N�AB*1��o�r�Jq�~f�^�=�/w,�c�T�N]c�D�m�ק�R�|�M���J�1�b]A��\/#���Jv�V�1���;���D��͜-!n�>)h[��lE�'�>5�r��x�)�FHr���2Yh�:��~S�X,^paQ�;`���U����"���k���={4�x%��g7JJ�*��u �˶��? ���7vIvַ	ҧֈ] �a�2������ˊ .�{�1m��]f������c�)�[�4'C���T"r�$�+lr� ��Q��`�0r�A?��
%d�O��I�׃����>W���������a؋��Z�T�o"�����]��:�6�0��H^R/m�:���&Yo=?��"̤b��Fw��."l�:����sIF(dTk5���I���c�����Do;�أy�!4�Su�g���1�:��n�^��9�D�!,1 �YF�.�lz0��1i���/h�*9ק'n���V��M�W���:����2����D+$t+�+z�x��]��D���͋��5�q���0��85k�>{,UP�ܑ �3�s���%~�Yͬ�@��qDURо��M�p�`7n�7�{V)�yϝ Hzt߿��%@�R��"��sO��gj�M�$䠎����1�2}t�W�u s�&��#Md���
=�.�kT��f��v�٭��*C
�]�}�B�0l���'jjB���QQ>�*Q����n��<u>s]�����(ň2؞K=�Y��E����H(�^�1x��(~q ���l�-y��fst�a�[,d�Ap�LiB������cA�sr{X��v��8��?����<�"�)���jiW�B�*�5�
mq�������ͺ�<�u�d�t��<�������~�b&!��d�2d���_�q�=��wi�قz�r�Vl�m����+ݜɦ!Ϫx5>q6c����*�D�o|�����^���,�緾u[֚H�CAR�[2L�^[D�"
y��M���B���wo��q��lv� ����	���_�i�o�v��*
D�N*���n�
�҂����$�l]e���A�1 �V�O�ݸ;�6�Ě!��F��7�(���u�Τ�����H���1E}����y!eD"�h9W��+���k%�-�FR�ϧj��T��{Mw3v�1Byف.yMMU+�����5�f@&�P(w5�%�@��7//��xTyw~ۧ���&q6吊����Y�>��y������Bg�!/[,�nh����ˈ�wT�������u��C�Ml�l�����-a �����d�N�ی:�kq���t��np3�n�t�~� PJOwo��ZsN��ˠ�V��N:�Dio5�U���\�����()����'�_���M	 5j(_%����}�'�*s\�Bb��؂�y=���4q]���9 ���sE��>�Rv"m�L��fƿ�K��~��Cf��:�@6�6��ϐ�=�)�K���M�쎆3L�Z��gb�*ͿdI:_�W/rT�.u[��~�H��źԫߣ=�l�� ������.�Q�_㻊��4h�!���>���h��̖�V��S�3v�<�?ϟ\�+��)��ZA���	� �x�����"nF�t�Wj��qᵩ����%(�?�OF�kC��^��{/��{�'iA��E��!R���(������ؙ�T��k�=�AqQ;�ź�[|pI������-c;}���7�|���5�HLI�q���D4?Q��ܱ���
%+T������~+��r0]�`�J���5��&�"��E�q�����ER�P�Sf'�x(�F�4���#����t�|x:�qc&�!3�6��٦P��D�2�����2J�|-�+�����'��I���|M���{f{	x�]��r7	ǆB�A�Rx	@��jlz&~04�-���$��N d�ڲw%���
OI�y�6�v�!I�O�����l�l0o%�#ΕT��ptl�4�l�Fu\��p`\p�T\{s�dUx������βā*�k�u8j?C�#C���Q<P����Z)\"Y��������w�B߹;i�1[(��Q��Q��m UJ�v�ՙ�H��	Xb����Y���4˩"�Z3�!-�J�KǧҎz�
 ��.�q�4J
����ٿ�3�7i,�8��}� ��EY(��xT��{�E^*�)��)���U��d ��Q��*h��3Rߝ]��0}o3�1�B[�S 	V�-Ԧ4)�^�����+hʾ=�"�aM��C���5 9E|h��feck�s?$��8I:o@nP�As&��ĩ�0�&t��<���tҟ�1�'&
�"aW]�̡<Q ��>JM�/�<��9a&_��V����Qu���FJ}�.O���쨳^��𓺪��@��{�i|�Y�z-�!*�������������{<!����H�b�#J�ߦ>*�Ng�\���[��ڿ��4���}��Qd=RcB_,�]�ksV]:������]�*���P��8��Yz��<y=��3�!�����1�����.�˷��s��)������3;K��;f����1��v.s)��k��j��3$�9^��0�+�W���/yI&���J���[D�%?�)���$:p�V�G��g�} =�*|`QU��`�S��lr�B^��R�!���,�I;~`���U��9ږh������@V�L�#J&ix���EyS�"��r� t�Z�T83Y:u������l~�J���1J��h,��#�"��������>a}d�/*K�k�i�`%�'��&E�8?�ڶt_�<c!����'q�r��q��޽�ŋ���P�LL��� 
�Im���UMQ�ө�8�+����ɩ�� z��f������ݱ\V��/y�Ptm/�y��d�$&6=��ͺ�]�L��'z�(����XlM���\#���^+�hc��E�)�n�g^�O.Y+�<�w.��36+tx�ӣ��˜'X��r���]�2H����5aK�ֳS�_���<B�d~�������UQ�g�#�{]�� f��Y�~7�Ḯ���`�X�#oA�u��,���t�r=�i�.	ʬ��" �Ou��`%�
u
\�q�n��se[[���i�2;�1yBJ���IE�0[C��"�6�A��&�E.�׶��$_줻�P5D�y�|/ܱ�L��p/ۉ�g��Gj#1�e�8��m���O�7���܊#H/���bw���e�+$�D
$�I|VؘP���Z�u�_�EU����b�	�+�D�6�ɘVНTݩҔ�Zwe�D0�vm�5?�!��b� !m/�nuJ��Wy�_��xրC{���2�L�Z�j�S�Ub�,h�����%m����D�42V %?$�D����={��5sه�9`��́?�=��-_�-���Khڑ����C��c�*Y��Ka��0�N��=fr����[��h�� M?�bw�{��9��f/丼7Uӵ�#`G�oz�T]��C�HC*Ȍ��?�"M;`�_�Yk.&�����5[�l{��eנ��]�/���
�}Zi7���v���0�!��;�>��=����(�Bw	��cq~�lVRD],:�k���b��Q���mJ���	Y���)��xq%J��N�),G#g?ؓ��h,wBO���^�w)�����%���g�X�,��s}������㬘���& Wdp�s�۶�����L?�Y���0���<�T>��o(T��&������i{_K�j$�D�*pO.?fP�O`��؛�j9p���,Z�fBʜ���1Fß`X��)�L4(�s\�1s3?�f>�����(|��i�"k������.z�ٰ����	�^��X# ��̑J/PAF&Z����dr��(�v�F^��T����K��V2�
v�YKH��#t����	%�N��v�sA6�3'
K���.K�����nZ*!kLB������]J�!�}=�m���e�	w�p����Q��s1���
R^���k/Eʜ,E�o+vDX�ܦ�0��i��ؔZ�*���m��̂�q}��dSڳ`}��\����d��{�g�����_��k�xJ0�m��g��
����:G� ϯZ�"�b�۱���+�#���4��B�����P�L�L��l-InG>�/�u<L��`������wo����!܍�B�'�*n�5�W��}�k�7�z<A��*�_���b�w�G���#О�rK|��_I�Z'��%<���=�m.U��~q�h���^���p�u�"�; ���#)�����4��x�y�m4(!���#7���U��N�_!��">5���}�C΋D�,���Ҙqս�^�΃� �&m:��L�D�uӬ��_�&(�t�\5Vވl.J����N#&nZpMz	��g����cv�s�q����o*��`-#�{��������\�SG�G}*�l����n��5���&�6�M9W՝ڤ�C4h�<�)ҡ�i���6Rx��晃�<��%8�uY���YH�)��������0��r5)*F�����v��렬L7C¯�M��"��5m�����i��KKA�q����wLk��[6=�Zfiʦ�y��0ub
%�)�6Δ��7�a�<4ަQ��.�Ѧ��c�����v�d\�űՋ0WFb�T��IB�슚��р�iʩ���c�C�F�Np�6�-]�t|�á�s�ϔR3�[��d��}x�8ĺv��J���8^�����ZSB*r>iz�6�狂��s=l�s�bo��&r�p)b�Y��>�nM!1�� dE2=}k�N,6�8Ǆt�<�V�_9A��y6�$��f*0r	�	�8���.�H�i3�9��r� �Np�4鞘7u����H����n��n��c
N'�r�v7y�G	�ߧ�l;7�(&E(�\����6���y�c�l�#�ͧ���k�xS�2)��_�x�d����W���LK��Xᅆ����ĩ�0�,2K/r�̐�f�gۻ�J }w �T|D!�iH�%��cL�����]�]l����-L@�����V'`},D]�x��lx���w�&��GBξ�K�
Vgl��#��H���$?�ÿ>�n�7�W�D����I��	� �x"�Iw��8�X=/�4��#��M��:X��ʌ�q�����K��Ny�~�ܐ��R{�y���RO��q����?�_�d�i���f��Q���3��S?�u�6O��d���/T��ó<��vE��.��{ɴ�h�n��>w(�V@(��:5�>J�Ę��)�7U�jA�XtV��I+d�Y<͈^���e��Q�h$v+��t�V5lA0t��C�x��9aY���?�2��PL�QO����٘J����iL�� ��b�8��)��M�Knh1�$5L���mX1���i3��$u��]O��_ϕ�G��DK��Vr�X�u� .(g@���'R��k�e�{/�d�3 &ز��*��������Yw�n>cPa�G�2�r_P*JI�V�2�?�:m�OzcN���t���>G�2�2,�'�$�:��Ĕ�
�ڂHJ������W��v�֬��Af�4��V���Y�����������0�z�"��x�x���Ͳ�z�qF���g�YC��%��|sVI���|~zIu��x�j�dT�:̹>l��}B�c�a���oo[4�A���2�G��a��{S=���_ltLzY-�_LC�&7Ô7�U�::���#����9:���bV|�C׼�k5O�ǐ�e����qc�����@�R���l5��*�B�sK}נwMy^X�ej�y�{,r3�R������t�e�<`-E�V�t��
�|���72��aCo�� �+��$�9;���Z��[���@d��z���|L6�R�&A�l��u˘�� i1�\)�qg��tk�[!$D���N�.(��3����Є���u��6����K2�i���E�fEcV�Ӽ��~�9����R"i�[O#�%��챂ͷC�g.���]'3��a��`��Ҕ`�$�@�[;M�����>��]�����^���b�?�U�!�PFs/xਅ�����B�X�G��\�H�ʅ��H���������륯�@�b�B�kzp</��ZhH{�~�����Y��0�7˷�*�;��Ň�� �r}15>C����&�B�k������0;LT�� �×k��l�o`Mgx�l���K�u��Bl���j7���_��:�:�X��U���O�dȦ��~Y�a<U�.'��=�	E�Ũo��� �zS��3���lNb�JlL�W)���r�)A!H��~U$�9�Cx:߈��	~�v P�65֓s�0 �q�*�P�$hB�X���JԚ���38ub��zk�!��9ơ^�X,
���q�JP�@����R��3�D5�a2#0@4&�N
��c���֊
���D���������8� �A�M���`����p���	�[���̂l��C�H {Ҍ@&ѱ�{F@i��΃�\+Gѡ��n������e�mS���M�O4{�����R�ͽ�6��'9#�@���i99��(�o>9���'�gˆq�����{�Zx��"v�e�N�PP#EƟ�*0�57.a
�[b��HՖ"��u�P�+l7/.�)=��)���B��@���TL]/�Y@AFv?�.�Im�u�*�W)�2;�#�ymUKjY�L���a:�J�tQ-����jj
�TG0mz�KdD~f�U�!����tVA��y�y��M��7���`��0J��a7��
�l�F�z˓����y���id�Ƴ��G�;\<T3W��\Hl��Z��RvZ� ��Z�ݚK~��1�!l�j�H��iP���Q����XR��ǿ�B7T�/y\�K��>�����t;�������a��,[x�t����:z!�c��!Lϟ�g�
��R�UkI�$�}[�g�%MW{�2�2l��-���2?��.�fl���3|�e�u������`�LRc,�� ��'d�Z$�u:ޯL�	oÊ��Q�V�*��N!O��9��J	i��ɭə_E�B��9�r<}�#��0����̍�!�K�ܩ�^k(b&KV�K��>b�@�ׅ�3~�	5H3̀���W_��c�D5�g[<X�/{���7��� ��ɵÿ	�9�\چ�?2g{я�Ʌ�o�Jsys����#�%D��W3��� ���XÁ6-D�s!2�+`��k:�������.����莄��
+���;/�����ك�?��D
ͱ������BA��̧�����V�T�&��Q����*[�䇧�#p��n��B�֐0P�<�N���d���@�������}3�46{\��D�L���^���GY��VYh��}��*�^�pQ�n�Ԝ�c]�1�-%��?j��&��W����M�Zg��"��`)�8�m݅LP/���8M�Q����*�������?�^���#�����5��'����V��tw
�>�f�0k��i��|�����J�6��-2����ә���ۃ4f��P1�-qב	9^cA�j����{l9��ɉ�c�i�eQ߹��f���C��O���A�U�W��528j1�Wm��}?����mI�x̾H��EZw���y긖i܍��m;�n6���D����;C��y9����NN�՛rP'r�G����qcI�;M������ZN�tA�rM���@uF���W<e&��R��vV��{�P,�ھD���Z�Q�t��\CQb>�N����\���K�6A&ta��j9�t*������m�`��/'��a�u��ձ9��_夺�e6�?5X�9e�!d��h	��Y㚁U� ���wN�_���5	�'l��H0n�r�U⎽���s��GA�D�sFF</�e���	!c�,z��ҥ�����4�.��*�8�����+h����Yo��ؐ�|pA�CI1��i��_RmX&R�D�,��p!��@[U��=jM�3G�V�h+U�@�a��	K���
 ��|��"��4����e�u-�8P\C���\|Svh,ef�ݡÉv���	?�Jy(S�t�v�˅����Y_^��BEv�{����|�O�uC�2����p��1/B�SS���f&�e{�-�Y'��!�>����.�&!Б���;�1�.0�f�����H�ힻw�n+��=X.�&���XL:$���B�/PrD�^)q>�%e�m�k�N6n���A�7c\�u-~�څ;/�������tk[{/��E�,��G��D����L�t1(�v�̈��M�y�[�+qSѼ$>i�2��/�}G9���+�]#��z�ɯ��]'"��OьEy�}�2n ��s>�.5�U�*�+x���[��Ɯ��$%M6GG���ǱoO��[�<D����C4�ǻ`�oV�J�%�� }P��˨枧��e�I�b����t�i��1�n�*~�]�!�f�D����Ԉs�o���#XHަ.n�la�~AZ�=|��xS�<�
�kV��y����y�ɣ��Un�ב��Ɛ�!�6h�c�S��~�jB����?��r�Őm,�A)����!f�wv �0c��+��8��!t@f�z�4�v���MzܔK�Hɷ/,l�Re:I�x��th��څ�jE��t�.�Q"��OGJ�i�~����g �Ҋ.VktI�6F��dܬ����M����������_e�(�E+ES�H��B k�� ��B7�L�N���4�WQ:͹��i�r޵��
�=���x���uW��4!��gw7��2� ��^�Cyæ=��c��rq� ��LA�&d$�3�zt#�u��|B��m���[��8�dl[�N��i`�n	��S&r���R�ћ��8�1zl�{l<
ӎ�c�h�B����S�̆Pڡ�1�g�@�8Գ঒��^�KB�Y1Ӫy��2�`��������H^���h��NE�T� �P����T��O�˂7�/��>G�/$]�[H?��\�R2 �F�J��?���>��є��,R�����PL:B�
vS��E�}��5f��"-py��?N#7L���Q��N�F68_f�	 ��.���|��}��x鯠��Q>�_�D��<�
<��Ƶ�����ר׫������\��UCf�b�w����~R�GG8ل�x�� ��B+^����[7n
H��UH��?]�X&-d�������!�73Ʈ�����(|���jǌ�Z�a;?P�TДCE����Uy�O6�	� ��M�[��-!�)���,��QI�����8gr*�-�ݗ��D��8��ِT*�GS�3d�b�'�ե������g��9-r��$�
.�;��-s/�����`�L:��*����D���-2��b�z�sch���&��D�K�f�y&�Meќ���?$kЀ0=�����z(P3YȊ���Ǆ�-p�r�AGn6��z����i�) v��Q��C�/��S�k�f_��z�.�`�l��(}��������M�~���W��iü�|��U���Ť(�%j/LY�Q-z:�:�@X���pO�cj�hOwI�qsԷ��I�p�S��기��;�Q��{=ԇ�������(�9Q�I$b�x�䋱�c.���"����)s�b%t�}�q�ۇ+��Lh�5Y_՘�W� �����!e����
.r�_e���N�k������)`�<�5+���r2v��C"�S�f���X)|;v�+���ʳ�aʿ
��8D���/P��B�v��a�D�:b��0a�\���_sM�]4�Y�Xy��ξ�|��_E� $��D�AA� ;�#��"�����Rl���mV���}ќ�(��I%j~�=���~��fE�<����Dgt�ѹ�u�䶐���q�D|B�����3���s5�����/�=��B��?\e8K�e��/��O7tD�B��k�%�y��@ڴ&m���JS�q0�}�`S�C%t�ɉ�
�����Iӌ��5�$������T��m��@b
��E���[����
͚G�g?�L >/e�\{Jo��W���G�7M9��Q�q0��T@�"�{�Xy���
r.:��#9�������[�p'A׽Ķ��Bơ���$<]��+��r�B!���nd�y٩���.�i:��A%恀K��jL���|| �������9׶��G��Q�*8�oy~��8��S^��B�gT��$c&��ֱ�?��@X%�����H�g6����Ł\����������,V(&�0�4
|]eg�>�m�8�RenЫ�[՗����q:�W�T����^
��Y�/�ϟ���~�Ja�j���s
]�b�:�;2T;S/5���r׷�Spb��,�n2f��:-I~�h{��ξ��əG��0��غ�Ad2�f.���yW]Qdq����B�1�]N�����?x��o��j* ޚ$�Ez�?|L��c��z$�OFk�~��7�zop�4��ft��RC=���j�.�)n�~ϢLx��9"ry���L���b��R�}5�k�[94����sѹ��&���0�U�މ2S�.��Sqi�W����e	v�h�*��{�݄�&�UJ+�w7v\e ���/ZvY���mz�����C̙i�ۄ�}]�b	}	�j��w>��&�a�O�QF��d�#q=
�i(U��1`�'ǔ�On�`��^8� ��.�������f��[���,�aj��XA7nw5�5j�L�Y�ǖ#a��8ddh�ӻH_U�aN����g��w'=?F<B덎��M����Y�ބ��]�7)�U����P�dA��Mɔ���=T�32}B�$�i�$����\P�@�<;����F#�[�Cۆ��3�7�>B�(	�x�΃�i{S����NG�x��x��%<��C���|��u� �� �:g;� @:�?�n��O[g��8��7�չl���H������Q�`'��wt��N$�2�9�d<��p/��N��P�S~��f�hZ��/���>4��&��#[�\�e�Mi�"�,�*��Xs��ms�;����hvI���GC���ѣB
� �CpH�<��򊽙A�6,�g��I�
l�Q	:��('B[μZ<���u��AҖ|�oI��-=T��w�-= ���ֹ�.����(�g9�gP���F1]7�
��.��n���7���4�������j�G�Bdt������F�[�)%t�>!��Q�O�3�.H��W�NQ�H��[.;�Ё�no��b|{PR>����ճ�9�m��Be�Akﬂ��S�������`}_/>t�È�d#�	�b�ŀS�(^ʹ���}Bn?g&^��AQ��;�m�׿�{O�ku?&�@��q@�@�}��$��Dkk�x��P(;�?� BK�H������D�}0\���ӭ�9P��.��۵lɂ�0�cx�/��MI=H2�$B��<�
�8c�U�G���C��C��6��a�ؒ-�o˱��r:�A:9#�2Ա�MgT�D��+�v!8*�'8�J. vF4�M��g=���
R����Uݝ��J�Ci�x3�2ZM5�!3�9y�J�~�O�LB���k
9��l`�'���L��E�<g���tnD�G��Ⱦ5jŰr����ms�0�i�t��t��>�Z*�F�9��?��~�-KS���,����Z,�`��cPL�oH�~}��;A�<��g�Hnn�Uǉ\8AeǱ/r�qh+�e��#}qZ��4�W�"?Љ�Z���mؗ��G�s�N'�O8fXО�n
��Uw�X"�҈�A�R�cl�*�����SߐɓxAi*�N(~��G7�Ģ��<�s����^E�x��� ���Fa��wvVi"s������u9�/��?9�~]�.FMFk p8]�5sf`�]"�M㴌h�^���7ڻ�.�th�T[1$�S��TOa6�G����~�Bxw���C?
j�K�&�nN�c�BL��a��a
�RH�P�W6��؈YX��:�ռ>*"�M�,՞6+�Yrպ�#��_��e���zݩ���0���z��GLC�:b�P+4<@KqaN��ÔHٜ>!��<����0F��}��Su�z��nP復E�K�#|���i�E�<�`g2�6&A�pר���z�B�d�U�X����4���ׁ���Ye&k8�ϟ�v��]����!2�.C�3��{��W2��W��H2�z#��Z� �q�zY�I�^^p�Z�Z`�&T�S��p�ܫ��_Â�'�֩��:��{���?���"�1=W��)�J���G�2��\d9aɿ[J����.���<YjS���;DЂ�50�"f���_KZ�`�2�T��vAi�!���N�fG���z�n̅x
�M�#&P����������\�D�n8�H��hF���*�r�ܕ{s��fg��� `�!ٰmg�>�Ϗf+9g�a"�Ǿ�UuZ�w��r��	�N5@��Z����3��MJJS���0���[W9㌴� �_[���|������_di+.	1$��l�;j�gi���3C�p�3�V�k�>�O�J&�WATqCŌ�7���U=]c^0S�{�,���A���} ɪ<k��� ���Q̐�?�s�I���OҟL^ҵ���,Ii��*cHՒ�A��Bf�!��a�(�(p�h��W��L"6�3���y#S�{�cm��Bp��P,�d��������߉s������E���ڠW�C��&�	#�;Y+����vA��T�u�[b�&�!k5��M�Ä9ESF��On[&�yPp�/�"��$�O�.���7��nw��R"o�X�%��	F�R��flX�o���>;焭qZUe�aHӊ��f�h�	��:EW�c�	&���#�<)��tʎT���+�.!���i|P�D��"P�}AO��p�G�%��t�	P�� ֖|������̳"�栄l����o�x_Q��)WR���ٜ�������"���sJ��_���2J���U
��4�'���ؽ`�Dnz
}��ZQ'H:Xp�]�C��b��a]��R|��>w�t|g�e?�M����>^1�Qq �;��ؚ���j���wra_�K�[{#�4b�O�j��Hl�J�+7�����y��F�]��AI����ڇW�K2��8�c�t�:�����[=8�wlb��!���j����l:��zdW�#�W�s������-Oj7����@ZSո�H��'lݱj70���kX�����������]m*5^�;���&�C3*,�"KO�}�����q��� ZUFӠAYm� U-��I�2Mt�ÔW@����A���<-Ua���5{h�{��"����e�2h��#T��+F��4޶�#��@T}Q�b�t-��K]n�4�Ր�3n-R�7+�L���F%�y0���CDo�=_ѵd
W|c,�bi��/>C 1`N�"�M.���Yr(���U�x�s��bt8��*bA<�%�~�,GkC���2�VFe�MR�������p� �)E�h){x���w�zT�����v2�����D
��c�dYS|Xڻ���w]Y�q���ҥ��j��'���e�G�*�������P��?��HCf����+��M�n&��D`h�p�/J\�'��g��6@�������4�nXaJ�P��H���O{���U!.;���F\2��=���2��^8
�'���|���ar �h\�%ˠ�����vqcUcXZd�rHL���>�>��y`����x�����"���M�ZW.�b�E�,<W@�-D���C��g�Զ���
��xV�6 c����ѳ�f�:��9U�Z@���B��Is���NJ��>^60!C4��u3�1�n���Kr�/�d	��[9�Q/�{X��U/{Wh_�BD�R6�b�~����}�{8�*�p�u�C`K���:�k��Ĺ���Yw�l��h]�-��祊���Ě�F�k�j�+�����s�7X���[M �)<��/҆je^��{Cye1ܑ-������S=�h�:�y�� �9A<�����F�[�S#X/ml4?��(}? ��%R~2R݅f?�`���GjJ���pz��p�O�uj�+��ӣA������G�A!�o�X��5X�ӱ��?��>���r58� �(u�%M�B��.S�%���_�"���y�ޞps굙�҆����s�G�\�4(�U�&N2S�V�)�ϪrNF��pH2S��v���/G�^��w�w�\H�T2���q��)��O�N)4��O�JGN6��+
�;|��J>�{�g�RK<�e]�6�s#=��Bg�E��*�@�YnS�`ZT�{�7*w_gq��$���\s�".L��h��z�FE�~��HK���"�r��_�� %{� ���;���R/b5{R�s�Ҏ��N��Ve}�a��W��N�Ew��4��v]H��[������/�i"F�;츨���Y�=�k*�X��i�<�G6�Ԛ��
����)/JZ�<�h��s[w��}��+A�q�Uk����/�B��M�=>H{U#��Wp.�"��m^hJ��9��$��9hc�^xDR&���1�UcfҰ4����jH"	�
��lϣZ�n'DKΎ�n���Ti�����&<�
��c-.��)	R��y�q����z2��lzxyo��e�y�F6r?�%����	韖���0.�+�����i�O9)nq���g���"��g��TOG`�F�+*�oA?�MO�爁+��a��/��M<�S��Wx73����W ����p�>�3�֜�ݭ�E�˞�#�D-k�:t&s(�{%�GZe�H</���5�I�$!f���r�%NE#"����0������Q�G$"����8!�����+�O�W�%���wZ���i�V�I��Am�=�b�J��9���a�qT*������&A�,vs������/��<�HX�5�1�� ���pQ�7^������!��\�](" ���!+Љ ��U�X��ۤ����\éOz�|DzA@Q����>��2��38":�봯����z1����b�h+�����̊[���7%��*y����lxs�PpH�� ����+��ٺ:�r�c�-�+����њ�Ze;��4GP�!h��41�b�7g)����A� Bc��	VKA����Ӝ�|�@��nH���JS9y��M������ȿ����������ګ����A��qx\��BOlE@�ƶ��O��ɂ�cF]%�0�j.�f�[�R�?c�˟1����t�@^ `q�*s� ڲ�8��O���p"�3�od�����s&C% ��"O�P4�)s,q��~!t�ѪL!+�L��9b��0h�#L��e���~�9*��u� ����h��e�v��s$*�R|app�ܙ���������B�^�Zmx��6D9_�%&A�lX��,@q�X� w8Y��ǐ+�'�/�J>�[��"4�t�b)�=-�Hv�ɭH�=n��L���ňh͠�R�*�
��bK'=�)M�+u����O���D49Hb,[��Ϟ�ς=( �p�J�=,o�y?~�.��i�����euN�� ��/�� ��7��_��L���EG��i�m=e���w%��UO�	��G5UGj��g�oZE˘}dF�F��~;\��V�DęvPT�9����n�~�ƢC��SG����ܨ��Ƶ��n��o\�H>i�a�&���|T���b
Ր���?������e���iū�$��7��j o^^%�z��y�FQ ᢡq䒵��1�JD�y����� ��uĹ;SWD3�v[hd�O�GZK��J9Ĝ�Sk�4n�{��s(�l�9#R�B<5݈���"�~���q��:QV��+�L�z\Ժ@\FHt�w�l_��p?W C$`p�M*�~6�y )�#�P��:@�(:�t`�����$Hj6����=���t��[�F����������@����B;4XeH�n�Z�Q�vc�O઀�p�XY��F5��[A1?JeN��2�~ۯm*WB��/ު��e��#"m�7��!��_�X���Zb�&z�aCb���mӑ`��m�����;��	�>�{�j��y/v��1�c� }�OJ��r:ҒץG��q�������Rl�0�a�e���V$�n�$=/$�kE'*�>���z
A�<���_����$jW������{V4!d�
^��C"�[�J��L ���������6K����6��	�8߶��`�w�m\hHG�Nټ^8kg�-���9 ��S�"ƺb�\�ڇ��K%o�Ӟ�њW�]�/C����~��S8�9�5ӭE:T�L�U�EDGF�`��7���o��҆(�kL���(%z���f��k���M���;�Z�x�@
XΞ�'ga6�h�N�|d����ԝqe�C8JOE����~��⦉��O�H�G;���j6�t�n�s3R�o��1�������H�4�����-H�#
� E״\��7ι�DAX�q|7e�9�ؼ�$����khmK���BSZ�6M��'��l.�i��h��G�� ����3���$�:�`_B����\���80�Ly�B.����OV ���=�3A��Т�n$ۑ���?;t@ʺ-_I)�ޮ�SC��y'�6�g)�#*&B����c�M�ܒ�}t���I�"�J���a���[[�Ldrm`݄����5���a�/�ť���BE.�Qa(�Ԙ��Fx%��`G�*K������k���c�n�N�2G�|m �$�h�` �X�oL�3�dU����Vڨ���-����'@_K`]��=s7 J��!8v��z��^a
�@�X)_˹��G����8O��Sdj��1��k�0���G%���D���u��߂K�4�H~��*�ň���UYs�_#��X֓�	@¢�n��`#��E�e/�X����xɳQ��m��$ͅ�UPk�u(�*sT�fp��R�x�m�'Ir�E�u�񉡚�pj����S;c$��¶I�I9���?Η���~!F�ު���d�b�^GU�� ��[�ӛ�՝�f�T�������sI�;w�:A������O�T�h�o�� ��Z��a$���Jn����7�s�����O(����e����&Ssȗ:�*�ײ�3B���S��k�hARV�c��]z�p&ll�t���-�@�e�T���a�r��Dq��}W��s'ƴ�}�W������s��G�l��X�-d��2���������읡���q�ae�8n#�Q/R{J��e���/�i�		�9P~4�L~�Ri�4��	#� �\ ���B���q���7�1u��v�L�򛪜?YS�,��1?� ����>�9{���H��J�ީm��rj�������=���)�����)iZ���U �h�Gy�w��$R��9�����+�H9VI�)����'���1vd��P��k��4�3����
?UH�?t����XC�@�r�4/�J_�EBq�)՞��j%��ord�ɀ���2��xQ: 1"'���?�+�C�F�0��֗��GY�d�I�80�Wo�Bb �t��=_�ˬ�|�
���g$J](�X�)@k!qZ��zM�읡��Q��@��sQ��O��OPS�����k_"�rb_�XaI���
 :��FD���`Z�*�bS��Q1Q- �0q����]F�=]�ka��������&��tpJ<��$�����"��zU�D�DdA��k�Ä�ݐ�e},˧GX��=���-s�W�9B�+|���%x�kY���֔	����T��xIT�B�4�6h
s	��O��B@!@ݴ��P��ͩ�7����'� ��CB1��j'������%y��[v�1�ɫr��o]���G`ię|^St�F�T�g�sz��
����'�/�J��pc*�2�ܹ���aZ�����D��� �,Z��B/���i��̞���1ˑg��݌P�d�����B���Q�_zf���kp���VL�'��֭6�n�KVD>��e������Z�b�7��%���(���hm����jT��vq��I�����wU9�����D"W|<8R;"噱����������c��Bv���0�Փ�]�̢�E�j9l�/��,of���J�K��Q��C�#ܓ�rx���뉚 ~����.v����ce�+0�C)��=� �<p[`���(Gޭ[�Q-胷J�E�aA�e���|����<^	��'�v+��Q��*�2��R��J�DJ��G��f)a�vQ���F���&�ۥ�� ���9T���В8j��b�d�&Ñ	 ��K�&��noXqG��cJm��E��7D�$�/���v���gc/Awj4E;��;�J0U�Q�	�s30�h�=.�����pW߬�Z��00�l�t���{�ͧ���f����7\����⁯B�7�Y�i>��ܘU�,��X��T�hO �luY��ԣYBU�"�E21����NV�n�	o����`�3Χq���r���8�-�k\}bC�2���"᩶aHe�|g��<��r]!�E���X#L0�����[u�7*i��(��G�:r�pBQ e��.�����*YP�4�30t���U￀�½�'
U�l����)�~/ 5��9��G�zl��n^D���
�R�h��L�w�s���D+���'Nb��t9�u/��YXU��f�v�W@3���$o���ͻ�.Gfۓz��OG��2�������gkm^��+�ծހ2���ê�|x�vj��^&8R:w��ϫP#�����5� D��L���%q�]����Q(��)�Yw�&�C>	��%W&t&�H���Q:���=b!oP��
�-�֑+�"�G( ����S$�Ҡ�$YNS�IBŋs{:YC��91� LMx@a=�V�d���76�r�3yζ�B�8c/؜�t�t'�y�	&�q�a*T���U*����/��OIcUb��!˼wS9�s����$Rx<!�pK+3�O��Kv�2�v4�>�q�nP��.�Z=$Ʒ��f	
�Ts�7�k"�k"�.��mΕ�����d��-Q��r�,���t֎���ĩU� 9���U�g6=�Ί�zt�^��TPMި�G*}\�5��.rƟo�5 �4��3#��s��-_AO~�Ft8�	FHoqT�"�m�.
���?!5���?�O$Rc
o���A$"�eŠ���kc��5_+˘����WJY����t���J�"�M.����M�\��M�&�����N�]\�5َIUʀOL�f��9-&�����f�I�3�w���JX��m(���v]I�Q@o� �!Ӱ�q��{��I�.�F���޵3��og�}�u�>=� �oq){�����i�F����wHd�����������bNH�g"���V�[�R�#ݤ6�o3�e/�6��m�]���.�� .	��S���eA�#Xem�ȑ5�[���Ş�r�ru��-��DFm�z|?���Ü`Ƹ
Y����M ��CW�7F���i�1)Uih���aCJ^���l�ߡ�X	�[j�h~T`ħ�A����w'��#�ع�xD4���e�O`��I>ӊ5�F��1�O�r3�f���� ��!�-��o?/�f�y�
���V!��!�	Uq@ScE�0�\��Ռ-�%N����� �k�^�Mn��DC-���t�>^4�_�SBYW+9z��q (ޞJ�a����x-z͟���X4�2>=��S�b�	=��'�P�0V�Ҍ�P�ڹ����Ю�t�
�^�Z}QU:��<��^�!��/`���8��Ag=Ԗ8�#J@`פ=��g��u��m4u&���b�LE��m�H����F'��M���pz2����d�GR�Bʥ��rgBYs�Ј3p9Ҋ�%��_T�'s"��6����J���v�$R�+��GF��>1}�;�s���T����X�����X�a�t����Sx�T�����<����-vt�|损������&K��fT_�^)�HB�k�����K�	H!|��{���CrK�
t��Qpf��+��#
6xOb�2#GոӵyWʻ	=W��� �o0�FKYQ�%6Yk(a��P��w���*�������%���~,_�-<�Ɩhd�<��a����g,_�?�cl��oD�RE��䨠Sd���"n�Y�D�wǗ4���`>x���ϡ"��D�=}��\��L,��z\@���Y�����6t
����bJ��yKUxs3%�m�D`֏�$u��S@R�g$u�a�z�A�9@�d�rA��I�}��������,y5p���.M4Ŷ[��qB'�e�N��æǉ�Ҟ,��E�U9��9�>��Fs��EE�Ŋ�:�E�I���3n�(��J#jX\����RAC���M8�Zv}���O�h� �a�X
�8۩��S�$�(ygr�Vё+��<qD�9��,��?"~�L�M�h�<<�)N����ō׳�zhxu��þj��.�9���;K��ّ�β���mw"�Qe��!`ᮠ�<�"�X7�a]�����zꎝ�&��Ұz�W�6'�� �c�{}F�#?�IL��%	ݹ��r���{�J%41��j���R�G��	�����F��3�����t�P�E�Գ��^����_j�b�"��aE�ӡ���Iv2	���{װ')�C��S�g�W��3��AZ�~ق��ư�����Ԉ чL��m�!����̠�$�il}'��{�m�`���t�,)��O(�ۡ˻b��ya�tuN	�N�x������E{"��v�u�����%���	�:"�$�$`j��hE��ϣnw���bڏP�B�u���]�� �G7�
�Qt�<T�~V(�.]�^O1���	��-ލ�˄J��14̲Y���@Ʈ�<��=�@� �玅��t��)
9��;�M�L��C�,4�̅�K�e�"����⩭�*ѥ_�	���t w�MLje�'�R�TT;A��jy�;�G�y퇊y�1�Hҿ���:�s�>�@C�s��5{1��f��#~
��{VWWa��?��Y���w���f���-�q��\�ya\f�
��r����d'���~A��։mv{�R��C�à�`@��c���7��MH	�r��M��qN]�?��E�[�,���3>#�׈��h��_�S��%����� 0�����n'6\�()�	֐)VB�U۫��L��?ڛ��p�ZJ�!3}b	������7���.��8*?p7T�A��)�� ��I�[+7Ќ����j�j�Њ]>EO�����s�N�O��Ћ@Q��v�� �4�]|�`MT)����(_���i�p�T��"Dà#;��2�;�G��4�9t0�ƃ��M���"k]��ǖ�$�>~�(���#j���rm	���ͣM�|@S;�w��V3�`��-��w�m�� #�J�գ]����L4㊪�q��y�w��c�w ����m�4�X�h8��̏*�&Ge����"��Xb���P����En̠������%)x�g�k&�K(�y��_~�������Yfƍ+�q�@�#��m��x��׍F���w��?�-�)�.��eQ�����8�JH&��<�\bf 3P�bp��;;��c*(0��c�Cfo��q����`������#�QN���)߂KZ�;�KZ�K�S�ٳTE�?.y}�QѯV�{��g{rӃ�Vg�8� ���;L�ϰެ��8Q�[�7u� �ʛ;��L;��WA>�bPj�N�3w����ֈ����Ӯ�����XX� \���'{u�-���#��.1�'�C�G�������nZD
�m� �͚��"��~&ZT����ivm�M�B������I���&��V���a�� ]�0=��G`	k]F�-ۗ!F��O�v�W���J
K�)h`�d��I?��9aW��V�2����I�k���$��+�s�t+�������`�O���J��J\����Wڗm��M7��>��\U��vGG�F|� �i����X�.�aW<�7���/���\��l���S����Zu��Hh�q)򢉅o8���@Ne16�ɑ��t�;~�a ��������)y%���x�e�%�I���o��6q�7�֎��K��	���d����Ι��v�u����"�>z�iA�\�zN�.�m�\J��I�_�m��F��m?�҄B9��.�b�q��Ljr���k�"wbz���ǩ.�x=4�S��/�1ɹG��'�B�,�z���,��"4��*�}?�`к(�趎+	F�E�� ��D9�H8|�<�A�/�V@�\Qς'�"�Q�\z��:�70Œ�\|0�aP��)Ʀ=˵�\#�C�y�'rE����o���'�L�k�D$x�p��]�9��-�$G��?��k�����)yC�
T=N�lpD��w�7`A���K*���1��@mB s�N]��Y����"��[�fCH<&����ͺ�.�ۢ�I�JTL1&���V�(�+��TQ7u����fi��������$^���
��H\���G뿌�Ґ��Z���P���א���K��0{���t�J�'�"���S	RЌ�`�����Ɣ�{�`�"�#W���w_ṕY/�I��q�{�5l�#���tj�W�Gw�GN�.kE�+`3ku�ɚ�����#��/o������c��ƶ+6�����J���og��YT������yJ�	��,���Y
9���N�-��;��Z�Hͧ�Īb�_F�V��u��K�.��O��b�������k+oK+�N�jL!0���l�Е��F��E#l~٪�VA�[�=B T]���S*C8"Rrif�y��U�׹	�����?���&o�L�2�����R���>��w$�?	/O���1�� ݎ
í��I��!�X�V�7��g�Ď�M��#)mBݾ�@5�{F?,�WP�l{'Pa�1�9�hn�,y�ގ��׻�iWe�r�7436B�)�9�z�l
/���s���FB��n]�� IAzQ�����;?b�<f���-��~\����*���4���P=8#J�C.����&�x��0.��g_
� �еw݁1r�g�-��l�Vq6R�i1g�0k!:��f�t�Kl2&�SJ*�� O�*�����v��PZ��b��P���7�]�,�_]�u�Ê��B����)bU.lR�j��>�UǝK�U|m�;�㱍]||;��|��[D�2K��e��h���nv�͘:vOͺ=V���k��b��9ڤ$����<�Mb�]jE)�0�Rr� !�x`l"�)�at���9Zi��a y���I���˸
�CQ�K�+Uw�Kl���-�����޺n��91���@r,�����Ug	�>�&֮�(��q��u=�W"���&pO�/.�K���N��}:�?u�ÔJ�JP��}�V��5������As�k[r=�1����ȡ�����5����# ���d��1ni�
�g���-�1��"k��d��.�}I�ڍI��-h��{�`�:K�S���x��]�����w.�N��c{��K]^�Kky8f�|�^����E�.}�;� ����.�%q��OÄ~�ӥ��@��`t�%�R��/�/�T�]`�tc+�j��D}������?G�kX�[���S��^�=�][Kz׌_؟�G����i���� ��=s���F=�R� ����l��箣&�stb�L��]��]�G�Eϟ�mQ<��T�p�ʸ�EǗa��W�!���\�o����:3�=)�c��be�bSѭ)���m���kn���n �{��l�p�HAjR�-�����41W���ѹ���� ���h�ewEK�\��/}�^)p^H׫ޢ	?Yko�Kr����B�ه=�����P�[G�Bu����(o;K@[���o�
9����Ƨ���a'Kj���.��>���8������|a���u�H�Z�l�Pz�����,je���;�1��Sy�/u��@��r��]iu�4���I!�Ic��5��h���PiH�}ag�"�Co"�)ï'װT��Sᗚ�%:;����t�66uΕ�"�`I����5^ς��3(um"�V�+�`���-�ݮJ���ʍx�����I���"�"���M:�ʧ*ñ��P��*�3:$��Uh��"�f)���Ƙr	�w���y��ҫ���k����T߇�#�� �F<6X.㮍�\��5�G�@O�B~F��n�q�\{�z�B�I(_�6$UR�a���gw���=y�	�d�9F�G n�p�O�J:ҹ����&�'���x��5�|�� �N�J�mn9�Z�Ȧ�.�9g+�L� X�ߎJ��]JV��������'�se���6��-v��>���1�\K�;3��|��`j�yy�p����][����"�l^��k��pk���	c���K�.���.Ⱦv�]il�ۖ�kYj%gf�+�R���[N��ׄ�s�q��~X�AcCG�'<����2������o8`��V���[��j�6��E���;p�I�Gty@����+�|�W��~hI�;���{����/S��,gZPݖ�}zts�ά�qM����g��%�)MQz�?m�<��LՋ����x }KF�P.�,Fk�l���W!��B�Sdk]b���wc��>��?��L�τ�;u@�c�����7L�u��xf��!t� S�?�-G+��̍C!v+��ۇeRYO��#pK�Njs ���b�<9�������~��p�>�����,���1��b�u࿨q��t��0��t��`��kp}���ɿ,� ��p�X\�� �aSM�/�64_(`r3�PfF�	�ѡ
��!�_o_|]�Z ��<�̣(ב� ��3� ݧ@g*(Y���ݯ<�M`�o%lN2o��MkE'�\�箆0IK#��E\���Ǡ�۩���f�,��q��j���ƌ�S����7�\�r������%�آ~*>��iy��;�E���y�p?rN{� '��q�3lUK���D9�� @7�A�뀪yV��"(�(D2z@��3����8o7'��8�r�a�L��aT`K$��Ч�0ײ�L%]o��}ʍ5ؤ4�`��M����#+��d�!�Ƣ���y �]��mc�bo b�����BUEw;(�����d�P�V��0��%�p�	G�U�P������;a�P�={�5�JL�녽�����]�mP��W�j(+̈z�6�)q��_
k늞���V3V+~�i0W�}���5u(���'ƿ��Y�����ʹDG�Ow9m�"�l-'��Eg�by�������o��M��v����^�QkY��cE/�{�[׏�D���X��!�>�e_`��ɄZ�z�)��H��)������^�k��wN��
:%������h��� `���%QFX�I���;S=ϣ��4��� h��h5����mE���h@s�
dY��Xc���YL�f�L�h�}_�B�C�y+��i�����vo2�5�g�����*��67��NZ"�h"��q�0��2UO~t�8��Q:-,����G���c��k��q�O�%h���f��(|M�*az��#�O�4�1���kq�.|Q���/�u���n	�4��;�ʘ\HHu�l�QdO<�m��N�Y�>T��Ė㫉��>�2~g�&�3�Cl�EV��S��Pd����L��\�9��z(�[S1�X���6�ϣ����&Jqi�!4��ݡB�w��i����Ŋ�f&!���b�d�1�i�7�g�'��Q��gG6�G�����aV_�ʃ�q��QM����r$K@�oa=�?%7�R�y��m-�$���l��mc�;n������\3�k�ӗtI��Z"��[�wq��D������ԯ��YVܮ+�l'����jJO=GWO�;��\4VF
���A��l�2M)���:>+�H�#�v�2�k +݌5s%xMn9r�6�2V��W
&�'%��2>��pG��V�n�_��I��=Dr��ͳSHZ� ʛ����u�ׄ��������/�*���)�P<
*EĚ�ηȑ%�ߺ%�������-3f�-��G� /�&��l�X!	���lNn��^5�	$��4;��P&����=8a$����r���WB��L�no�Ү��B5�i�	x�IWj���������Be�\�t�J��~ڢ(S H̄��nǕ�?���L�P��u,0�S�~���K����ğ�O�1�D�F��\b����b�&�{TA�Az��7�;j��}5S���	VHM��þ8Nt��T���f��e�Z����e{�l��~w�!*�l�/�=t�L�,n4�s=�@�F�����Oz���W����Z�CT2 9Yұ��Caksu8���cIH�̇T<%�x*�t���P ����q� ����r�E�:E*҈P-/x��f��&��p5[����u&g�<`�s�[�K�-%�+@�WX��
�u�zp�7��
�jS�_�J�v��%�9ߠ;P-�'a��*jf�"��Ë�t �m�d	gg�b`%�1���@�
���g�ΦG]j�8+nJC1_Bk����]��G0�lu�Zp8����;�זӘ!z��4����tW4�L���\��Lt#�fk؝��W��x����7�	����S��c_�a��V�Bz��V���:U����a��� ��x�vg��:ւ�'��u�A���֑B���{��ψ�e�����ez"=�ELQn�n �N�f`�=l��*�?�X�����.i�6!�bu�e�3I��7�d}���MUyߪ'��P�rd�2���]H;l��I� �U^����t��$̠*I��ȴL{��#�BڠlD13�������8����iR$�^z�k�4���Gu^���E\��Tqr��D����'y�uqh�o��5��I	��%�I��;�y5[�[w��cc�ѭ�)�i�X��F6��V5�}W���)��(A7�d�y�̶Mt`��خ�ߒ��[i߿�����d�v�#��v�B�%j�Xd�j ����4�m,a��I�&��䌱�ߴ��Ǩ�G8
��'�2GZ������@��EHB	a>t}�}9��һ��ѴE��^p���I�B��D*�Hޥo�Q߰�A�NWa��ۂx}4"��B��b�#͇n�%���(����փ�d���,jU�+�ٴs]!����v�%����3�ˇ	Q�ذĤA`L��"xl��9C�K:e����F�	d�� x2�Pρ�G,�Ν�WQ��W�F^�P�oM@��}
�N��( ��n3QE=���>�ۜ�}e�M=�隓��� �vSRUk�]�%)�%�-�.|փ�1G���v��ϰl{��\:�Z��ZE��9�[���!�i��0� �f�3��ү�����&�)֤_8J�ܪA$�Q�ד��Z��R8}����U�=x�.��]��?�Q���^Z��udHC0�R���^X����=�o\7���g��l�����SdGh���/Ԍ]f{����|$V��A���n�}���;x}Y��`�Z��Ĩ��{�� ���0��w��*��|q��fB��k �v��@�=���Vl��x��찳y�����,�i�s]şP�[*i��2�Q�:�q�颾]����):X�}�~b�s��b�=i+�q�C|Ѝg����&-O@��kf>�@90<����kD�F�"f!�A��C��������d��ٛ<�a�9�YJ<�(QN��;D]=���Ƌ�c�;+�q�Rdڞ�%Є�ͷv_纺F=�j�d���X��K���f����r�7�����#Y++>#7Z'E�#v�ױ����F�}�	X|s�c]��)_&�ЍIP 18=�`������v��h�]�/�M�7$�P��j�{���!���|����<��,���]~ɚAi��*m&����ɥǧf�����fJ�C�.�C���W"j58����)u����
*�p���ޘ~S�,n �d���\ݳ�ꥴ������@�0�7�~�W�U�i?�(�6�иiB��	��%�X���e0B(�)�X'<�5�s����|�=�q�1-ȡf)�}���/+��HH��6�7_���epf�f�����4	dzG��!"�!�����i�,Z��ܗ{kp��`U���S�ؐ]�D�:�M:�)�����fG�ʛG�#?ʥ��#�wF�/��
R� �:`�g�8l��yd��k�.7���k��������SЂX=��y��&�)�+��E����_�Ϣغϓ��D�٦uƒ@�5�UfOA{I.��w�����8�P�$�N�5�.`���	d���+�����i:ڰxtUrڹ���l3j*��k�SԄ��TG��9V��/um|
	�Xs�ho& E._;w��G����
Ó���D���c���!\z�}I:��r�e�}��T�bC>�4BW�ux�[g��νkh�:�\}�9�*ַ���2588Ј^z=sh���sy�U�n��?�������	-2�l�ʫ��)�xi�WU�Z�HOtL�u'C�I�~��n����g%ù�9U�Dr����s�`���=� ټ��75��Qcv{u9"ɝ,;�։�{�pr�oF�����tg�PE3D��hS�(�&l,� L�ޒM} |�F��LT"~�>�F�Q��q��,T��u)?+�p1�ǧn���9JV����3a&�i��LI1���c�s*�8�	��v�/nѡR���9�c�Z�XT-r3��p���l�5R[�%�z�t��%�E�FaO�胩����:o<	KE4/@�EF_�����<�ݼ��yȜ��NL2�K{'����N���}v�&�S�Np��!
/,�y.5p;��?�}�q��oG�%���:+�䥅�u����3Vp���]b&l�l��_c��|4��=�-æ\�z��� -�U��c����xO�(�B�������7~�{�tE|���{x���Y�:�z)}Z*r�����.�����Y.-dь=��$�fc�(Mۣ�3�Wxj'g���w���Oi����b�w�i�DP��뮸J�e҄?;����4A�|0͕�>�'�]+�b�OY��A���$F;Z��B��Z� �|.pЕR!+�O�SrR�gV:�	��m�J��*V�^V�H o�:0
�`�*���D�Cbf��}I�ɵ��h�m��d�Ru\zuDc�������o
+�"��E��}�AQ�Gհ
�RJN:�Ç�"���W�DA�! \^�;�x�7��ɷؐ��h��m�.Eؒ�۠�:�����H� ��^���u�FDf��8�P�B��`h$�U8(�H�Y���������o�4��oE'{c>��k���C�8�O�%�֌= d�
| ��P����(�٪2�K��,�?�����j��D�R���
��������h��Y�voge:,
bz3x9�r�����>9A��'�G���L��}�����A4c����OnT�����ۀٺ�\�=)���5��6`jS�O�5�su���}�L�TE��o��!̘��m��c��T�8�9�NL�Pݸ��Ϻ���p���\vS�R�1�lXHpUf��Hph3��c Vs'w�Ģ��ˋȔY
�ʶh���]C�ޱA&c�+��R�%�WپL-����^�3)w�:=��T�}�3Q��Y8;0��:j��ٴ �&��xx��s�U���o�ց�_I8�l����Q�*��E��>�D�2�yH�#(F�RΥ�5�ޥ���v����7@�GY�|K�捕s��D��Q�4�Ii�U�d�������Q�AE�BU���w��P�&��d�����ضj��՝
�j�rI��R��j�%>"�o���
�U�G��5S������7XY>08zhZ���q7b����B_@�wD}�I1�m��EDD��q��N9���>?���)l��Elw#b
Rjq*��"Ώ���u�8��w�F���q������g�v�&_�'r>OMe���n]�&��R��]iU=m�ڃq���7�n$J�i�tF8Iԩ)�Q��S����ľx~�-1��H��A��}0�3fp�=T)'V�Y<R��V�I����f����x��I��������:�Wd�L���S���G<�dJ�b��M��D��-�ơn6�q��x�I!�>:zE^p<����m�sH!3Ǜ�e�!���>%e�'�U{R�E�ʃ�؏iT�$�I��C�Y�=�n���݃���Q%�Qs����.�ѹ��j��S�V�;��\�]�j�M��W6�AԨ�|�H��f���ǹ�S��A 7��"�zX��|��Rd鯨ju��׌�g4NTu@�����R�2���!r�I�%����g�����·�k��AOZ�;�
�]I,�GL����۸��|�-��V�U�v�D_��� �Tb�P*PZ�k���Y�'��Yu���DE: ��~�?�+�E���3�Ñ;n~Q{X��m`���s��_}|g��b��+4��ʚ��E�*}�F������ ��"�"P����ܡ��Z���Ρ��gbG���௨��l|D�w#�����ٺ��	x�d�Y�b�Bp9�aRv�C�>�9��&��(4 #Fڏ�L'�Q�����@s(	�0��q}�t���	!ɯ��������Mn?�ޏw��DB+N�y�#�O��������J"K7�ZaY�5Fj���`�h���]��'�0_���^��&𖐔����hWg�J-bx�O&�'������1���%/H���&��!�wj�ϲo���� ���x_���
��R �i⧖q+
�Mt�
2ja붌E-H.����ԋd���V��ؠ�3�� �?l���BNr�bjW�2!�/ ��몐���EE��\�n�G�pq�ꦅ1sy��e�n��b<��h}B�������Y��) "�b�qʰ��e�;�a���u���y���e_��u<9�d�FA�������y�Uߏ.�m��	,E��3����t���ԋX3J�$c���9���B��h���s���Y�Ζ�Ô���j�-O1[Ό���Ml)�H��k�I3�5X�6GeT6��`;P:��6�c�襀���H�A����?Ƚi8�/>!������=��r�R�]���#��mί���ĎmR�4g��"G����ֵ��b�dB�owWM�������i/���rZ�\��VS��ԣ�v<�1�+������c6�<�w�`�zVu�̺�����@��U�;ʿ��@P��Nb0@9S'�h�Z�;��V�r�]��D����E��	CӚ�3��hR�R�p(szG�nƪ���� �.[?Ѭ�������6B���#�����k�#���K��Rq䚱��#�+%��nޥxYSx~�>����r�r�=�ӆ����r�9q��эHF��8��创;,[���r�k�pz5��^o`ݶ
K�榲Npà�i�\��jכYc�۰�,�y���&�q.�h�T���m�QЛ������eJ2�ϦP Ut��B�͙���4���#�۹�Z+_)�^:O��!6��_�x��.I��&��ݴ�LrN�ki ��j���/GQ[����[��6�8����윙3
�>��vO������mj�m[�l�jH��)X��i��;����� �$��,�����W���7���h�,W����<�
�c��>��'O]=%�=7�ˡ��(^2P�"�Q%A/�#���h��٨]b�{���R�=ø�Ez�S��B��m(k��̬��R�g@_��S���/t� F���3Ik����H�g
(�8��i������C�������~%W��ι�g!�~�!��CI�n�W��0������� }�7���3Y����Ws�J�X��_�n��P-,X_�@� ��ߑ������R�#4;�� ��J{Dy�D��lb����]k����kn-�2f��J^:D�_~JX��.[�%1���y�G��(�ur�N;���+L�H�7<�zr)���a���r.*�
�V4��Y�3�ӈ<��\[i�K��xzyJ2�y�Nd�"�9��	��zg���K\���n�Is�~���(Y��]�nή����*��ioD�f+�fS+��ͳ~��ܮB��4��3�Ӗ���_����'��k�r=���1�[���&Y�D���6ڬ�!������7�uU�~�;�y�(�A�Zh�C�1�=�r�&������>9�:��=�{T��Q�!x�	�c���Ru'J9�ӵ��ezE�ݮ���R��8
��H(L�E���E[Btza�<��d�Y��<ֹ�,ݰ\�� ��d��%�IS�ɧr�<���Z��h�}dj(�D,qR�r�蔋)*.��i���$�4T���1�+d���� AK@���"��.�� 8IHD�;�"��) �}�+g��&;-+޼�!!{W� M�z;*�ߠ�9��@J�5���
?�@j/4Nt2�U����3`��(���&'� �*Ea$0K��b�a4dʯ��O��*���!ֲ��;T���Q6p,�w���h�Ye�L�X<?YsU[���KR[�싑�^*Dũ/ӎ{:��8b}8ZE�ZC^Ec�y��p�\��B�>�Iw�6�Dd���]�0�h��,��2z�7E��n$7� 5�X�oY���p��Mf���鳺Ӱ���#�q�:Zۜ��3W�:��t{
��н3�gz�KY`~��FL�6<�YDr�] |��o�.V�"%/A���,c�[TM�jLL�X�|����/(���?b�sJ@��nv`��Z$�mW����WƸ�P�Ԩڞ������|]c'�קz�(w[��K�lߴ�ɓ��ܜ� $E D�GOg+��VZi�p.r�`"��|'���EBjDB��2� �W�t�+����oso�I/~�;d�`G����)��z�����E���
��E�k��L��OB3����U-��T~1��d����':e4,|�$���&u춖��7~�M�}<���pe�la�"��S��@�Y�,Vhf��y�w��u� ��
�M���h|?J���p�TM.E�
��*����?�����S��/�g�cqޡ˥��=H��Ys֓s�|œ�f6��݊��ם/����<ũPVdbcZw;�y�U��}�2�p�F\;�!�y�\x[�5���S�$uH�9����4G��r�*F��&i���3+�_0�:�|#{7�:�S*O��iuuR�)���1g��W��MR�o�G#��Ü]���U3/�6=b�����:��9��x���%�]�<�Ʀ��I͛��;;y��|)�P�{���ԆWQ�ȡ��c�[����I�]��"��P�`�7��q֩��|����Wm`�L�Wb�G��(3���I��dXB������c���l��sv�JGJ&����K�Mφ��D^kM�h��&���_�
�u���T��/� V��,�X��Ea�G�^���׶w�������t��8F�i[}K��h��}�#fl�xoO�_��y�ew��$�*C�|Lx���d:d�;I�st@��ܿ���0�#�M�
@Qe�J�.����pnC�a�e_$]�Eﴡ01�C�w՘]��*C�EQ߁k�4���>��&�ss&����ۻa��KZl1��ƵZ��y��6. �A��{�Ք@OH�)�'ln� N�����b�б�$�����\90s����ֳ�M��Ո'	���W�l��:��;jgb��L����G4e�M��B����}Q��pt1�f�C�>���0s��.��ט�x��f[ ������ƫ�U^��pb��� �b�"��������{.8���:�����b� �=#�N�D$|i�'��I�h�wjǐ�ܩr������O	�;��o�����JGV)�J)��?X����Ø�!r6��'���f�j����H�=Y	�%DZ:�{Qx�JyR�Zu5[��VcN$�@M�_(���2\]�Ғ�^^�*3^�>VA�\�o�=[Fnu�4X�G0j�'�8�n�Ş�}yZ��8�Y{Z����m�	�����v��w�s�ג�-)4&�%$�L�婗��r�h�����������qibȀ����k?l�7����g�5&DWm��>���h�/�:d�
���S�y���"jԟ�.ڐ�}$�+D�1�����:�И?[�P}�S��ɰy_Զ(� g�i������IMu����m�ƥ�XИY��Ő����(�E�|���@巭�"��d��2;�߳S6���YP	�@�^c�����8�& 	�+#ߨ񯥉�?��0�K�=�?6`l��8+�OKL�	N������w�|#���{��o�s�-�˔�iv��<�ɓibܚ�'�#)��U��ԧ���h�'���f��,_J�$W���֚��C��@����*��2p�$�F �;����Z����	Ο�<'^˵�ϓ%TJ���T�0H���:�H@px�h7�!�Cu���Wk�zѽ�:"k���"��b�o��ؼ���o��D�'��g}��(��wc��W��V�E�� �����F�	9���]�"C��=�6��N�x>���Nږ�_��<�f�����y���G+#���%X�@��0�Q/��N"?0?����E�!�lS�r���� V�Iv/����q'Ooi�o�T�[UsS̕��p`vT��t����\y�c���nԺ)�w&��CL��V�W�[JXeA}��V��R?�#�y�������U���(��K'F�_
�'eƣ�öʲ/��)��������Z��ͧ���k��k��N����~[
� jP�Biz_��O�XX�d�Mԓv?�$N,���Ѿ�xx�Gku�Я�C_��T�f��A;�`t�PtW@-+o�E�S�.~tU��8�t*�[Q�-�4E'�Δ�6�c�Ft�N�eyB�v��9��w����&�+x@+�$���
I�y��+3��hj?q[7�o|*9��⭳���ME�B�g���H��W���8����n�Õg=u	��ȼ�~�4yj�tt�p]9���OO�zi����:��!s�w��X�?��-����: �����,Ȩ"y�+Kb����µ ���6��c���0��f��&��%�>vz]��P.�������a�+�C���c�,,�A	�E��A�I���&K�d�	�A��M6� ^��f�'�i�v*KD���Ɓ��6�v�{�S�x�DlD$�� 7��@���1����^|����M)�ɶ����K���jc�S|����aC'�^*_聍�MYg'�T�FF�m\l`�چ����(��>�[�X&o���pT�F��4�-f`��JWl�����P�����4��eҥ������W+�*�>QР%�,�͒�Qj��T����A�p��z�^l5�᷼O�݁�/�J��e��s���v�8ϟ��G���g3��jIb�t9��*�gFSHYB�[����ʑ+|&pҍ�����l�N?�2���Ō!#?��S{% ���3���G)��ok��:x}�#u�KPn:&�H�b<�6�l��T�#gOKtk��ԗ��B��cj##��f_��)�E/iE���i�O�j]�*�=#\*3(��UJ�<с(+�9�G�, ư���I�3��������ҍw(I9���x$�"�ڐ�
$79�V���n/ �����?~��n�=�z��w��+�SF�q S��|���!w��֣$��.}�:K�.���2Ư��o�?�/��ϓ^��.�!<Ф�E�Z����u3 xpoU6����,l |��D2A�XOp�W?��/'�}&^C����V$���Ț{��"Ƶ�0�)�|��w�y	-�5;����t"��Խ��UA |�*�v��D$"��6<���y�h�h��R���ˋ�AX*2z���L���� ���a��3@Ln��݉\4�$C4��k��s��K(�ߒ�@�L�C	B����f�+��Dq4�q�9�+Sf�N���+�p���������S�y���A�GV�`K�O���(NSJP��|"f�SF�}���6(�3
��!�萱H�!b�o`�m1���hE�N��:I�r7�d3�Ayg�`!7	�|���R�i�G
S9B1w0����� ଗ����ӧ���t%Y��/F@�uM���3�@1��Ci�5�E7�I���®~�@��c��������.z(�Aew��G�Юa��R#�A��I��u=����Ot�Z����M$�^x���⨽�Fa��'�n'��*���	��k롬�"|5W9::e0Y�� � b�`����z�b�n�w��SFy��Rg���f��Y��*���)f��=AV ̌�:&�D�āߙ��<҈��|@3�Q�G����2���U�em�={Ґj:V��Wq�k��N7&�D4PZ!=Dg�@�,�����v��@%�"S��Ϗg��;6"��peÙCU�-d �ϫR��|d�w�2춃97�`�B�O�T5E���q�;P�cB�����BB:88DrV틡�^�+��m�m������r�4nf4��h�9�"Նj����k����� �V;�{�@A�ll�W�vE�eR�h���ʭ	�Ѵ�Qv<��ڢnx���v��*?��2��r���B�6�B��]ף)�ɥ]n�@�t"IRo���ϲ�,���p:�r��l�{�4{����2�;����<.�k�c$��a��C{�=���W7vK�)�w\���up�zp��А��]�	��5�M��I�Q�:]M#�U�'&�7*��������Q�x����Q�2Vb���xؾǺ���o����m�r���&P��t�2m<Xg�*a��Uv3O�CV9k�f/l�A�W\�²e�gpB�(&s��!���Nd����-��mfOH&���{�<}���=FC=�7��$OL�����Z:ɠ��v2'�t�W���:$���jly��>4����"} ˰�vۤ.�.g7t��!�z�uA���tڔi�QL��pQ�(�q�8\�\��F��? p�� �'=C���cH��ݶ?��	�C�Y��=��I�Y������T���\ǆd���#�o�aM�ݧ���Z��O�M�l���b�)�߲w��?A�&���+j��c�{3�F��6So�6�r8a �'oG�ސ��R���B�qT�����HKJ�q4b �����4Xg=�����C�A�������7u��L�ci�^%x G�j{�?c8"%hx�d��y� ��d[���ڙ���`��U���g�'���u�]`U�7v��`��`��{�xB����!~k�WT�P^�H�	>�#�-=�7z�^��D���so��c��9��^� �CYs���!�(?�_�6h3ߋ���Իmh����i����4��]h��?	��.�5�C���}�CA�)<��d�s�V�Q�ׇ wCx
�e�3�j6���n��������D���ěĤv�!6�1��|]_׬����@#�6Y�힆��<�V{���R��߫���,'Ɩ��8�@�ETN�̚z"�!���,Z �E�o<��]Y���%V���X/z����<�e�*���TşI�فgpa�[fx@H�Оs�Ҩ��#��Tux�y��!���q��'at���r)dW4,Ё�"%f��qG��G�N.�7�rD��c�rDJU��8Ĥ�Mi�B<��˘xF4%G~����䥧�49`���ݕ!��ll��<-z�����f�r�M?<F/j�J�m�r�h�ZFU��ط���f����
��^""�(ћo���V��������Q��q"�U�D 0B�G���^!{�v��n~r���ιs�)�,�G�2���k0����V����y�@W� ���������Q���\-]$��eYT'1A�,V���A�B�[ኼ¾�bǬ�1+I��G��5'D�}�^�p_ܨY�!�^�I�'����Ή<F�O�����޽�1��8�_[�'�Xn~�|[UОi-���?߷�Þf��C.*��L�1A����Rz���p�]�R`�<����<Q���0jc��9m&�"�8���4��{4ga�����;r*z�Z4Yp�Q������a����hYߟ �@�c���H�����>�ӱ���k!�}:�	e�?J��s�V�&%�mgq�҄�ϴ��QҰ�ˆIJd�g'�#! ��X����2FWW�����뎐�ɺnᏯ�����i_-�^	�^NK]��p�_�Q����bZ�\�J��]�q��YGu���u-��ͱ6g^��[��'�XE����Ĉ�'n�����W�t0�%�f���$���?� ��T��D��q�|$F2j��}=X9F�e��Y�Q��0�*�Q�£�0B���"��w�P2C@R�{.�^�u��~���4�#���S�t��I�U�P�$o�^�M���@t��N���=��`�#"���b(֧�܃���6�4=naj���u5�T����!Iv�o���Z����ƅ�`�d7ଟL�Ӈ�s#t3�?W	KCq�j��%P很�CaQ��+�t>>�]\����lh׌!�_S@���	l3�UL���f�)�$�)��؊y���6=l����Wh��dL�7�� ��s�@��٢� z�BX���)�0���l��x�fT�'��.-OEKt9c��M΀����J� 4���0����n��k�O�)��_�V�����\����xc��K���Ge:8����?j~�Q��x�~QkH��z�]l|��G1�Q%<���ԙc�U�qtJ�(�4��-��1�$�<댅奖����)��ĎA�j��Um���.S� ��_�;����K,Ө�f����d*U��m�8�Y�����LpD>�\E�z�l�k��L��.����>�źc����螐
���C���/X�X4l�\y�&�P�������0��D�|L�-���������l���E�+�&� >p�Rt�^�➋��X��A��>t]�x��P9���Gl��-6�Rp��&ay��$��Cܬ��W>�0���{��^������e�濣�>\�e_��[�����d�YT���߀��jzI�*G>���p=ɯ�k����12�B��h��/�/Ksӣ&j�Q�����Lut��ԥDD��,2�:}��Yy�dF�����RQ���xs�nF���G���
/�]iK���9���@�Ԇp�t�D:~�Pdɑ`|+:P_˄�;���Ҝ^Y�����8���W֕v��#�쿀i�mKɅYW�UV��%6<����d�RO;m�?�^e�M5�N���	���\P�n�R�t\2�x��N���>��Z��#�i H��Fxu~�$�W���M�ii�U)V�Q$Pj�����8cJ�4�B?��40 �D<k��!�Ct�U� �3�=�X�@�&WLz�GyM��n �� �
�:%�@$#�� �Ǭ�CF��m�O� z��Ö_�#x܋>d:'�4;9�7M`��k����˝�4���Jw(k�qx��&��ͯOj��sw�����/SۦS��4."2���}e��G��ӷ�g�:e��L�\=����}�kL#�ʯG������դ������iE���_@0�-�m�"X���*�'�3�_?8�;TO�>�&����{��?>�f~����e��OQ��Q=�!��dm8G��ֳt)��,
������dRV{|w���~�"�2���Q���˛i1���r����UPD��m�)ED-Zs6�dE;5<�P����׶4���!�����ZU�bۻho�ֻ͑���OqU�8���[�c��]FwE>&mn��s��P<EreE%�B�J�fz�	.���+��>5�1Ka?�9�\����:е�,yz�e?�j4��sS�
��<��MY�1@�D�#U>gIϬ�8"���H+�!'\T��`�Îh7��&�C`.z�]zq3A��C�(x.m驌��n����1L�%��@�?h�ךƤ �ImE�u�~��9��G�~e��j4�{C�	��r�ɪ�E��`��vT�ra���=�Z"&�w&2l��\��&��y�����=�z�X�Ma�����
��5r���&�"GG��萊{j6����9����>��8w`w_|����JNؒO.�D.N*ه�N��;<�7̄<�u�ds&v�_	�Q�v�P���6�^�k4q�<4�_�u'�o��[r�+�{Zq�7n&R��᝔��giJ�D}Va�Yr	I��`�Z���e������q������X=��+��l�zn�2�,5�A���
����OJ2ц!OL��A �����O�t�&N%!��\�%z]�w�>B���m>�^�r�RUg6��N�T�?8V����G�l��<n�4�D�����$Ï��H�U���FJ�>�9$ �ś]UTS�p��������l���.u���0�e��m���&ƪfh�q^��I��/�~���`>VV���	�>�ݏ�|��z�Ȓr�Y�肜���b�e?j��b�<׋"�ޞ���՝x�؏��遹�sG�)���(�Ã�1R>��;n���w�f��Β��!���.m�m��ѭGe\M;�ku�~�seA{+�N���+���<u��"�I��tw_�w#xr:��W�k���{A�̦��Ћ���<1�� LYĞR��Ǜi�񒫗\�����b��GX��%h*�t&�1�`,�S�p���E�\���U�!����r����a�_���p4(RJi�ߑs�U��uE79���d��O�0ӛ�tR��S�,~�9KP*���[���`��<�g���
Pe'(�ù�����OM`�Z��n�%R[Z7���94�ɭb?��7����T�!��*2i����!���BҪ�O?�P܅�Ouaͭ��!!�8ï�L�T�N�͌BkԨ���w�5�j�˂>9�Ld��x\�Wz�6�z�0�~:�<�����Psú�Յ(ҳʎ�7�YxO��+���:,�#���VI��Ҋ��vp�B'v�(�ȅ,��w����Ă��Z�)[F��L:/2w����������έ,%�IJ�Je��)���x�j��:���p��p�Bp�E�V7��ZuOP�>�� �AIx�ȗ:4����#�����~_y��Tsq�0�\Z�>������\>Tr��gE�_�C`�mǢ`v��}�h�f����z����HP�'�v���1p\�P��+7�k�;�䨘=#��v�W���[�G1��4�(�Ob�ĂHz���LJ�(h�Ͼ#/B�*�#���N-i��@i��n�o�ċwL���SxK8M��f�ޞ�X�Z��������N�}䀦���C ������F���Pʹ�[��	��)k��B"���M�B�K@�$�}=BA-*-�����5�E�ĉӌ`[�NR�(H9˒[V �t��|pK�u`���Y����J���`����'.K G	eS��p�����H�5���u�纱jj)�������'���I"Dqͽ�~*�*�œ��fLHM*���I��P�+�g�沱`���$�t�+@��)}-:|{@��~�s���g�"n)�q&�LCa./0�$��n��X�z�9�=P��;&N���#D�{+B�
�����4>��<�Zɯ
h�����}%�GB�f���HD�tho��t���	��C�I�9f�G��:�(α�n`��|�B��t�����c*�sc]���=�N�[}P�'��GX�&�U���6�� sq��r��;�(e��+���1Ŗم	���a��]�Q0Y1��ֱc�N]��M�М�.}ԋ�y���?��Q"���w}3�($b���с J,m��3�1hv�߱����v���{ ۦ��w�~r��x�JV���q�*ٓ�2jſ��NƲ��ʰI�Q��������gJdN�8}̘����0\"C���#מ�	�L������ґ�5%@�y������.��K�Y��v}?`%�#�4��.��o�a�(wC���
�E!M�����fָ�05FhH��J���	��+���6��LW�#�-PY6AN�r�Y;'j(�o��z���:w�ш_����?��{����;eqH��Ћo�k#�,]��=U�f�J�<<���\���_���V��I�)}ŨV��� @s���~�i���Fn+rڰ�T��xxpK�F$�b�1�.H�8z^�����B>J6 ��^�T���`1��>��e^9��$-�H7p����K�F!wvd#�W�5�k4�J,m��M���qC�e���qD���KsXqϑ������
?�=��i4��V|v]��*Nۍ�l��	�G�v��.�rw�Ioe���s�7/n7��s��Ff�F������ϱ
�y��O>5e��,P�06���p����a(���s,�TUķ�;�h��f�{��j�#%�2��"����!t�-[u\:�����͌��0�.��L�EHa���������LOKA	^�7J����Jl��5B�a���_��v!l����.�q�&��/ٱ�*Yfq,8��M�6��N�z�s���i�5	�$2��vnƬ��[���o{�n��$1x9�����v>���SΗ^$Ն<��D��b�.v�p)�~n^���yN�r� �hp����*�s}��� [��3/��n�R�$M��l!vG��U�Qr {-칮+�Uז.փ��Q �29�}e��N=��0����V�`-�i��k�D��c�Ix�@�QS�8*{:Y ypf!B�=N��^¡ �.��@�����; ��/����q�|l�8�*� ,��/%�
۞��f�z�������M��D����*^z��$�]i��6ң^��)��<�aFJ~~O�ԽsY��ء|~�$E�+�5�ī�X6�}��h�.G�OpA��y��Qg��3�Ji�D�NF_�3{��#{�[oɇ�S~���3�W�u��m=�|<��:�)f�=�12/ 6b_{ز"��!�;�#�J�'܎�47c�5zbOJ��Q}l���=�	��M��Z� Szi2ͮ�;T%z �M�f|1~��g
*a���Dm�����T���h��!�rQ���,�����q�3PΒ/���;"�
d�N���%K��=�傮��e��TSC�����{��UD�����SM2��yDPOI���K�O<���̦��;��l\���p䭂^����=����{7����H��5�k�8�3���p�%D���$���͗	���w7pE3>�<rD���!΢2u!,u���/)6�x͡�w�}��2`�+�R�U9R.*�V�x��ol��g�%;���S��~�xI���_]��X����',SZ�!|@㊬3Ée=��UY�z���ٹڲB-��9�#1��r��_�Fu>l�,�<5��y+���<��QQ�E�$�hbR���#�������)���q?<i��h�b �����Ժ{=�F.+?��U�ko��c4���=2���s5��5�R��d��}A`��Ң���S6��%T��Aډ�γ� "}��
���u��ѯ��.��FXf��
J���7��/�#셛*h���?J �z�|�qk2�EX roE��� ���{�l<�G�.Q4�nf����f�
[�C|�m9�/��7PNb2D���}�(��� <�
q�/wJ#i�̐�h��*�:m���W�Ɗc���#p�q�$��<`�J���;�6�IEd����D���(���`dr���9� �t[�z��X�U��QXk����\�d��Q�7�څb���
|�
����ʤW���Z��P�^��y]6���6@%�NX�=��2����B�(�12A0pĊ1���ϴ%a���.cP�X���z��!_�H��A=�X�:Z�@�͸⟶�X�fq�e"<!������5$k�ӫ�*'�]ͥ��x]�������j2c���|��D��!�GͪPw��!��6Tl�_�2'�w%�~�
�o��X݁�D���tb������רW�&o���ʄP���K���H��C����m�dTy���o#&o�1�v��J-�(&i��M�f�P�>��c,s�Ws�8�R� !���/���SJ�e��l8�����Mw/Z��v��O~.���K0eIv�������I�u׽��Q�w�`��;����<�wO�\��G�/�����exצ&����
٧^�"����n2S&�mn�%�5����)�[�ӂ�lD3�`��GB[�a�YX_;l���\�<�����%Z�����bW�T�ЯvU��W,QQ��GHkG��,��FGVo�1'�K��
Dn�0_�[z��V��P&����E#.��-S�LS{
�wr��3��f�l$VL3��2�m�T@�ā����B~F:����q'���e��S�!L��u�T���|g�<������"��U�>}(�C-g^�t��-'1eqD��.)�䗦mmvL�$��m_�-(�<��i��
\Y*`�Q�R��w)����Q�s��ڑiiВf�(��ls�̫Uu�8�0g��Q�� �����:+!�+����_�Jo�Z�p��*6�(֭���G��Yl��m��ײ��#?8H�/ޮi
@���͉q�{?�Vm!̺Y�i��$"��{vF�g���m��"=�ޅZ��	��F�t�ӟ�J�8�xnz@��@+/Dƒ�t�=/0�=
�m<�����4�L�)R/C!�j����L��Ɉ��;K��F�NǿҎ�)DF����2�Q�r����=�`&�U6E���:3W\�lq)���]�F=�W&d���mީ֋KDA�:��aXF�PQ��9S�A��$I�SΙ�۰�}S&���:"(�C�j���	uHL��j��( ��!�̽e�7�L��T9��vkB�J�ϒ�Z�@��:	3nw%$�^�s<�6r�(�[�>!��"�����
�=��6�,������=��]���i��ń̽�2}8o�
u�V����f,!�_�n9�n�N���;�.�-�i�}f�|\��z��T�y����CB�3���i{ӌO����-.⼐rAhT�(���gl
o�g�J���.�Ҡ Gf�l��Q��ף���#��)$��֣��jFd�U�:sP���1X����Sf�em����[�!�:X'��~��7�y.:����ͻ�yFӻ������o��b��z�O ��Yo'*-%��{�֤�t*-��CX���� C�@v���гd>ԣ�}i*�V3�T"�?6_��]�t/A B�d��T�$�y;#P���bHe�%X�zV���K�Ȏy�Vyڹ�J���1{�'��#�u�8d0]�e|�m�=O*���g1Vᰖac��4�"?&�gӆ�o?���mE@B�ʩ���Y N>����!-�[&��*�a.+V:]�rp��L��g�,���\�s8u^F�\U��_�kQǬC���t�F��>論4�<bmR�����<���k$�-�[�K���_X���]��0��^� �ЊS���	$�wЊk����`���@�mqҏ������>��ÎEcd"Q��Q����W��~~o|�� ���|��X�I?���'�n��o��m�6_�Gwͫ�
g�!�Q t�R`�N���MG��ߒ>EL5�05���P���|�,�nb/Ƥ&�9�;�s����-��B����^2��U�,�iժ{9FKl�-��uh��X��=��� 	�1�������k�h�Вm�����	}Ws�V����{�>��e
��x�T�UKT���_���Tٟ;LO[N�v��&��Y�X�5�=�	=�����8<��L&��(��E� �M��e���iOį�C�Z ����F�v��۠���.�����
��u�R�a��He�-\4-o����!v;qo񟍔 [�>_G	{�R��9�4��	ao,�6�G\� O��N�l��(2g�1��%�i��٫s*�S K���b����V�x@�&��\qU��s�g�VΓ#_gOֱ��K����V3|�_��o�|�^�sg�1�Fx��	�p}#�&��ag� C�IDs������{�����
#�r=b��\�Ma�/�䮆� ����P�����G䩻��P[��M�
��_�!��@#��I�@Z?� 2��j�  %���f�%��eah�OL�(�TF�Z���8�"ݏ��4�/�eL��U�B��Y�`�k.Z�+�	~�E���y$�	���L.�`&2���o��8M��S~���[��?=�<�s��׮N���2`����y���)
V�*,�p�P,yhxc�֣w�KZ��{��7�R�`G"�T��47!��>5z{�,2'�� .��%-#@��m�aQ�{ -�

e�R����W:o�!=�gƎг���Nl��+ʺ���J��Gd@	�=�Y���^�5�u
?��+�H�+�*���݋�F�u�3�l�a��s���d�C	�%u�$��!���MҺ���V�MZ��_4�vPH7���m8���d,ds��:���iTh�n�3HG=ȥ��!P�LU��n:X�i��,��|J���d�����K��/�����&��+��߫5�>��'f��	�F[0.�� m&�`�bo�4�\����7���`��	;Q�ˆF���1���-[Zrq8ՠ^SD�G��F�-/A.��=�B��晬HǍ�X;����݅�ݍ���H��THdp��)"
5����?��O�[1�}"�������o>��a2�?��\7t��i�A�ٲ?z�1�d�Y.(�Q�a����^�>���udL!A���:2�_�5��H������{�UL��c����GIKq�i�y�ǒ�,�b��ч!l��b�?K3��?��$�=������'�G<D�P��c��e>O����o�'`���i������[�O�E�sw���𼲑�����o��<���@C����3�����W�A��ˇl���-���3}<~����p{&=�:��9r-ÊN��ҫY����v4�Pֆ E�����������>>����Z�J�hiʪ�F#MK#��Y��H2��$�sU�-�k�UVw@9M�AyL��oJ�47�X`�^x���𸮢�Em&ү��>f��IӺ���8'4"'�q�pOKM���v���G�_g2��~��֙��b0RW� ���`���5hm�s�ّ��.�C�:^��c�����׾��>L�[A 	�$N�uAܾ���3��@����ǻW�����ԛf����ʪy������pFA��6�f�"���(�/
B��H)ܘ�]#�!!��,�>�	�##r
�QI뀒���B��ɔ��Z��E9 Y�(<l�$L׺]�%��WL2���6�UD�'_�l�14��{�<
�J(�
�
�p�|	���U_�#�#'�r��a�?��V�L�$��|�]z>�t�ᶳ�H�q�DQ�T��N�*-���́5�Db�h�d����!�������v�F"1�T҄�ʾ�LGI
��7UnE���9Ý�u�w�&���jM�W���J'���0&�w[�s�?l?�e��gPQ���4���"��BFz�[v���ra"/���=�;!�� fN�,�#Zj�Ƣ���6�w�m}�َbFe���|�t2߻���a�97��SD��6r��������@��H������Ggt{$���pP~w�j;QTf����a��{JS��5��]�r˭S%����
4�H����n��0C�-/�L�t0y`�ɖF�	��m�/�P>�>����T��"�8���+m0�!�-�@Y�1�|.c��&�5u>�y�j���Y!A�(.�IXBc�(Jq+����ʸ�=���c��3�z������%���nW*�9�n����N6�>F���.��k~�pxRX$c]����)�%]����#B�ʁ꾒�x�f�B��zV����*�j�y��0!5;�}P�b#���X,ų���JQ@K̚I��;� @xa��&N:g`Sg�z1f����>9���w����i�zj��X�{���N5�DfCH�㦹�X�*�����1���_'bÌ���b����әVq��zD�U�!Tg��B�?^&}6�]0�A�.�����Z��-L�ښ�	
]e�啍�������ا1T������$t=��4���!Ke�I��F��͖L���m��՛���h�bT�3=�U�TQ��� ���m���Ǌ��)4�y���pI�Ԉ���uh����6��w�:5v��Ue��=Sި� #tSN�\C�Bv2���3��ZT��L� phW@��6!�S�!y����WW6Vϧ�^�B�nP�lXM��4h��Z'h���i���ӷ�j1|0Y0��K
	㥽O	a�� �+��#� ʞT*j��Q�;2Qa��P�(�, ���C�5T{~���'�Kb� Ln;�d�������Ð~�K��O�4��-oh'��6f� |�V��y]	�X�� ��U�$!���`�5;��q^p��Vj��r�7��L5�!�y�;oJ ��ZA�{(���2��/ܦ`#�B������QU�v��<����eԜ�7����FV+���T�5d�h4�hJm�q$A�(������^j�0a��*-� tr06GMYȓ��%��2�(�Ve��o���'Z�޾=Y�x�0M�Op�XjK���dۚ"˕O�D3AY��!K(��q�i��|���°��BU���L�Y �)Un����sܩS���h�1��>Y���QF|�<�F���\d��ʸ�*8�"&4��L�f�P�8W�� �Kn���>P�c�qc��4
uʦԹa��xvmN�O~��U�䮥I�;��ɇt��'�i�<4h6>�]̔Ӝ.ڀG�y����>�z}��Q9e%��3z��]�ٱ����Z��Ɨݙ���؋9D��t��3�RJW���R�O[���>���𳿐�D�?D�E�ke�.:�PՁ�uA���k��6�/��)G �Q�b���j���W�Ĵ?0��GŃR�_���Vp#J�[�~�a�1�T;��,���3�9�32�J�z��5�26�ܞ��{_���g`@ȘU/�;�#�u�o�R ��RBSK��� ��Y',N&��L>Е�ƌ	@�քk�U���)W��֫��#��h��ߜ�?;qO�կ�Pa_�O�yط�eG[^I.���"S ��j�M#3�es&w��+�	�i��?���Ӓ��nc$�A��gv���-��&RȪ����W&�L���?!�Ĺ�5�^��gL%K�{8e&�9n���a6��f�l
3��I|�MІ��-��%��մ�Ā[�����6S����l�y���G��:ۿ�Ḯ�F��jbT{ɷ�^�c'{4UV�H�6��p�^MG��y���/atz oVF��N*3�;���8N_�(/���[���1�Z65�7`��=�yw,�R6[e]��h�o��V�`�M�7=Gw����L�똡㑆�l����"	�R��Q�T���N�i�v�w�:��}.�"��U���Ɵ#c�0�"�|��������Ֆ�-��]��b�O#��p�W�N{M�ԉ<(7V�^�K<���J��Z+��ã/�	^`05<�"�P�Gu$�j'����=4��b��n�3ʟ��#yŝ��6�^�7��Nы�Y���߁%�ԫ�'܃(�/M!?�R5��h�ﯙc���f�ƏyAW��KQ��yR�pѻ��W���x*'Ub0��ŷ�h�t����%���Z;���	�+��\�UGE˴!DL\M�4̫[�O?]�h��F.gOޏ Mk�	~�u4s8I�G[!y����������,��u�q��~���n�s��gJy�MÄ�>�U�x��8G�߯��h+U�a�S���N=dXM�N�o` �Vh0�NJ�������z�f2o����ԛ��-�㜆�Eu��g3x�|	-O�η�4�Vr�Zo�n�;�Q]M��e�
n�Q�E�e$��c�?�.��/�7QQ��Ađ�O�$���#!�~����`�x���&�p�Åk��cd� �$0���P���(�l��^�!�5=�2��z9�5Y��<�qq��ϡ��Ѕ�$9Oy�㹂K��]��-��D�ߎ��Q�V�/�X����	�	f�S���e�R��\�6������(~��g���s�����Qfozk-7wxUn�K�F_��}n�#�
�7F
z��}��9��zD�8��lga)��-κ��6B?-�+fb�g	X[Ը��i��e2@�2�|06�ɸ�ϊ�����ģ�0�?���}ͼJ[j�A%���jJx�A�Ps#{��l�b���i�A����43�H?:�*��?QW��470B��IL[U��mW��^&	}$���&�!�Tz��qr�q���L0�#��0�vI/�1Me��{�E	k5����(�I�V�x"�d���,��W:�R���/���jL(��/$�@Pﳾ�on�HdB�%,1D.7de�	���+w�y��)�X����dq�x����s����SFEbz�Ҳ2��8�Ќ�N�������*�J�+0d�B'u���]�ܕ5r��t�`/�x.�����y즩]�z�u���5�~-�U36�"�۹�Pג��Y�)���7g(kmu��aM�-��	i�7���'���Ք���X���>VcP�Н�[w�-Y�t���Ȑ��I����jk��ill�r�}�cn3m���=��7x�Eoǁ�N�4�Y�O^�+�I��0C��mM0~�1
�R/�E��J��ƋL�l�~&�����r׫F���[KW��+؆6�W�����Zî��8|K�����4����e̕����V&'�^@P�s��B���@ŧ�?%�:�q����L�ZHC�VK��:�^��+#��g'��ן�SDM�sq���c<b�o��H?��Db�i}��Y��9St(U�,{�-*m�c��&6�$�֦-�|���{"+���ʹ����,�q@�7H����u6N�5H����W/U��/�a��s� ��7V�Ƕ���ɢ�쏾�P��1-��(�q6˰5K8���JaZ��Eew�hn�uǻ�, �Sy��.��\�OJn
F����azK+�.�o��Җ:� W1�ߵq��|�I$���;�l�h>[� _�X�`�(�`��1!�>𙱾������ڛۧo
?�z�����	w�O�r1@�a���FL54U������T"�j��u�M>��<�%N��"P��Ò�h�Zƞ�ı�
T�����U��]=Z�&1��Q��i{S')*p��$I�(t+�W�94�/��P�ˑ
mC�3��JI�������{��21Q q4AM�����28��P�
�r��>������$�
`S��Y]���ʒS��<ē^�#����5�[�s���8aFB�:��x�+�>5�A8����h���#h�7�Wզ�D�5#�����y�:�6�Gc��N�@��A��\�e��8z��y���\;1I�u9(#�=��w=8&.��jb���T7�#h�����?`��w�()_�YN��_��
L�9o�r�� ���@�b��="���yԆ��B�Q�6/?�bW����6�k�ݑ1|����`��־��Y����~:��qn�Z��rm�^m�|�DZ>	�Y�3�cȀ�X�!N�_6{�)	"d`���������uN%�1nZ��`�����<Z��[�x��7������$��7,'c)�� f��4(��t�NxA�b�#������i�����.۰�UDD2^��͇��UXdS��#���r��e���ө����J�Ŋ�F(�=������ 2p�b-�-����x�P��W-#ow��'�w?%G�L�W�HAiO�?=mX��\��O��罏��r^�F?/\1�O����%=��$���Jհ�%���-'T�ީ�1�c�_����tr��p_�M��,zH
t2%�b�p̊����~�S/>�^����H�%�֯���O	��&i���1��d�vf9Sw�dC��/�J�糔� �~�\�̊Lh���5k�K����-2�#z������b=����ýK{<nt�]L����j)��+OQ�3�^سH���,?k�[.j��B-'9! n�AO�Z�0�e�xӥK�挆�Lv�voe=ag灑�e����h��C�*+�R�8,�����ˏA�yS�}��ze���q�O��ߟ?dU��j�{1ϾDT��X_W��>A�Tjw�z�!�6s��,f1���G����
f'��+��.�Fe��a�ܩ'6f�S��=pK��T���
Z%��oG�����������o6����N�v<6�v�h�I�I�B@� ����j���f�;\k�-���PIi!a3��e씿5iN�p����AC�?�g+Eq����=T�=p�!1�o��2aȟ���C�/|�ǒ��?�?W'��9x���TG�!���3�i�w"೺W�[���VG|<�Ld^'w!�uk�@X�]р\�V�bI�UC(��d$��d�@���й�l
L��њ-^՘9v����m�3wWY<$X�������|E�_�e��zX�F=ڎ�Пv�v�L��>Hx�v�`�$�c�G��OQ^�X��o��_��~�� �*c��g����9��"�b߇����
���&l`	JC������H�c�z���Q��dde/v���ռ�(�=P�D�����al,ZbZc�/���p, 5�����0�:���pj+0�~\(����}m�tv��E�!q����rIcjw(���6U�ѹ��/���^Q��j�ݭ�\��I��3�I�F�����
>�+��@��_��w,��.�!��˖e!�ٷDZ�[Ŏ���/p���$k��P!>��,�횏�1�[Z����P���%���v�v@���w��O��q!]f�񝙷;�m耗!�	%��g�V�P٣Ӏ��m�֖���M�L���v�>��D��;/��u&q��!������>��Ї�;��ے��;p�~�e��c0$<[f,�R��@l�j{M�j�����(�P���Z߽�B�U�ꅂJ@J	k����Dl�0���QFJ����Wa�:q:\�)�b$��|�Z}�y[��-�1���n�����s?��)�k�^��Zk(��>^	>��vsNϽ ����k�]�����W"�C�!����^���O��Y�
Bdvo/�$&��o���� ll�rE쪂4�U e�(`B�9�>��/e'B		��Cd�V�Ռ��0F�\w�g9}�TO�����:7ve+�6B��A[�a���*47o�/��d�}�
�e�Z�{(h,�5��Ueҳf��k���[��6c0m�̛a����;���c�~�[��y�?�)3EpLDeu�/ɪ��@�@U�A�#F��21!��׮���=Z�J@g!�>�ʭwѡ�ʕ��#���s��^ ۮ�LL��Ξ�Aq�p��$@k� Qn�+ɠ3�~�C�_��AA�P#���_�trZ &�`�8д�����
�G��3��钬>����y���s��*Ӻn.�B��������A����\���q�L��2r=��1a��1�����$a�3�����%	ߡ�)��O�Bo���C�Z�j�%q/,f(�`��u"`S������mkN���K��@�����]���aU71�C�pZƤ����qujhe"��R��G8�퇏�'V����Gؼ"A�c��>���8k��s��KAm���k;e��Xq���}�� #��¶ߒ?K/��7�<~X��=tmMC,J,�W# W7�"m��G;���g��d��w�^��=#�q���� �A��M^����lMIǃ	��1�]L�U|h�����D���P �B�k��k�9;����⎔�TA�c�pĸ��o?�2s�]�p��S��X�I���((���g��q�q�i�,/pA�KK�(��o:��/ S��+��LcHv�NM�{O�3D���ki*�$P���:�o�������_�6�1nӝ�?&�o[f�O�>`&5�v����� �Y��e���L�x�����d\���v�pM���,���)��(b�p�>y��C� �d}�f\��_CK���#�S�ʖ��h�h+Vy����Ob�J�a&/>sz0'���?7	�%�#4���_̈́���+��|��"=�k�Bd��~���U��s��,�+��,���h��:^��e׊<Q�O[�wy��'l����χ�=؎��n��O�߸���1����_y� �$��CT@�g�ݩP��-�n��y̅�!�:�+o��x�E�X���i�C�Ӣ?�n{�~�����Ī��h�*���Z�����B�y����A�d�FI8�N��Q�H��𮷘sBpn���	C;�%�k}699�*,���!��v{c�,k
 �>d�q�TBi��8ĕz�]��L�)���k7�؀�!o�w�d��a������_��ZO�Rg%K�������U�!������F��5IwL���f���UKz^�M�a��p%uIPT�ʓ�N*�?o	��/AE�v�L�Z,���7��%kj�%�J0��G�3�SK�`������2��l=��ܛ|�c0���YK��Ap�D��jW�1T_t)��*�H@��AT���Ę�:� �PN��ة��ƙ��#op]��~칾с!䱇���7�l�_����H<d�׸?Kx��i�$�w���.����gU���5�B�|D�o�o��r@�v	W<�X�\ԋ"��:O�y��ò�̆����Y��c�Tm�r�t��v�a>V����ʀ�P��K�e;!��ޫ���,e� ���|>�2�����/ҐA}�fza")d� ������=zpcuQ-;�3�X
O�����,�ݕ��jᬟ3�	�@	�I�(�d�P��P(R�y �zY�`���#(��ǟeA'eF�#��q�r�&�B�ȑ
��YQ�XА�,f7=%��QU(f�KF�ęYj�w�2֝"y�]����|4�$7�\׎�O���	�^%��}���%�SR�QdW��s�4���_��sg�<)��V�ᬉH�3����u�d�5C�<+��{s�D��S*k?�>�tL�ç0�3�tCW\�j4��"0�����~`���a.,[d��//����^ee[���;�9D�&��96=2��GN����:x�qVH�u~�tB^����#�NF]zthF{_��{J՗H���zT��aޢRt�]���ʃ���mh2걳Y����dr>����y�����v�3���s�h���Lt3��O����r|��R=��e���9�� 1�SL_�|��#�1�33��[��c�q�^�B}��Y�����*�����?
�hr��9���7��:k}@�ae��*���`g*?���r�����:gFP�)�u;! �p]d_�P��r�G�v�-�hKM�Н2pa{"�:M�Y���,�,+��_e��q!�x�U�1΀ +'���x���8�����q|��ro�o��gczc신�la ��@P��~U����L�k��'ֽ���� J�����|�#!��ˆ��Y�h�ڤg�b gX�L�v�s%-��jx=�|��a�fu1�9?�^�fo����Щ,ܼ�M�tX��@=$��/G5��t���8�T�NM#���k��@+��09O��7C�<��8͢����*�b�G@�6Ւ_$����3<+����+fI7��6�)��#>Պ�?5��m*��{y���������z�Y��G�"0��N�y�0M�?ƍ��R#C#(�x�Mʳ�M� [B$4���03K$��H��k�*h*�8'�MT�G���5U~���R,����Ѩ-�I��ѓJB�uJ`��+�!�-��`��De7��'ʸ ���BFofډt�K����o�ɡݽ{e�^�ou_UC��^.ߨ�ty�O�E&t0s(�M����7U�����b�D�{�c�W��2��Y���Ab�&��ƪ^��p8�z��n:@x1���j|R���m��`v�����0�lݯ�%�S􃅕����gN�`�v1,@O�h~����wb.G��߬�<(>��i�cv �9�'�8�e{��8�Uhv6Y]�ܥ�B�˩��3ZR��8���VV����ˢ/��0��wN��$u��o�4Pچ���讽�&����'�-TUp�2'�l�G��W�1Y49s]��{.u�gC����o{���&�+͒�ܾ�§����w"�����٣��`��]�?Hy�`L�[&N�Dm&��z��W��P�գT^Y�N56"��F�q��B�(��yI }�O��-i7nj��E���M�D2�M8��&���v��O�60b����.x��Y
��Q��wSk����5q9(�nw?���;��VE�U�2�C�;��{f�r*��6�W���u]v�Ơ]���fB�<[��l#��/��$�r?��uѶ1���~(}���u@��/�A�˴&���~��׻��%�5�4��;��ɠ��I��7��$��Ͽ8Lo�H�8X��,�d����r��/P\�p���>���$?��Ňt�J_����@d���cX��i6[��p�.I�`���y9�~�3/啎񄞧����� �r=s)������u���]u_���$>�v���M(�u�>���A���Ef?��7��a_:��l�7v��OAQ���^X�~6ΆD��z�v�b��	������]ob���.x�7b����gY����	��2~TE��G����y�JQ]/��?$ބ湦@E���b�/e.���V�[gR[��.��{�
)t�l�w�'�K����p�/��c���c{,,j�=��MIzzj��^p34�K`
~���	�O|d;�I���~��*\�@���j�C�=��Mm��N���N|4���g`P	��� �*��P��T��~9����k��F�=�9� �ՃE�>�9�r�]0�VV���Ļp&L��ʖ��欵�{#���<��(��R�{t�Q(e�;]�����Ѣ��j�����K!5�R��)���Kح��Qy /���c��s��/�!�+?��䫐���3_��(qrwxO������m���*'�����$D-�\��ۆ����t!���a{�>鮻�<�c�،9ч#c�#��HI���.,�m^�W�mz�?RO�>3N�n�FoH��MPns��A���Ĥ>¿�Z�&��K)v*��������G��V1��;w����UU��oz�(Lj�c���V��5,Du��� �r%�K�n��'�������u��g � ����0c�?�'h�Q�x�n N�M+3���)���1D�l��2�^4Z��S��( �x��k~3"$)s�N�H
N���Sa¦����vW���ؗ��
J|��J��'�nS"�#6iC���.�jયU~Qg<���`��)|��h�QP�gr��~b��J����f;/t�ԟT��J�˭pS�*� ��g��Ƕ�,AR��[��]��5H�t��������R��h�n�rA)�_7"����
�{�
�j?}D?�k��R�˦���7�����o���5�J�b�Р�SMC��`�ƾ��WSO8��;p�"g~�g ʏhJ|��7�7c��=}�~L(�Y�^�2�~7i6��{�-3��y
Fn5E��:�)(4;��rk�Ѫ�F,���J���Ji`ad���Զ��}ں��%}�Ί�w%Ɵ��7)��S�L-w"؅#��,z�u����?��m[T�"���P�7�25��v��AJ��Dck�WǦ���g]�!���G�y}� ���zi�0o�'�rz��,�
��<�*\jC����&"�eCg����~��b���1��ƴ���8�[;��Ц'�}M���3�H}ou9@�w��C���@��^��xn���w��*�G\e�A��s*�VRʮ����m�� +�'<�t�js�%o]��	�ϙ�u���]��T%c<Crz7,��=��ȡg\e�������f_��h�Ǡ �)�\D_�*�JA��k��g�+E W�ӗ"0������.0@�}#�̭(��D��1�
����*�?�z)n-S���e�h�c0]�4rɜ��.Cv�� �B`��	����Yo'e��7�}d�{=�[�>?Q�L��#/��h�^<��|�ܸ7����fy/�Yb��L�B66�U���w�,K���ǻ���
ji�4�mɘ�W��R=g�u��2���M1�)(�4���4������[U��|�޸Q����^_���(A�?�O�϶�v{,_"�ι�!���D�L�x�Aas���UA���`'[(^D�A���T4@�v��N��'�ލ�õ}k���en�@��E�tV%�L����,3z��?�0q���b~��W�c��YX���v��ب*�/�Ӑ��+:y��tg3� B�O=-�#�hR����) ̜�t��9a,$�ɸ�0�����6��o��v���ݽ��M�fy�:��1�����B��b����9� u98���s+�v�|���,��cؖ�eQZ=v��2+��
&���a��!m�POi4V����"� Ӡ�(��i�+�r�<�N�,o���sD2�����'��T��{��.��u�$�☍D�1O�ص��ر����&��O\Nx���+<���[y���)���K){�����1���l��<������u��J;��x�I����|V���s<���.Iq�Y}];��Be�Z���v�C}r�W6�2[@�fS��=�=�b�1��RS~6c��o${��z�ປI-��j�__� ��4��1ܝ�B�g&�~��?�M;M�)DQ���N�)#���We��充�Z��Z7C�t)ry����j����|�Fh���,�q��v
a������{O�s�*_�+��o��(�?�`-�5]�@�$e��|�k���<�Hu+Ӈ��\,sSa�`~\��M���c'���4�F��)�$J���:����}�����@� 	����Vn�̔3��LĬ�ݱ�0��u��O��(@�W�
]�Cv2�����Æ�Ɔ	��|`a���ܡ��7{Uh5��-"�w>���l4�Ԁ��j�E�g��Q.��\��C&�<k�Ψ�؏�΍\�v`���c�����7��I�
�l<S��V���5ӡFS<<{hzn��� ���c��y 3�inD�dp��qH�4�ApBN�U������+tT�Ct�s�0�<��²�!",�i�V�X���HDhp@�H�X��,q����
����� zs�$���S�/^Z�����L�M���./��!��3yJ��=�j:V���@`�1i
����B�Z�����hm8�&q;`lz��+\�><��~G��H��p6��U"����Z{��΄���u���4g@�wi��v
�*	��$��.�������{�L���몈�n�̵�i�:HZ�q*����;�E���״�l�[����dHj<�,�?ֽ�x�;�1}"G���� 	q�d��)�.�5!�t�u���0}�����v�^X�i9@�?���D#W�h�)2Hv�j�D$�O�0���,���c�<6֠�����D��.V�Ƭ	��BE\����Kk�!
�j���tk�?f����^�N�3���^-�]�-����-C��9?�8�X-O=a5�	f�v$�������6� dy_T�B���&<V�� )ۯ�1:����@. ]K�孨1n���t����\������֎��� �m���8�b��5R��x�x?��)��g�ؤ��W��,���e��F�pN�}0�F-���������<7�M<DpڗD��vK̣%>l�U��B��L[�{��X�:�_s�,�P�:�ab[t{$s��Tޛ1��Ѣxs~!�b�0������� %o>����5���њ���۵�� ���>l�I#+ltG�s>a�H�No=i?z�����-�{(.߼�Qӎu����"�����@zҟ�a���*1��\������#c{9�����C��n�����0�h��S�"��L��{/�1V��}9[l����#L|�����Ezm^��p�lK1S��*����w�8CmtM�-s�ժxz <z���2�r�|(���Iy��Y�d�/��D��(��ݤ�@j�<f��Itے�Ծ�G��
d*tϔ�Dз�'��g�J�w�52��8}�p=� �˲2�	��%@tߧ�?;�9�3��5ܩ߲= ��\?��';���X2�[�sc	��V9`��"������n�Fx��K��,k<��
��^2L#����G�R��+z;4i���(>p4�=p/ׁ^���n�\6/Y`��b��b�����C�o���������{�6�	�ZZ�|!0��d"�t����7��-�*F]�$�Ҏ�QVv��Hif��l��^��uM��MN��ǿ@�'K��f�~��a��$!*j�EU(c�҅�b�}�a��R�Q~T�sF�y��K6T]��ա�Oll�V&x�ilZ[�Q�@�Ͳ����c�d�f��j�L���zLk���f��!��%{c���&+�V' X�@]��\)�c?���G���/�3������O��9[�ю�}�&,���9��S��*#CF���**��iz�BէYX��d{`����pN��NZB���=�`2�z瀃�'ά���88J1�w�a[�q�z;�nmw�l�K�?�pc x�{B,���m��	)�;*��?���[��A/��/d�>�%����"p��\�O���G�C<$90��:��b��ly,܉� �aU��>e�;���܅9\�eMx"tl��x*��#4?4u���k_������o5���J����t�\:xq&퓌Pܧ"���1d,���D3�H�n�u2���k[n�̘*��<|}���#�"��c��i�\zd*�����+�+o���� �N���3��\BjR�D^�����jHz֩�+���~d�����!��,Y�q����� /,!�-�X�p��ڦ����9�~k��z*w4�ƹ�?p[�2eE1���t���"��S������)C� .�|��E�(rb��s�����!B&��`䏫[/㣍�l����]W�	b�U�-%G���Ƌ/�x{'�PS���Iz���?�Bupa� �`��ƭdVݚy�r���h7�A�Y�0��G�w%*댍��m,�}f¯��~�D���h�W�MY��s�^\c�0��/�PUюV|�h��� t��|���@�j���W(����������
$�k2�/>"͟ V#v���k<��N8����e���Ϩ|��$U�}jM/�#G[�&�Rڭ���� ��$�c�ő�<"����CN����ηF�:(�x�	1�)U�V:��Ț�c)��B�m����:���������e�OY�V<��
n��o�V�W�eA��oH�T��1�ă�q����a�d�h���æR���pfq_̗�Tڔ��m��;g�z��!��f��ur ��n��ġLi-V�ֻ�T)O��1>�#`�;���M����鉬m�����'&�Y��S0�o��$X��qD:�>��* ��8g*�H���^����ޫj���~�l9�(m�G�XM�F��"�T!���"K�W�ߵɇ�	��m��G��A,�G����[�dl*]R]%�7�����^e����<s�f�{�����]����@`�J�LX$d���d����|v2�L�?�����\�
�-B��lb)�2����[�D�!�@:��t,�I�ҁ �@J�����{����zn���ʁvJJ&e���u\}���*�?�P�V/Aպ�|�v����;7�u�3V#M�����I�Y���)����J����=��կ�����Ѷ��HP�%�p��J�尃��/ͻ�tԲ�1�IC�����$ ��4GmB?��+��N���T�m����#�y�?ܞt&�#�п�� �A���\f&
�ʡ��b�߮�D3|�*6!��Z�[�7i2CDb�sh����q�����N��P�T�d�Eޕ�r��o��G2KӠ \>���Hvi`sN!��,Zw=ڡ�_�̹ҍ��}�U�G�� �e�}���>M����l~r68�t���H�*蛘�vy����گ>Hx�2�ŗ�Ar[��.���|K%�y�-��"�S�7��,���V��K��B���nY9&��8�mB|.fv�9�D]�����v\N�!����y�6�p���Ď���� �D�}F���z��Zf�	P�O��U���B�a�[ ��+�����T���HVK��MA?���8\>�`��L"D��W'�<���S )b��s�yf���}%tq���$��5
���?��Ё3�q�${�M�k����l���*��Z�Z ��Cv���6a���ܘ}�ϵ�)����͒�Y��Aae/�4�qB:f�%�q�^��}�g:������ ��4[�W��T�DF�0be��$�&qQ&�1BMD&��R�h ډ���Xϝ�ZZl�ۭ��Ñ4��_x�Mc�`tL�
�a5¼�͇���zx�wu�2�'W�'"�?z��ߤbl�a>�dx,vV0F����Z//v[>N�;W8!ȑ��W@G.K�k)�FM����O�!���o�m+>ҁ'���О^��Vd֌�Җ"q�h�G>��z��=��	�G��tò��>���"�b�0Q菂AI�@7PR�!kWOů�!�%� ���rE��g��9����v
�{=F��'���>-9�Cx�ϻ�RB��3��J?g;- �����z�S��>��ÉT�Y�qOk
���Х���Y�'��0y��:���{oi��*3��90��:hE_��c@��ƞA�nS��qn:KG�4%�{ʃ�8��9'�s�\��V�Ko�6���[7d2��;�C;�>b/t@�ȼJ����Bk�!�'��U�r-F���W�%�Zs��Y�Dv���w1�e�xF!(q���e���P�������wt����61~�O<6�9K ��$�<J���)���ʙ�-�`�_-�?g:�#�[I��� �0a��8/��,���~"P��F2y<���	d��Qɂ��~la܈�]��>�ъ���>&?��5��8�4��5M��>B5b@Q��f���lGg8콗��m��d@��$������I(l��'���Pƚ.��L��w�P���]����J=&{n�}�8���I{�
�y���i�-�Ř��vw�lC�����1�"T�n�?�뎯xm紙�#��>O�� ��2���}��{�-u�
�m]2o��0�����1bȧC5:čXg�o��`���o���[���x�.k{������Ϳ�+D���(�|���zѫ��Y��R(�qX�8���K��Ğ�A��+�B���,�=�mgq����X���SF�; �Ӡ_�+ :B���2�y���،������GsCy��������_�S���r��}2�h/�/�Ъ�G�ދ��g�v[^�t:؎9H(����\Rw6�VG51;]RwOT�?�\��k}�׵Ģ�Mu9�w��O��>ȥ]P9����u8^g�'"��~��z�(�>8�>ak��Y�U���C��V�{�뱚�di�/c\�m*��]!@ls:�fZW��
	k�F�@�Ni���`A�c���{�5�����)3;dz�2��a�+2d�g�S�Dv3�,� �!P��܇�_rȳ�-,��8��b�ĉ{���(�.J��H5c v��"�b����@�k���+*��߰���s�%�<
Y��Q��wC�Ƚ<�rx��t6��~�"=�IL�zy^Jp��s��u%�" ��&����*jNS�O�ݻg>��Pذ�:�[=�Scd�B����;�z��ti��gz-IK�#꟏��2��Uf����� �z�4�}2��T_{/��\�G1��i�N���-/f5�=w���@1n^���F/�n�bF-8y�=��&���_�Y�|�3�1��oT�O���m��D��L�6߬\�ӌ2�������&IoM��Pv��|n/���F��W�{�%���$)/���¯��;�P/r���?��,�g\�T��V6�T��Cp&ݖ��g��?�M	_8�����x�
_`1��v��]�X)Ӄ�>b7���n���8Wb0�w��i�B��W6X]'a��`̏��E[-�T�Y��p�8�|LL!������Hr��Q��
���r��l`d�����'��ѻ���!�:��F��A�X��c�g����朮弍�I|���ٙ��D�ho������vB0S��&3h��,��s�����frp�2�F e�ƪ�����K���̮�V���۔:C c��B���2��d�{�[6��D�z��l�Xvd:g��p���s�=��HV�8�n�.�c�����2�LwBҳ�kt	_":�"�����.���5㠦���D�z��s�1A�t{aƳ���4i]���ӃY!_�QqD�y�\��.Á����5��U��h����LT	��9����~K�bzViS��A��F���K���f4�c���JTRh���G�m4���R���..x����(<��B<��!��}I��4��bcX'q��ӝ�����
A�5���	t`�kʑ�W��L�����|%5B*��P�����]�}R�`�*MfSVm��Gv[;�pw~�Ӊ�����@�/�"b<3�x��yu�NņK��]�4EM�KE��X��~���Q�5Fe_��l����0b-q���2юzvP��?~�t*�h�&�%Of+S#lVK�&�*:�
�n�j�t�����L�G�I�D�/7�m5u�w��7u�(�5l��W�b��$��&�Ec�C��`����vµ |����>sT9:�߇L�C��$%�5�==�4$r���3�>g�f.�Zx���,��^����KߎV��p�ު` ���x�g%6����2X�_����1vf��5� û��C0�!��U����dޚϑf���,Q,�3�d��$Nm%Ec4��_��(^�)�f��p>���\$�U�TC������}��в�"V��~,��8R�E���rF�|�.����a�&���zqJ�.�B���&�%z�us�uh�:ͩ�fO]���_�;dA{q�6%^c����C��z��}�p�G��^b��)�^[/"8��wg�H��Ύ���-�6_â�D��%4A�ܶ�F.��LL��y�ܶ��z�R����*0�O�4��/�(<�}�cك>��7���FY���t4��p��ɥ����ʻZ?L@oX��\Qa[�"l�u/�H"�7Ja�2���M�ޝ�.cid>Q݇sa;38u�G?L�Mc�U���c�Vp��Cm���Vp�����F"y�}�*�
Oxyu�F)k� 7�QMu6�jQ&�m���Y�^"�>������0㢊Z<WI3 ŅXoݦ	�8N���^�^
f���h���<�::�ĳR�>u�j�y���|�.�dL���D��̈́&��P�
����V<�.ŋ�;��n�6��=!�R�ØE�^�4ZKS*�Jd�3Ԗ�{��];�MLL��%��x��AMs�Nx���јƺ�]X��a(��Q�N�u��m6��W�յCA!�eؿI�����K�(��ǟ�d.�5�O�ļ��{��Ȝ��?w�z�\�G��u\�,�?A��d�w�B�,�ESɛ)���q�5�w�i�ύ�?� E|/��WJ	N��*`�m�bRZW�F"Ĉ=�n� .�K�sMǉ�$>��$ ��N�*�m���Z��T�x\o�n�'�#4g�0��D�i?H���:�� \�����֏�l�Z��/2����y�9��).�?S&�n�*ߦX��:�C:(�$LQ���+?)��)�2rf7[�Š]��KYf�j��,�9}r�c ]�k�ʭTN��K�UbP�jWS��,x�v�7� g"]U/���#PErDY�j��{<�&=�"�?_�+x'�B�	��\�����&k�&T��-� dZ�-�XL���������MJ�Co��D`Y�۔��	���8���p�λ�ˬ֚�1���E�
w�ě�mn|C�bH����/~�t�����-�ӝFR>�yH��)knu0 ���?Pu.g�~�XA[w�$.g�"�IG��L���
��o]	"Ҷ3王��ˠ��陽�#�xC����v�G+L����7�h<�<�h&�lcqǻ�r���tL�$�X�_q�\s��h����j���f
^��+���F�&�Mצ��;���ys�� J�7t>��R�D͓���<ζ��̣o�Lj�6������'�Ux��4W�h��#qꠈ��AS��nY���FV ��v�V'2��Ɣ���+V%!�b ��E���@�LT��!o'^+�Bǥ�,n)X�'Z|֝�,�͸����{l�ı��6$N:ʿ�!R��6���MN��ޅ�v�7���C��n�#D��On-���w�$�2�e����>��4��FWKF�
+WH�9%��_D}*����S�J�v�o�JA���7*����V���/��=�}oIUh��X�H%��e��V�>��6��ɻhw�[VE.#�Xb�T����̰��
�'��{�C#��r��͉'J�4�iB�ҝ�6@ǘ�`��d��i���x�7�#Z�NiIF�Mo1�d���vm���ߤ��m�*_�"�AtP�Ú��dW�kz�v	��AI'j*t�mD=A�
��<�^=��]�=�E�%���Y�O�A��bx�D��l���f�Z|J���r�!#�:�]��ޜ(�Fלe�/��n�5�M(-�ne������CM��P���� ���cr�فo�#���pk`�<m�Z):=��������;凫����)�iM�,U��a~+�>���Y����M՛�b�]@Y��t��ɹ�e�a�B0͊fa� �e��De��D�t��\퀣!C��b�6���H/Ȑ1"�ɔ�(u���s�#m����}'	��^��T�U�sH�v��� $����:
=s�۾	�����T��|hu��+�N��]�%8ˁ��:���49|�hZ����ѱq5�Z���ݭ[� ��:CDBӃA��AJc�ۈA���P�[��!�%B��QW�q�]��E�A�⃍ޔ�K���A��h����0	(�5��tlN<�Bh(�h*�1��f���l�1���?1���Sr�K�4��3�\�1w��6W��m����0zƬ��Q�j�;x��?��E�c^'�NЯ%�Q��	|u�SQ��t��P��5�a5?5I�3�� pP�S�ͭؖ����[��'2�p(
���'��7\�����j���q���؁;���	M��E�?rc��U,�|�"�16 �n�EJ@	���'�@����b}e�X�v��iV�~PLa�����R8;>2�c�v�����
(M��ы����Е�\�h��zP�e��u�t:���bQƃ$1сH�r�m�y����%�{��)Yy�g�u׃����Fn�f���k#x�F���듬0Gx�y���oH|w�7��Tiٿ��c�v���ͣ@�!il$� ����e�vNş�%]F�@����(a�	$0���8���xu\�b(�l�r����7�$�P���SJ瑉:�2�D6�5��˩M�i3��x�,�=�c�.�eq�u�V�,v5�J��ۥ�~��;{�T)�e0_=a���$1�H�]��/�XI�	?���z�R��ߴ��2�[�@��wn^�;p'n���:�a3��ʅ���G#Siؽ�p��?��(��D�}��f���Ϥ����(�Gc'�{>���a����`����/<�6�a7V,M�e�Z��Ȭ�+��"s��'�JoQ��L_��ZƷ�ow�
����[*��CۀrxLC].{��Z����H�4D�K�i,��t�.������0���k4=����^Eoa��w�����������@�]:+�nR�D6#��WȚo;���Gts@3?&��L����M��T|�Ū��~T�I�!�e�Y�مHf̨�8N���Î�I
��3�UVșv㚳��OU���|��Тpϥ������a"��+��|���B�a��hd84K:�~�������
Bm�Uz!65<F&�!����!�L�{RV�2}�W��M����UK-aݜ��|R�ǔ=���b�}�� 8Ҷ�4l�b���^7��j&i|�"F�㰛�R�+�#�	�I`f���~,��䗄V�f���W<�4��H����C���v�[J�Hgc���� ņ��O�hx\����B��<���C�|����;C��V��o��aC��WD�E����g�ʬ\c�ܤc��ؓ	����	+נ�B�+����-+繁�4����x�m=��~FÖ���@Z���ht��tί��KSȢ�33��l�1��R��ֹ��Ҋ"��C'8��*/Ku�����љ�i�����Y �R��Q�����2C���ýl�i��8��8E���)�M�&�[�,q��g�˩m��;\��SZ�,�,P�>��|B�H'��))Fko���s�㟗`����7��@~�k� ��Yi������^���T �Y[$��DDSIp��=�h�,ZQ���u|ʪ�=��!����8nP�U_/'g��y�w��v����n4Aq��KЖ�*���<&a�1��dc��������ь��'�6��SL�
��!��1��r2tq��HIw�Zt�p	�9��HPu�K�(�����W�E�b�8�_뷔��K:Pf| 8�׶��Xdd}k�)�HY�&�+�o �ehs��H�n��x��@�����c9�d�Ǳ��q"6~IDu�&��JX���2%����{2"V�;��!�+�b��p��%H4��I��h{�=1���Pt g�'*��dLb=
P�֐~l��ҷ�`��U�ҵ�'D4�N���u7"@ɇ�4��֏=&�ė��o�	<����
�s(��h_V�#��6)�*Rw��;�k�qۦ�"C��3�[S񪦒R�H�^tud"�}�zl,���d��(�[�$�V�?���
�ή�t�.3�d��7AX}�d�[�Պ2+��?ã2+�e�z'��ZZ�c�m�_��Q���h��	V�׌S�
����v9��h�@��e��U�KS)���]��ݰf�΃�9�|jf��D*M�
�VH\��J�7����o
�[+�1���-����9�3�g�H�Y8��?��08=�3��^�$�Ԉ�NK�8� <Q���7�df6��WT��Z�^b�{|N������Up�Ȼ�,�p�w���\.x����J�����G�0t���ygc?�wU��2��<���R��vk̹2Q��끸�o_�
�hƇ�g|��a�yX�ۖ���U#���j⦽����cc�2��I�J{���&(����2��=��-,�h���㞀����F�!�Ɉ�h�����LF�7�"V{�<��Dc�Σ�oq����r�$����z���
+Ŋ%����gL�ʋ�H67�)P�6,}���{뽳��Tz��҃�A}s��햱2)L�~��gj�"�ȟ���A�G������$��$�Bf��`?���:��k��h�Ѝ�<á� TR�ȳxJ�}��qo�}�!aÛ�
6ǵ�a����^9�9aU�r�eSw��2!�S�_jL���
綊U���@�*!��.�o�lj��vj!����4��z��%i3!-��j�]�tF�cW�;�}!��r�o=�C�/���&㚍I�Y�E����*�W%����3+�+�k�-���9mT��`:0g���+U�&�my��J7�_����{�~k��t�QN� ܺ�o���v~a���n�[]�{��_sQ~ �jĉ��D������IhD$.����a��Q�.�E_�r�x�0>�q�cJבq���m��^?� �RCd��	&f=}/��ר�M�$�y�vr�p��zR2��8�\1����U>F$���A�fN�{��d4���w����h�)W�8���y0����^ba��� D��}��G��������ʹ�" �P'j6�"���7@m㧮E���$�7�����ǁ��Ɍ�!�mh� _�daA@��O묉D�v��f�׭	t�E͗�?��7{>AН�*�\2��'�����ߎ�6�i�UX*��T%vn:̟B�ă��Q�O�a�(�t.Q�����>�3蟆¡e^戨��"O�1=���o�ȯ�
)��	���Z j-�J~�#v��r��t�<��2ȧ�����9ل��v^�������O��<M�~`�U� U+T�]
��e,u�a�����l �$����?�r`P�!�:��8��3�s�*.b��kG�B���-��
2��ac�w�M�ǫF������Zcۀ23�-cG��)�Ny�?�#A��H�~MQ���
��AɆ�[3�W���<�
��iK�i��5��%��'_}]��:f����]~��]��e��G��o��}�Wզ�07�p�ZJd�D]e�7��7�'(�vs�q-�J�Wbto�
���v��(�(�3��;g^����ģ��3�_�gI�\�GF@���/�PS�@���8|�-t�<jó�Ц��);A���@�xeÅ'�XO�����d*�zA~�"�%�!�:5�cT��WA|09dN4�G8�A8�;~�^�8H	C�V�A[$y�8�0�v/L:��䏥1=�w��5��>s<F�A��Ytm%�J�����G�W�A�m0�TP���1�ゕ�c���ܦm���ϻ�^�X
��f�i����$��E>6A����<�����Ӹ�0(c�o;���h[e��Ϙ�3���t��Y��;�M]�8a֗�*�WJ��!����>���<?5�1�;��.n��
�4�=�r�td�!+ݘaL��A��e"���G��l��%
�LM��.}�C��e��WzӐaI��w�H���߮�J���]4i��N3�Vし�y�Na�p�Q�G����e���������֚����_�h�+��)euoW���VĦE�Hs����]�ݣ�I῝�o}��6�ޅ��WQ�UK.+��ڡQ��W��vo���U�5��8+����XxOԷ��'݄A�+~�o�;�:� 	ԓJ��������=ϑe�P	�?�lZr�W���qG�֯��cF�\�1�~�/E���������k	`�)���9T��V��E��<��\�A?���R�1�d)08����.��.aZ�%��ī�a̲'���f蛖y�vٿ��������a���6:[���}ۯ��E -�f+��_��X�M� �)?j�[�\�na��:EJ��=+��%v�$e�4�kq�X!�٣s.#�0h��s�X�N��8����y����;V�t���غA!xG�\��5CO�w�C��:T�;�uDPu1ߔ�V�f�*��N�����d��>fF��� �Tw"�Tv�bOiه�N]�*yڟh���Q�.�:.3���!xz����Ua9��(-�>�5�]�B!'�b8&�!
X��%��e�Y�M�{��
�'o�3/�%!�����Z�
������Q�<.������3$A��6�����@����{0����,r�z�s�ֳ�1���N�d���!�=����S[�p��~j���L���&K��S��K����`S ��l±��u+��y��w 6���d��
� ��x=���c'�qB�cN5Š��9��>8zyc�'Z�r:�NI
����c������A��9�Y����
��:��dVPH$����yh-I貈�7��	�~ނ�}NYJ�'�_)Ï��B�<��*I��½�;�!���\Tu��|'�w���KM��H԰��EM=<�ӫ_?yWxwf)�b�)&��z����Uo�^O�N�Ă�����%�����Z�� �ݓ]��9~�Vn�N�s=}]���F�W�ͫ Bm{�6:Ԥ0	,�=W1e���Z����HMqjG�����+��tFu'�����ex��n��U ��ܝ1$��V��ƃ�ݰ�L��>O�´I�3�ښ�c�����"s��ȁ���%������<�\*�>/�Q�h.b�9犳�	'UA����1��{��*���D+~`4o�]������B���C{����q�|_M��H��r@}WvO��(k��}_�|�n�a�����Z9)��"�l��G@��B���߼��j��N�79<�l�(Nh�{��Z�\_�,pɷ����4���6��NZ�.�8�jöӫ5�N�Kq�N%���c�>�!$�68���k{[R�AN8�֢��ݯ;��l��tĹN_6c�b(��O:	E�(-����c̱p,y�ƿ�۔^�^5#�0D��_�Q�H���q�^l��1��ߧ�?�=�y�-�ne�ݳV�Q7_���q �ꘇ8pd}�^A��������^��ؑ
xP�I�0Cx	V���V�_4��6�~�b�|GX_���6���Bj��_m&���ۨ�����I�l���ԷW�k�wt���8t��8+3Y-�j1e�m���	#T.<3��8�N��H��$x
8�}��V���ꧼu�]�����n�b�M^�Z�z�[�z� r��*�24��T��n�FZ������$K��=�׹�=t���~z!��5���蓟�XV4?��w<T�?���"Κ(�N�ӖN��r)3�э��g��a�7��;ކ�6�R�\�*�`v�;<ePD�.�J�Ƈܦ���ʼ(y�~��%;���Fj��r#|�ο𘚏��\��šsAx�����vW�����z[+��M�x^V�I�6�'t��SR��G��W3$+�6�����m���D�D��`O��s�c��(U%�-:V�g;���Pu@�NKy6�C���י�8ݎ��hK��g���{#{�ߏ)�yBFJ/jS�z���WN��4�ڶ��<�e�����bb��w\�^��R���QU��[2��h�	�o?W��aw��Fd��}&�8\{h�׊���R�dp��&z�Ǥ@�,!1�=���F���=�-��Ar蒛�����L���L�����ݽ91 *���b7��꘍�ڈ�]Ybs�R���AOlr��t���^a�m���\���[XG޹���6��nK�����/�!�������>m`�F�ǋ�lA�����l�W��C�՞���׸ڀ���y��̀W�:*"�[��F��j����G��rJ��c���cB�~����
�3�?^�]�p�</�Y\=�,�m��rE�����o�rZ
F��@"�.A�8���f�����[�9���')���Z��Ym��.�3Γ�l��Є7!�����n�
_��Ћk0�J��]Qw�oQ{�?�ƍ����`��U�I>�Vj�}[CI�A~�<��I|xP�~���C�Au�Q�O�JlT�y�������\FR��7�X��$�A&��5�(�S��~��eu�Q)ψ�HSP����W��7#(ac� ݜ�՜�,H� ��T�� nKܣ/��-�M���U�O��^=i�Gd��r��V:����	�}FkWߝT;	A?r���C�-���4{+�Du,��h�r_,�������*����nbԘ�=�MZ(��:y
��IQ-D���� �@9�,�X7�}mPE��՘8w�+:�Z�U N�O�YӳH�mvs��Rv���>c5u8�}��^ys���GܓZOO%����>R�����0ٵ��<��ߤ�&վ��Sǉ��&H���G{�a��`���D���	4%E)E����DhPI��̏� �n�_	��ɲ9��̩����TIH�״�� �?����n�yg20,�<򻛌������9�,\���s�e��ۗ�&�N��,]7Bs�Ŕ�5ي�p}�aq9�1����_��w����V�V�0zm��>���������D�]]k�B'���S23�N�]��r�=�X{�:��j�C��	������a~#]��x��AS'˵���Y}� 6��'�X{�l׷<-�.A�{�ʭ���mp,"0��ݲ�?c/ó�Y��~-����'���d�X����z^�I���0)O�WR�CQZ���K��/6���{_t��` ^Q�Ɉ8�$����{�bн#mͭ)�î,|ģ�����3��j2���T�&I�W���KX���W���-�E6�l�<;D�7�M��a��F�=��ɎCb%�FG�L�=�#t��[4i���ףO�¯�]�h�}h�Y*bb�, �d6����C)?`q��_(U���u��������uś��Ȃf\���%����S'��Bf��ٳ�D�
�k�!��1�'��t6�� OHP�T�����50Q!����X�V.̎x��NϙhM{��O:��A-k^(���v��|�w�xT��~�Y�1��y�Z�)�q�ƙ:�fb�ű[l?�(W4Ot��H�@��5�;��,<Xԓ�h����&���UΏъ�|q����W��R|�U�0�ߖ��{ۀ�Z���4��m���t��F'Q�K�]�(Y�+?k��b����9bO�������~��:6h|Ni�t �I �S�^(�2�C.�߅��#�2wI�-X�9�ɢ=FY�4�.ߪXs��D�9G�A�d6�V��o���+��[z性2�7ѩ/z9��|C��!
@��LZD���z]6�����C�#�d�$�]�lz�=���t �F	�!]b�G�{��Vf������ggQ2U���
��1|M��f�G����`'�rֱ�(���dp���~�Rn�E�y��/��4�δ�X��ZM0Mȷ?x�,� �Q�[�>�E����ΏNf:����wrȮD*��cy���#��5A�S�e����<�{<����9�z*s�,g��<��W�;+�Ȍø*�`G(ҳ(�w��/^�"�̻�u�٧�5���?c���7���bW�(e�-^�XI�@|K�7���&Z|їhT�:��N��xUj�SHͧث �x��Qǲ�C��O��w�&s��	���o�4�ĝ�����=�i (���s,?�n��A3�a �y�z�*O�(���,��Cqayw,Z������'�4M��v,�lo�a!�]ڋ+b���jU��%�u]<��Q�y� }��� c�̑�c�Ӯ�![�g��m��I�*韟<�Ƀ7Xj�H�j��2��S�DB�u��ҵ���B��(��K��H&D6^(�鷄���@d.w��(���
AY{.��Y�J�S�����R��T}9��r2��A��߹>`u�A,��q@��F�������[���n���<ռ���N�@�m�؛��~4H�6�R=X�G	�����g�R�L��O_�Ae�yCw<5ƲvwrEw���l������C����x�ˮr��D��ipRV�[��U,������_�{3Z���{�=g&���@�Y�}�oy>	\f��)v�yBSHT�7T�����iߜE�2�f"�ۡ�pޮ8T��{�E �xԓ�Nu6����*����AE�dW(!��,�)D>�ÐJ��'����('Nȓ͔S�r��~f�zqV��u#�6�l}m �G��=g�9)���e�a(�H��̌%�C�e��� #՜�3~ԝgQN���" �o��>lD"����Y*Y�a��iϦ�����5�v1�F㛱����`\�Y-O��{�L���_:c�)�8(��ص�婃�s�w�~�+so�O(�k�4ܒ���ُ��VY�Q�A��;)���C�8����-R؇B�>��*p.���o� �B���')pc�
b��n4�~G�%$d�nH�G1T�& ���G�&� ��~\������kN��w}��e���*mB�Zd~D�w[�F���1V/�@r��5�T�=Y�)�~�)iFN���XM�'��Xj�pM7�Vt|�-��TfG��t��Gk�!0��0�Q�Q�cM��i���x�Ox[J��~<��_Blد��N뿆uI@@��9�� i��ra��8�f*0�ͼ��T�F,~��0��Wtw��Ǎ��z�/�O.V2�#�5���6��C�?�/GedEei��i�S-��`���j	};�B]�u�'{R����ڃ"K��4P���C2�ߢ�I͔�U�f	r%����i�n����l�&�r�+E���󗶠*�� q�����ã�!�����r"ؔ����9���z�%�/yާ��%G�9����J1?]u]��)�l %�j�AD+D�)$���k��Noˈf�csd������q��4+<ۙ���7_t�FU���= ������xS1����;v��p]F��3���y������B��cSҙ
q?�f9�"M����lS9�盖>L;,>|��p>E@��֐Sf�A�_nr���ܹ�yh|)�������̫��
�Qs�P���a�\��qRv^�T���Ib����rV��u���Π�{!_�MWI�˷̩s�):�`�'?����7�>�� hv�*�H(��˞�����ٽB��S��ej@~��m��vlpj ����;�{�x��B�Q���Kǧ�0�2 �!U�F����E�6	�R,�� �0*G5�L^eK�ļp�f_���,���C�s۞j~=J��.9)���/\&~���!�1DX���ϼx�m�7��Ή���wHZ�Ӫܟ�h���9�2 �c�ǡ�/NXw�.�XU��x�܍�@H|2�,������|``�-�Ɨ���x��B��V���h��d~0�&�4�3{��	��qw�>j�i{���h3Fe�	�5`�x�k��9���t>j�h��]H���h[���6��̫oI�1�,Kwlu�|�u��^��Ք@�E�50���x)ј�-ߟ0��Ș/nD���Y�z��f˲�e�Ϻ�<N�j)W��0J�I�&1�G�U����]��JPЦ:��S��q�6�]����KK�9}bҀ�SL�����@�5��\��;���u���y��v���0#�"ӓ}��Φ��X?.�/a�ƊΑ3f�N�	�CU���\���n��$ؽ�'	�R� ۀx��^��׃�lȤwI��#W<����CМ�����Ͽ ��S����9r�0 ��Y~��c���$��|���֊�t2y�~�c�͐bNq�]F꼜����o��iì���_m����̭���ǆ�g߀,�`��^'������������>w��3v�ϫ�������Tt�"�;Kt�9��Ak'>���Q�J�v��+��-��`A�|�)��"����fK���S]����lw��O�p�����WdQ	\C	e�oӶc)����$8Z"T���p��I�<���@B�*!�/I�$�YU�U=W�$��d�CυhHuW{�_�,��
؏<=�(^��G����b��<O�i��	V@��je�%3c�q@5z���`MF6=����$�`��B����x^��|���!��/�Y�P��Գ�����9�I�R!`7�7t�44���kj~Jr4��V��ъ4O��DR��	����H���2�wJ
Y�t��Q�&U>32��"^+�������|3Z�0AC�"�xk>�L1� ^�v�{z}����5�����9ݾ����y�I��G�zqՎ���L��&n�ӭJ�p���	�&�P����@�!��h��sZG���Dv[ O���v�����5y*���ir6�o~76�dɱ?�������Y�a�y"�g�;l�V����_+�4�U�;љ�u��C���`d���O�_�ڤ��t��C�{�1�Ι��(�z	U�Q*��S�zH�:�V6n'a������&,�5t ]�
FGz�<�ۄ(����A��/)�_'��=��L5���H��I)
������]M� ����F��tV3��d��:H2y��;�������N�Z�N�C�$��7�|�2Zሷp�0kG�9v�:���$Q3»��m�W�|��SΪ5X�,U��S��ׄ�����O��'R1��T/9��N�\v<H��|���*� 6����`f.9����ˡ�ir$$���M��YV�x)�ʻ�HYcM �Kvxg�v��9lC�<�I+.�d��Lp�eB�w�o1��!��[{�5N�YI�6r�v���L�d�X�3�3�J������}/9ll�I��� (�s�d?T��J8�P��*�Ӑr������(?� ��!m�u��uf�ў��CZd�ivy���g�y��ZW\���/��E��P��O�tr�ǽ�'r8�`@�5+�X��mom$ۀSKM���_�̡(�u8���_���W�gI;-|���Y��u�v�M�D�k�NHfu�P�'�UV�H	�c�e����IO�<���_.��(��^^�&�|�鏭:�d��A������V"�sIܮ�5��:��v�v�0��g����t����(�7�2����)�W�@*^���w1n%��*Y�!A"�-�4�a�J}D��N�x����t��3tV��yլ)��I�� �$Q�ƻ@K�"��Щ`S�n�@\GAɶ�Pֹ��48��X��W8Uf�V@RI�W\i�>�N�t�J��)�V7y;�8������U�N�+�F&��0T�b�=��q��?�����^�Kw��E��a�eѮ(�1ZQ��2�	��R@�A���
kȕ($�J�M��F���;�G��GS�mE�=�P)���	Jf%��_I�%�-
����˒I�:�3%Yjw���ƖZ��I֯>/�*���2!D~T�,}�M�}��PE�ɴ�lN��ap����-��;��@4�������.~r�UZ�y�ZkA
���M;�2J���e5�ke�R/v�+�w4u~�l,�� ($��6��I��PgE�SГ�J��-}���m�h�� �1'�i�ֹ�rCc�vg.��Jgeߧ�^M����h�H�G]�Y�xr�7%i���P�8;-��~��V_�T��P�g�_�������,?n��B�0yp\R7@�vU����	
է�4ɒj��6J�((J]��/���ӝ�z�
4�_�!�ܟt}(I?�Hn�������'8�I� #��9t :��s��9�͒\�tɼ�	 jhx��)��A!h����٘���-�2/�@��}fԶ8�S��b��Bñ����H�Gv����/���K�tX����<!
:���)����k��l>�����q���$Y ����{��Q��(���"�lF�fTΰ)֏��/[#r����_)�W1�-z�9F{�x`��c�j��r0K ^C?!A��q���9ڵ��HF�KBy�T�~�uұP.��5�0 �����h��"�0���߂/<q�~h�7��Y�&V���'�E
��8��W~k�7�j2��_��(��0�f��~+N��|tf�O�	��`�J�dYzX�r�]~3Ѝ��q:pM��n��3��A
2X�/��E!���q�[)2ߞ�2�h���0v�O��Eo����@�e19k��g�B��|`��Aަùژ3q_��
b�K���H�n�A�d�I�O�:ѵ',Z��#CYBC�� �PdB)7K���>$2�p�QQ�i���	�ܓ��'��wP쀤]'����g)�߸#����*�^�,jO�I������zg�EK?��)�_m)e!�u������D���s-t��ƫ1Dˍ���7b\,+O���0Paz��Y���H���{���t�8����v��[��*�v��O�-F1� �h����ҵ�-i�&�q��hn�ډBY�l�cj4JﺧQ�}:ePa��I�n8�+˻�vVҋ2�x���
aSK`������X��|L�=���,U+�n���B��I��h��7Ƴ��ћ.v3�e�W�(�5_{�3�"�t����{FZ�k-�����[�������sw��`��Vuo7(M~f�Oi]Pe�˪���Z\�}}|�"��<���a=��]׼6��W����V��P�����.!Ne|�w��H�������.��������l�3MDטp�R��%�NB��;D��;��)��^�3��I���r�9'��<�<�-�0ܾ7K.�EB��.�I`�4�s�2���
�1+iעk�ħ�����7w���L���i�;b���r�vA�����aW�W�bD-9f��&�#���j��c ��L{��[���X��}���Kܘ��Kϧ?*�!zh9�TE��q}�K�"*R��*RW��l���b�r�YP[�ɢ��97&��ٷk5WK�C-=Y�l/�Da"���r�d�J/��(�P._��'[Ӹ��A6,!�\֡Up��I!CY��غf߾���9�/�� ,)�;P��>�>��Co��'9�����HwU�r�S������3�a0����~X�>��W��
��G����f��l(��~g����J;��:���Fg@qU�����aWu2.�'O �����˟q�i�[�$��8N�"3��ȷ
��a�G�_�	�Y�ŠҾb�@�<�VM�pm�k��q«�V�k<�f�7�Ϩ)���oh���.)x��36񀑕��.�4:"�m(E���(�}T�/<a��RoEk�� ���J6��\T���	��!b�߃N&l�P��T-�Di��^�
�7ä��u���olb��R�N�n0)x�*)8�aqf8���0������5���>Ce�A��<�cH�������K,x+!��Pr�����~o��ca��kG2vX�����*�-�\�|�
 o���A����8�Dӹ��YS篦h)�\���ǣ�Ч��Ɉ���hD`<�a�ȴG9�8rEޛ
Ow���N*|�ݚG�L��g����?F<��+�02�[��鬍��E�K8���hiZ����cT�IW����E=�[;�L"�o#&W٣ܝ��y"*��LX)0�`��|m�p��S2�Ս�MhwT�>�(؍"��!w���̇�8���w�i�SEW��7(�����/*��`�|�֊Gm=�.ĵ�֨�?8�r��T��*�}9 �۽�lB�k���$S�Z���!ʫ�}�+�y�`�I�Z�*ܾ���3���/{�
�Nl����6���졯�<X,��j�	�B��H"M�P�o8�=��ye1�����׼F�/�~�����^Sj���,�,�q@�V�1ާ��+@0F7b|LVu�Ȼl�z�O�=� �����1��a&��P�IUq%W�r�Nx6�3���S��u4?!�;�݇��*��?���9��7�U�+���2n��ʇ�"�g㟙�P�s�N�!��հ}h�D�b��էy[vm���4����0�\�Gf88��z<uQa�&�����l�;�'Ls�M�� ވ��c����ֵ��]���`{�j@�f�^u6�����"u/p�z�8��ցT$�r{�o��X4M�/a�Ha��:9�@'�
��z�]~��~g?Ox��^��	��蓧.)�X�	�h��(1��~Ȟf�~_�x��͚f�:!����ۯR�=�l�����rx�Ks��Tӕ�.
��D�,U�P��u�Qͨ��$5�DB2>�M֚�8���ϳ8���e�k�QE������p7�c�W�<M0x�\Q��l�[ǥd��|WC1i���!�@Q���X�j�@����1�`�"`��n�I�|���iH��k��ZY�_���q���.�h�����P��Õ�zv�	�L%�R<t �7�n��(~�ګ�ªf��h�W��Z�Ґ�&a=U7�����H�{k��"�0���eV�ձ[����,yJ�9���Oɣ�%��]�0�eΕH�yV�f+-�ɫ8}b�̶R��6;D���W�ׇ�'���/�'|�ϰ��D����\��aӝ���wX���J�����a0���9�eU�O��\��:%{K �J��<q��o25�''���}�R�p׊5%a�"C #)��|u�KD������Z���}hI��<	_��ŦD?D��#�A-G��ʣ������W.���Ҵ��Y(��]���2��Y�X�8�I�mA\��n9��G�,.q5���l�0�~Z��j� p߉�`2�3H��V �O�T�}�7z�8^�s����@&���}+�R��K�������������?��Q0���^i��d7���9�!�!�ݽ�qĭ���M�#�*L�N�����wϓ=��'&��i ����������b�?�f�k�aBEp��0�t� l��"x��q��U�c�.�������i���FD��#�AÏ�{%��9*,��G���,�, ��wI s~x�h��&b���:/��R��lF|��Rg���`�N���U�����kG��%�MG��DW���+m���:X��Z�D�_��T7��i�k�1�uλ��]�� AfZ���JM!mݚ��g3S1�qIn�1tr�s4ZQD#��&I�9���W��K)�h;#����٭�Z�Ь�j��;e��ﾐ&�ʔ����0=c<Z�Ŀ����)j���gJG����AiŇY���y�I楱�%2�j�}6�%����+�i"x�⥮���Y|e���W#�e��gs��$�
�򅇼Kr��Q�����&Y�l-淁��{-|\(����[����E���@�#m#R%(�1;�Z{\6#M�)�d�°u3�$��g���9wr\h�R65i��f��=��@�ϛDR��xhlE/ݏ�A�kxr��&�#�eΠ��A=�K�U�t�ҭ���g8L��m���x���2�:��߷�M�f,b1 �J 5D[l?�������ia~�F2�,-�t;�T����& Z%���K�9��ꃤƅ�r�BwO^��7�/�~�n4��<0���۱�I=	BZiv��S��1��e�����%2љro$�����YQ����D�
�#�ć�c0����ln�\7`�8�u�h�A���!�GBĕ�Y9A�\������o��Q{⿳�]���	)#��f!P���w7�d�&O�͛h�I�2,2�=�6���q�B.�ғ޴W�dhz���}�G��+�/�P]�zw��(5%c��E�`���m���1�MOf�pu8�����CD~j2�I-O?���������2�zK�_����B�B?<㫥B�ђ��cp�Y�nW�lΚ����+6r�奈I LT�huӏgV�ķȄ�"4�gDj��s�ӛd��n��"_�Ώ��+���[�������3��^�b�,�+��	���cs���/i=.k�xk���8�Qi%)�ϴN�]��l�YG���=���0��|�!p"�6��[�3�k�R�[�#\8O_s�`��=������ ��ZĶuX[*�����{�[����18�z��~
����t0cx�쉸m^1񱧠��ϒo�:�����2�������j�����IC�L�Wز_���|14��<z-�@=ME�y�����%��� ���`�b�U!���5ԓ�S�ȡە��f�T�@/�oS�_~��@XRBap~+�h�D�JM2^��ڰ�5����<��c�� ���f3F��nF���t�h�}��;�C����o��I� D�����.³涴��(����.~F��GA�=hN)��z$g�kR/��D��kp]�5א�x��%���k�5�-?�nQMW�;	�T�f>w|$+�[�+� *ܡ�{?��v�A��ɯ�(*702�uR�볺:H� LN���O��~��ȕ�����wFR�Ti\�������l�#} �{��W��B+��O��`����q|���.�bx%�#�8�9k���νS�m�ǌ�Cp]��yt6I�I���:���*��j���_;���q����B��ı�'D��W�W��(���t�o7ڝ�;�w�����"�4acT?��A�l�;�x�\;��8������}�#�:T��T���fSj���]����%n'��q;�S�z�tF�.D��r�>�:�=�Z2#���r�э D���!*�_D�9QĎ"��W�������� ���v�ۂd��v ���}cDu�3�EM]���w$]/�B��[a��l��
�~�9�F6۳װP�����BC:Nh0��z�0&�^.�a��ܮ��Dc�-&�I�p2�q�!�Ά�����2�;� `k$`����o ���-�H�Br�P���̦�9G��������$jfG�'�T��S�pV٠��)8�����s�Ɖ�W�(��v�6��ς��)]�[�L�kG��Sf_Q���]�
��>����N���%�7�Cd�YWg��Kz�E��5�h��I�ߗ_���vI�:F�R0�7m��V�"&�¸8���_��x���0��^{��J?a��!6��}��tAJbPw�6U��y�k�؏����t5�>�}o�\�����չ�����7J.�&�'�ȱ�VAT��,����@�.��]1z
�7`H�`ǝYS�ݐA����u2�[�C�a�Ϳ����.��4���΍�4KV��(=�aR�}�ʝ:���/ع��?r�wg�*7b�V)R�v,1Gߤ3s��$�M쪴Z]����w�a:r�Ɏ�[�@��_-�}�"��_��(�H�z��Hm�̹�J�܉����T�����P]�����37�z&"���D��g��pT$�V=r�=M���Fc���I�[Z�浝�Y�������$]�Q�%f~�K�?V̅��-s����o�n6���P>a�k��"�����ɥ�vAp_��f��m��mO�oVKF�y�,n��CXo.��ǴI�)it/�n�!cظV�}�X���ʤ,�n�f��`D6���m��JH)�����^�{5�,�E���S20�Nt�{��n�M6,ͧ�r�߱G��n��a����g�2��"�L`?��3�-G{G�^
�`���{��hѫw�=�aX���>�� ���ͦ&ĩ���1�h$�"R�6��ыO&[�5t�_ӰYx�(�<��؟� �9w���*8����o�TF��5p�t�
+\|�z/{,�F���ẓn�ۚ}�j{�0>*O�6�撍i��'���^'���Mq��j"��w`��J�Y8�K�"?�^l�r�8�p��sZc�r������-����r�Ǟ�#��T�U���zyq�dWI���r�X�u}Fvf�����p��:Y�g��j"�m�m�q�ǋ�C�Z횝������m+g�
���_2�N F2�?˘TH���N����� �
�A/
���{4(��,�����ˮۻ�?~��y)X:���%�PD��T@A�I^b[0U�,�q�%�/<a0kXs�HoY��JJ�:~��rd�.��s���B�ћ�O�� �P���A�gw���@��Sk���E�@��Z\�XG�|2'��_�ߛ뀟��Գ�
��R��W�ui���f�����Τ�z+G�n3O�P-pf��cݯ:چ����_L-���d��F�Ks��,Fo�]�{S�J�Š_\?�~���V�q7�:%���A��6�Ru���:εRj3�]=�I��2.�ڭ�&[�N�=A"?��GY������u��V��p�>45-^z�F��@�?V�|��w��$ ���޷��b�l���K�W?��O�Ƭ��w��1����7�g�7_L�������t��%���.ڇ���Wy0_o؋��F}laܷ�ЍV�����EG��)��۽���c���7���#'y��j��؝"����<�{H�W4��g>/O�i4eؖ��Y�.E?�ո`u5o_K\=�R��Z���iC��n�B9LZ����9�^�����x3ߵ��P��_0s���v��]����g�*`�#U%��O���1(J���^oTo3��NFMC�3��Y����N��䠱D���k����6���_���4��>��y��=�c�d1N��3���]S�?�G<���������o6��Nz�/��^ŜB���d��o�YaA��#>����5�T�Dã�m���Z
<�"�C�����,C�9aF�<��ca��]�)�09')%�U��{��!��d�E $穹��%^��c��啕B���ɓT ��2��~ጼe�[��c�h�� ğ�.f7���u�-מ�3bwC��jc�es���f�3�̵�'�~�z�!��"qFf��\�.�Z�-6�}�F���z�b�(ˀ�l���Q�zx�$%>[U����q�����7:����.z�K�կ֮��|�!)��h!FE�e�_�O獠iq7;���R�:�8=M ,��TQ쐮w�\���g�D�"�����UL`��F(+s��9~�`���F�	{�i�O�2m�^-=d�ԁ�N�<I��L�}��[_��8�zs=X�
���oD��+maY�tO��ĸ�l�����3�0k%h�(kѵ����gab��|r���>��S@
�-�~���iGz��:�a2���nAC��2�
�)������#��)¼b����q�喩8��ڏ������-�/�M�i����J�w���	 �3��H�'o���F�4�$x�t������U�!�,�hN�Y~g�Y��9,n�~� #"�#
@��Z��V����P��z�s�U~l���)�u��,n�Oa�l�L��F��%���i�+���_��dD�}҈��M���Q�<�[�3D���o�[���k5n�dJ�H�P��n�]���^���m���5y4��q�t�R[09 ��Z���y�|�uQ6����t8�W��&{T����B����:�*9��I>��"$@�w�ۆ��3t��&=�-{�-�)��5Z'`�ɚHY)ԇՕd�O�Ixk�e�U/��o�]�5lHv��C�!<qkW,���L�e�1İρ0W\�v ��5�~�|�P��U~����I���0&�#��:DJ���9�X}��Y�^�3T�n]��GG�u�.�s=�I�l�a����"M�4�f���WEM߇əE�X*6��OS�BL�{����ez� �k��^
���n扅�(H��ZjSuO�c�;,F@}%N�J�i�6V������$���P����9�
�]�~�2"�J1��j�@�p�3 ����4��xG�'�i��M�x����lڑ��1��M8@?-z��E|�v�#C��g��LD��gq�s<>aNlJ�A�{>5
��P�l�A����rK�-ڥ�;|�\���`a�E�����r�_�9Q^oԪ̿	�k�9!� /�1�P��q�C�I��B�ؔ�5��M9�Gg#�*��m":eG�s䭛ݯL����m�{��@���s���̫���"�ȫeJC�A�SU���?�J��O��8��x����M_|/ա��,3����>t7_��c����ǿ�������ѯ�n��+�Ѡ( L'.�Ŵ��T%� I���
���̴1�Y9eO�cZ��T��$ �\�'���uV{*T�sˬ(����{s��D/�`����MK�w��5C�"*0�f��Jt��WT:��j˚�_��+���ڍ���8
����w7 }I��6l�
X���������Ͽɬ��p�5��G�OP�oTvr2+	p��g(�ԏM��.��}�lS�9{C&Ɠ��t��*�����"_��L���":��!?_��	`�	Q�@���	e���(.f����B1�����h��V����6����+�D�Zf�Wq �I�w��>Orц���Ց�͘�F	�AVuB1=ꡡ��Y��W&)诺QJ^�;�]l�-��QX��R-�b7��ę��mXx�Fh_�b];ށ��]\&r���t��� |���2���X�d2u�� ��1��_Ѣ)�*���yې�خ�f���I�F���Jm��%o%,��5�Fʱ\�\ѽ4���KW�;�dQ&����K��}����Nxٺ��F��Uf�����M���h��͈��A�"q�^�E��<7�6���^̜��-U=P¥h��#�Xc�LU�#������Nf;v�zI�,1���t��5K#m4��Fc-'�I�;^��`Z	C�{:N<[^'��/�*����㑂m��?�F�{�  b�B'x�;}j`���j�H��"��Q0�N�m�������Ci~YшR�=@c��V獪q�uO�\�)dS2��߷J.�$L}[����b�/t��}�qQ�W���a��s�t�-&h�WV�(R����}�4B#�#�r'�	ٺ+K;��m�4�-7��i�����=��T<4��7,�C�o�z�>F��T��H=�������7$'Bŉ�jr��'ܐ&�c�*u�+�,8N��)&�y�$�ԯ�R����N�?\s�J��U'1��Q���j���P�\��ln9�N~����PoV7<X�S�M�7ώ��]�t�%�I��m^3�Y����}6i"����~ʤ�7GR�F'�;lm�{��k#���l��] ݆�T���7b~��p�bУ���&��;]�Ϛ�����b���%�]ؒ�I�qi�U:�L�5�N�9�R��U�,w�nR2�l% 3)9=�J4ͧ� ����I�t ����Ӄ�H�2�+���Ğ�,eE�M�	(��-�L/x��P����
TOC��|d{�e���I���@�y]e���Gl7�|S��z�[sY��VQ����3� B�&A�Ы���n��"��^g:������E��tN*��7�:Y~�nm���<1@D�d�i���� ���v�D¹-����Px��_���b�88���>�� CW|��+�(�3���������h���0�L՗f�34Կ}���[�p$滘��ӑh�u6{iY>Y�����X�]��V	o�'ĚY�AG>�F��,�!B��/��DLL1?!n�Eծ�֪{�v�⢑g��"]���f�R���Ŝ��^�1c,&]<WM��x�er��D�&����	j���ǌƋp���H��;�"ٽ�eR�7�JN�镁����2qUߘAgb�u�^�e��d�$W;�L��pLŒtT)�k��1� /�@7Zo�I����p�ɱ��\�W?F� ������.�!�If����/I�%�A�X�2��{@/�y-�%B�X>��k!���gF����}l���C�*N�?�,�>��M)�)i3��m�3E9�Tb��(`�#�3�~ع����hR�"M�H�tQ~�FqXP�U ٶ��}9s��A:�$HrLkxg�$k6R]=/�%�t�`�;^~|$vE��A�<a<=gߴ���ȜĩR-�ڣ-Ny���1-� #�;,c�۴��3�7��=c(�=2V{pZ���eE��^��,v������9��?r�3^@�hJHߞ�ev^���q8k�_ݦ�#!����nڠ� �˚Ȅ���_buR+8���=����m�)�����9�ӽ���ӛ$y�3��h�Aqg���]�?Ff8��II��-�Wͽ@�ɤ�M�;j!�&O'�^�N�:�� ݌=�z�N�;1�20�"=:�S,d�ו��8�[�픝�a��{��I���Xa�p{�(���CW���s(_5�D�*�?�_5TW������
f���������*r�zN�k����[U=�S���A39I�(����3��H�^����*B���{��n/��f^'�j;�i���J³ǎ	P�N�kXl�J#4����n� �1Z��*Tː��n���t®9��3��d9��z_�F�� �$X���!�P�����ø>}Rc��ꍔm�)��L2���CT�"�d���B	���Ivt-(�>
Ҍ�h�?C��ٹ�t���<e߭#�DMg>�e��ӐX�ʗ ���ȠuB�y������+����X�/V|�"�������%_��@n�g:Y�E����6p����ӊ�q%N�4� ��{�Cr��҂��V�?L
����;.�&�b��A~[f���@~�@1��g��+�C�HX��7T�5^��y볓.�����ls�n#�3/V;��������E|j��K'x�&�F����Jxq�[�6(�tp�Ĝ��p�5�C�(��.5��Fu�b*�����WgU�>C6�hu�h��BDO��Vʱ9R��V�K��kTdwΥ�٥��C���tX -�3�f�<�����\�d^��n?��rv�E�B~�A��x��U�����s~�Vf��;������(1'�
 b#1�����?f��B�a��_�O��@@����cI���H'E����
nZ3��2|�Uɘ�9%&;��I�j��[�G���x���`gp�.c������c!(�t$���	�KvR-º�� ���+P�� (��p� "��<�4ٳ����{��.��H,Y���:m�WPY\��U;�U�agH��5|�M�L�LT�V^?��8W(�=2s�u�j�KS__�W-���%�q�N����l�$�	�V�����uWvp�.�^��U��A�v����C�]J�>�9��OJ���_��#��Ϡd�Q�^,�������� ޮ��վ>�ه��w/�jJ@�9��.y�}sxQ��.�N������G�#�J`8Y]���'Ԛ��!�W�lK)^�̼ҟC���4���h@��Q2(V�VS$��/�1���%�.�U��K�w�d'V���߄w�=�-S�`*��r�kI��eNS	9]��C�0�M�Gi��2& n�˃~��aD��<�����6.k+^Y��z�꾳@�ec^�����=��9�G����U]��P̞#�.{��5����iO(�9{Q%UGt��1�ad����r�L�B��*�$�Ǔ��3�GT�1����u�mSߴa�0
KZ1luc�V~�Y%��u��fa-d�=�2�e�����j���?4ͭ����폲��T����;��yP?�.ћ��,n˥�K�m��%�	��ǿ����OO�O��[����Ku�܇܏���	�$;Z��xp��=>�:�i;��Y���� �k�bޑ�~��ג�����F�P��'P���a��/����O a���{٭�Ġ1I�n��w�Ⱍy��MF�� ��g.�*�wqhV���X[��x�#�//��Y�I��4�}xwL��aC��*�.ٓӊ	٢����س�@Ua���ꜻ}�{>h'���(Q��q@��^����62�1A���"��=
�b����������j\�0�C�X����I{8�]"�<�A�.l���e5T����c���d![���Af7&��* �en<d�W�>߱����w���;�j�v)ɂA9B�M�]���
F����K&D�V�����\�L���+�ӈC����p�ߨ�D+,��_�x��}Ob�M\G�-� O��8�j����#�'�����7kU贱�@��9��%��k�RRƸ�ő-�O�}<��gb�^7u1�}��S�0X�w#a��sx5�!���������f�颬
�;�A,n�������O�}�\��x���V)��'�]�c����ңRM����﹄��GY��|���k���޾�tM�E�z6]7�4X���!�(�p6U��J�B_�v��|��'�r~k#���5�0�tՔ1�[�9u?��z��[��9u�휁�w�?r�ȶH&���T�s�X2��T����Һ"륩���PgU��KR1H���a�F������7VnP��9;�ߩ�����Vv��I�*��Y��~b����Ji��ܘo�-�k>�9g8]g���9Ĭ��ӻMrs)��i;�@���SA������|�Do�;�"5�I>��1n��'a
��zJ�`C�(���6�ٮ����"@b���Q^e
���'�+E��v�;�t1����	ak�X���h*�_�����W���r�ٌ��s��;d����y�!�`����iV�أ�H����JW��[����S���~ޖ��W����WE�d1�C����L1�&(�qe �p!ۮ5���Wٶ��~�d��x���7��e,N�p�\���|e[Iǥ� +�N�=�{U�<Sтg������gd�E/�����q,Ӿݑ�?au���T=VM:r��,������r�M#3��u �ۮiY\�S�X,��YX��I²ɾt b�6�c
%�UX�-����Z��W�&���|��Q�;�֋�b�C<�K��<��G��-����c����A��YTQ���>=ڏ��۽Ty�e1Σg��Ŋ}Q� ���d~��Y���`@z����y�]�vc�$�A��m���N��2G���Ȥ����(����D�&�����Q�u�ɍ�=ǭ'7#,�p�����f�1V��h�b�xUdR��%���7�����v�^g�w�|�_�2�����^����`X��P��F�kg�sd�%���`b��';R�v^�]ct��R���k��O�w�G1��)r�Zi�ѰnɭW��@\JC�bt;a��EL��3'�����D��LA4ύb�M �[����*�_T�ձ4B�kZ��k
���+:�v���\W1��(nҨ��I�f��0J�O+���*�jm��>=c{��m�=T�W=��{�!��6Dm0���n��NC�^�a:���Q;P$�B3�yWQl�/�
��;�kN�\��V�+�<3�C75�%�Z~[S�LG����K��v�&�\.��( roH>sD:�x�P�
H�մ�
��5�!�nY�Ѡ�&1Еh�_��+IV��>m_�o���!��TR���2ƨ����8�����Q��\�Ӡ��?�<��JT����Y>� mz~n�|�g� �G�;�
GQ��kڼ��
��Ӡ��U/��|�N
�Yg���_�ȳ/|�d�6���~�ؠ跞/����b��Ў�
�S��`
��v�.Z5�C���8��C�-ޥ�t�%b3%�ʧ�Iz��1X��և,�# ���.m��7�]Z{��:Z����&rڲ�c�\O06O8q��w�$���vn��w��:Ջ��]���!|�N9�����*$J�9�;{Q��ê�:,ҍ�M��#�'*6�x�����"���]��Jzء7.�Wl'�]~�@�b7k����ReVGj�Fk�W��$��M�
)�`9�מ[�o��^��T���ǿ�w�7�r�3v�Ċ靚���"���f��5����f���UN��G#��N;:)M���`���塙�Xt��7�&����%د�q\VЮA��˝;�P���~
��C�}1��0^�F�ņT��e�Zq �!�#l�=���v���f���xR�6�&d�':6E6�G��2�r�N+�.O����S��z�H�я��ٶ��Wqb�s�t�Q�G��Oa���FM�e���,f{;��p��g'�C��J8�wh4Q�U:Z�����e��K�ܼs��D��T�����m_�O��l� 1�3g���mU(/�))-yx'�ђ�~�c"���	�[�1�^�؛�5T��H�ؙ���I��,��k���㑇�|	��x�y��L�g������~�h��w�����q�}�fC��1���U�ᴦ�r~���$Tt0[���P�(^K��t�{a�l{�?x��&J���鄺\�6��9Vޏ�P9�}�ۦ@0�[˕๰��,"�|w�������Oo��7��:�2�bTnEȡ��3"�I@�X�EKR�ɐ��`�Ě�v�an�Æ�v�¶�z+�@[�+��j[�IYx�T��PZd�d���3H-(�ٝ���� ��e��u%R����������L�O�.~V��Ѷ�O��F7M���[*|�ar������oo�1끨���у��֕��p~4�ࡼ��B��}����įJ��jkpUN�P7�Rھ�����L�!�5�GR�u.�\���v2j�y򽂥�߸*�ʰ`v�?��	��L�F�۸���^$Q�ol�Wd=�IF�os�I^���	�����γI��F#�3��94;���CP���H?���R���0|���pRT}����ZOF��f��p���|CjW�\R���� �/�#ӝDH��5VX����`�;��s�]�5�����*In�qϸ=h+:�x#��p�bl���B�	��9_���F�K�B;Y>�j�������(�D��M���M�'?���8��;�!�N�ޝ��9���kBTb���Җ��"�<��~�i��A*yرV1����;��8�"'/����7݅=No+&˽�|�,~�N"��p��׬��fR��83��8��.v���B��ݡG���:u��k��O ���+��?)\������i��+5)� E�2G�3�TlަpMٽ�e�P{E+�!>�'�`���n�	䙭���ݨ���ǚ�\�H�т^���Z�.U`v?��{�C��W���]�gr�~ڭx�p�%��=s��1�iH����!GڐI���@N?otcSsc:�TX���8x���D-3�#��w�%ݒ���]_?&����En�{�f2ͦ��~�/ߴLA�z�
�YG0	�D����;��K7�c|L�R��f�lb�.��:��q%��}9���@{�/[��I�\�w'!g5�d���K0G�@Ag\�ج�>�Tsu\�P����]b�3��c<ZB�����B׮�4B���������L�O�[�e�N�Ɉ�a�x���en�s���[�|�M�w9@~��.Nv� �I��g�х+�M��� ����z2�g��R���ǩ���.�|[ú�E!�k�h`�X/;^�#֭ �2���zM}J�d?����qĀPl�{�k4\��I{��8��'WʀZ&͋�#����p=�s� ����~�|��a�*�(h�m�e�C焤m��Q�f
-7�NB~�ӡ�j�N������4>}�+�r&ES���B>��y<0d%�]�k�t�<�țQb���y���� �Q7��dYO���G�ɩuq�Hw0����S;�z��x�/����ȴ��ٚƩ�+��|ٟFf��ꖭ�Q[鲱��^~�ѽ�����2�0L{-�P��y�A��_=�����f�jq��'�94�!��`;���}n<H>�|�mٻt�h5���w��<Ճ�u=S����S�=��k����u&�y�Tv���jyr)r!;��:9�=|z�Q&�ͅ��h���o]/�grY���
��.��K�zw������/BsXoT�s�= /�zq���YY�1޺rBC%tˏYv�wۚk�C�I<�7r��q;������y=PN}�Q�^g�+h��:u�����r����'���?�|���]��&��,�̧����F��ŗ��	(��q�*_ˉq̤<�cq�S�mv���gR��p��G�60�W���
��`�j�O?f<�<��
�%Ť�/"�B֥�~��}��c����;]XT�� �^��h�Cp���Zy�GRe�U�Ob@�TPa0�HF�L�̅9i�D(��\���a)�j
ev�q�T؂ZK#�2�UԐn�O=�T:�-6i�TO������v�펀'}O�m��;��F(��E~{�yOE����<S�$Eow�`�q'Y�F��� �ۂ�ZqN$�
a)XvfM]�?~1�����黍e�OoY�U�����"ޟf��y$y�&���%/X� � s�R��f3�V烙f�/h�&3pFS�-�H�S�F�����!�������8�9� �7��;���c�[8�/v�+�Zu����`�`�����S� r������%C�b/����N<UN�0w�BS���\׳��D'�^=�	�0ֹࠠn���!�\XT:��DE�)UW|O�p}�g�;�����h��8B�e�����q�a�BJ���q�}�k���8jz����?*l_
	{�)K�8#�H�d�آOj��1Ќ�	��]t~�����ǥ��D��O`�&y�Qd����dh
�8��#�Fi0ad���͑r��Z���+���OtJ���k^�p�7���q�����hz�7�A�m>�ܔ�Si*�ƫ�'�&^�ﶁ�Jq�{��s%���֮6l:�:w)fݩzAwum 6d���^��a(_����g4V:u;!U�;˻?��X����9�(6<�OF/��r�!�~�`V��X��H�%��y�)�g+1GE6��-��,~�F���5�r�LK�$�`I�i(�=�����s�FΔ��J\8�G!�Ni}��g��
L��Qt��P|%�b�m˰r2	eqr����g����9���M (.�4�fO��0�}Ć�g�Db��(g�wC���a���u��ߔ����rU�ݜ:�i�zY`8�Y�Ԃ�gau�̌!��?"(in3��v�H~.�(>�pM����u;$,�K����L�ok�� ,������=�<�.�;ki���c�a����E?�K�9�;9�N(1�P4t�z)�8�Ē��0�L0�V��RLEA�@���we�P�Mh�)�U���*.m�<� ��y�T^��vx>��3j��t�o����֭��E��ߤ+���x�y�� 3;:E�,P77c�Y\M��c'�l���<%�M���ސ]|atUNEB�_��ۑ�{��jU�}��
u�u�+制�֣żWϸ�j�
�,��ޒ�x�,�Wd-Q7�����>���9�-A���{6�j�,g�D��F�5XZ��oإ���o�y.���L��b)����ʴ���o@𷦬�7j^�:�p,X�?H78Xd%TP���sa
>>Og7X�8�������=����g�ΰW^���9mƚ�)
�uU�EI�ۓo�(O����=�j��`�O����y�آ@<��av3bo4,`V�N�&#��� d s��'7��{�}D?K�b_���rQ����g�yl0�{��%�F6�&�<�ˆK���'fu��-k
'$t�,;�'�)[�}����ϙ����ě`�r���^�(י6��zO�����0��E��i�������N=�1>*T�v嘀>�:-t������������b(�A�]�+���Y��&ɼ�ULTϞ!&�Pı,�%�(��@��$��0��� T��f�	��qVH��O���[�T�Ԯ.3���+�얤p��f{����J%|3"�9	D�;_�΃��Ӏ����{��^� ��*B0���E�Ldl�Aչ32����T̜Gj��fo��}�cB
g���TN�-Nhk��,�0����N���r>@���I�M��]"�k'?���]��}�
Z��t��d����*y��q�E�y�B\ߨ��*���н�[To)H��ji"��l�����9L��@������7bdh����ѮH��w��9?�?��>��w:���3:D�RZN�6��5A�6�,8m[�J�Y?2�gX);�,�>��st�{h�l���V��`>hǫQӟ�����sc���༇���R~�*3㾑s%����(��gF���;iZ+�DIsj
x�hS:��ź?��r��֌���\���/�y�� ���]���󯶏��dl$���A�I��I^99l�j���0����<�"�O����".��Ɔ	�2�l�O
U���Q8�i�D��z*�n>V�?H���#���p1�x"\^)�u^��	��ɈkN����%�bRI��n2T�ܴ^q�j��-�pf�L��)#�(�ㅰ��@Z_T ��ee�����c+:̊v���X���bb������_ �3W�(���RWE�1a�Z2Ll
"^�C� ����(�ع�<R�Z�ց��,�&��9$�����)Q�䐀��s8s�ݎ��t�9���h��#������ݛ9tvtʆ�X�Y+9�|~hL
�N��:ھ �;�0ɘ)98�l�F�;���M�goT��u��_���W�.ы6e��r�o5���#1ס5`�9]���dwT:S��S����B��+(���ie �P:�fQu.욡VnC"ڛU5�v���b��)yg����1u�7��������0���A�8S?׌z,�B�b������?�g�"K�k��a�� �0sqa��
=P������v�w����n���oWY�	r�+��,]6�l����%�醈)�U	r;(����b��m�vc[@SڋM����b{|��{���J�6����x:|{�lg�ۧ����gXpN"gK�����?�z�#�Q@�"�5� \׃?���=�T͕�q��n.7X���@c����[���]�Ó�can�)�L�qS�C�q�� 4��il;�a�l@ MN�zQ=�^,���9����d�$�t߲��(C���0N���}�cpIo
è�wOK#8�AY��&8G�F6���Z���9���f_�AӚ���lϘ[��2��!
�=!������.j���ɟYo��9��1(A���Z<���2�/�`��vgq��7c�� �o�����ex�8�^�\�b:�8��XB�zm{5�{ڗ5R���3=0�!�A��Z��G 	8����p�.���EDa�0��t��"#ckI���nV�Q��O�C~핫0l�_�x�v�EvE�����q��8O�T�}��\,"�q����p}YW㦰��&�3gI�&�7�Ő<�Ġ��H�=���j9�W�c�)��R�F��<��=@ZzW�G�s���J����8�<W30��&�d�\-N��F�
���A���A�E��4!�Gҍ&9��SJ/�m�!! R@f�bmB�~�X��DE˳ڢ������[e�ǌ�Bu�	᷊ʹug������b8��\�;#]$n1���^��dQ#v#O-���c�}[5�JG{>���-��ý�u�U��~$"́�C�ِ8�J���
�Aa�q{�!��ڛ���3�ċ߄$���i\	�����^�~7��,�״:q4��,m�� i���A�p1�����,�]�(����!j�>F��D�%�h9�ED|��IG��(����o&W���������OS�U#�r7V��RX8�[��H��~���7�I(k'�2H���
���+w�����̀k���+o�6k���"FD`A��ߘ9�Τy�X�oH�TZ6�0��53>�T���=�8�+{l���>��~�{O|a�`I|5�-ƅ�dӑ��p}RdZ �e�S��?��*�3۰���W�lr: >�[18j^�x���s�T�T/#=0�8��+�2�G9T�D���w)�@Sl�8zr�ख़��V����Kk��J֠f�U��ՔwY��׍��ȹ�i��{�q�@J����z0�ȏ=J���!���k����F�N�с�u�5r�ũ��Q-�Bƅ_��oc�Jy�v˔|�	�2�Lck���q�ʚ'qz"�;O���N�%܊�~�?)�ɽv=�xD��?�J�&�,Ɗ�O����p��&m�=������������ ��*�>[��1IP`m�Z���~"j�����Ƴ��L*>��u/��Џ W�Q���%��������n��5/`Ⲑ�M�g�����`�B��膔�*-+hV+ )u�绵l�T�bOh��rX���fh�B踺c��6�B�	]��ɟx�~d������aJC�w��H� l�S5|�Iv��!�/� �{��;��<����U�X���h%ek-�!;������?��E�DD!���ɩ�fk�KuL����(p��/N�>�B�,�)�"D����p�W���I	o\��\��z8�`J~�{+Y~e\FKɽvZ�h��� �4��S�ю$�Q��U���:r��B~���5���+��{�?�*&ʯ?�����3gK��ъ%�'�7nzrZ�n���fQ���(�	�"B��M}O�W0��#B�Cg��'c�(8D^�p�L�b�jAeo~�օ�D	vL��n͐+�P�=NE��{I<Ԩ�X�A�ǵR��O,:NE�{'i��Ф�F]Ɇ��j'Q�й�	f�r2��f��wǚV���#����e�Y �ڑ���xR~��GQ��r�G���Z�Xҍv<��Cʸ�=aq�w*�%8:u!
>[*�I���3e7w���N5u���܏+^�)��|w���fC��~l��W���rOT��a',��zG '%4�R��
3w��e��p2�fS�a��V䌗���J�A.�Wb� C���}y�q��NG3��s�a[����N��c�h�Jr�,������DCj�����ϡ̽����Bc�AgЙ�>�w?=r��@�����gDhi��i��Jy'ֵ���I��p���w��L��-���k�i��^'��ۦ��Ƞ%�-�Z����b���B�h��¹��ۡg��9��:,p+�_.��WZ&�e8[�x@��'�EY9_�<��#��k,i����P����/��bR��r��V[��#ھj�(a�p�4 r+�d�������"HbX���r��XgJ:LG߸7%����~��ا?���n�-���}��A�Ѣ�(7��	���0)���ٴ鵏8+�}l2��:��V�w�Tk��xh]q�R]�<�n9����Cp�7��c��o�2%w�)�g;LI�,�;��`�cvw��&�δam-ݵP���A���Ĕ��د��ub��B��Kp���h�7��+7.l���\к�[̏Fy,�\�����/yw��5r>˿-�l_ �*��.ӊ��D!�"PFd0`����+�1iM{=�WW�.䗴�05+l��u�ǛAؑ�(���n�9nmd�<�"��q�
���t��e5_qW�J��������)z�8�����PtQ޿L.��@$|A^h�V8�v�p�;���+.oD"!�*gl
S�W�=��'�c�E�s��잽>_�n<��	]3պ�-�����u�Pr�wK"�U^��0� ��H�7��!^��gRN�Ll�v� ��=��}}�4��m��iYR�i�)0�k�9�6�lj �}�!�3d��3&�M�}���uL(�S��'y�ly��:����@'�k1�Ï|�<��=?g���^$��G
6�����s:�-�P%F�@��[2�Sc��Y>�-������Њl�&�2�~�����(�Uc�hd�u)ӫ����8H�	8������	�E+O�yj♄q�@��G����]�k��^���R��=G�J�~�١n7�}�0��[���nY�!�XO�۴]���\�ILӚ�	p'���Ȫ�9��;|�>4L%w@v���� ?�!z�w̱'�5�{|�R)�#A݅��\�������<W��!f�p��'��P�T�aE�����詝$��;��U��	?"�aP���!��fu��P�8�H[!��#�d�A�F ��\
^��@Bj+��&;kD����dM2vI��~V�w����{w��0aQ�*XD⽫:�|�P�-?�� ZP���"��vn�5��H�"vl��v}���<RV��7��f-�gd��[��r�)���X�G+���u>Q���A���u�/<�Jl����>�,��ݟ}��H��n2��� �4�!!o�/C����nq��=�'�:H�﹘7>Jc�����M<����Q�|v��p�J*����֜�A�sf^�ɫ��%
g's6~��}X�������Y��<��?�Z�K�g��u��24(�2�#
�ش`��X��3��Z�)�<�T[��ҍxh�8|�4�Hs�M���[���g�3��p�Q��k�@E�}.Bԝ�8�2��KfTz\�\F@ɨ+$:$9���ܭ6iU�$�:"� *�0��:�,�>�����V���V	���V�(�cA�Z1S������a褧�9nzjʍ�pm+��K�P��V=�Q�s�b�O3�H�t~��m��r+��9g�X�!I���;�i`S��3s�x>�FzB{���d�䜯��ǕJ�����U�k�;oE�����X<c��g�G����<d8�/�$j���Q�1Μ�+�����[� �z�0�򭌶�����q�qo�T�:����XA�#���$�M�uf�а��)��_z�Y�R�N��������WS�JC/Ĉx��ia��=�6
)1螨3�A��`��53՚oU�#��N��9�,��yY�����-�?=��y�ግ�"�}��w{�{\����qM�;�����ɖܹ��(�)6Ǜ�#��(v7�#��8w:���6s��k��Ć+��ݥ���T�G�;p��Y�G��/Y�Ff�D�5{���lNfH+�~=�lf��	�y���-R�B��'��a��/�c���J]����z�b��x���ҷI�D#M�L5�F�k����މ֎S�Y�EO��>Ғv@��¹;���4��Y�����BnU�sK�:*�K����W�c����Q�Z�UkO�8�ρ�S�P��W$R�˵�#��\\�.��� u[&X�II<��M�O���p�!ێ"+�On+�ݘ�C�"i��Z�&���՚<�n��$�"R�l��#`rj�=��܊��M|�hX���*�Q6М0��ɗC:������ ��=�����؍����W��LS��MSz�Q�_��dӸQ����'��cW�����뾋�4h�����u��t��U�Tʩ��G�i\3J�j�מ�y��h��;1��ۀ������+y�2��UV@E�OX3���y_ճ�3m����Y\���e�d��#'*��3������h*�e�#{��\6�`y�Ӻ$yeʵ$��8
���3����������
�*�"b�b=�|�C�St����C��Bu	3qД��&���ݦ�e�*�O27��G$*�v��=4#��B%���0|U϶�y�&)�|�����C���A~'n5�!w!�y�G����܏I��&_�M��xqo^��X��� E����ko9g_���Q+�k��M���g���WXhθ��}z:�}_Ja��/K�7czW��|��w�
l��J���Zf݄k��m�/�b�\�	?1Z,�an_7�-]U���ݨ��/zI�PU�&���%D,MD�s���J%Yu�[�O�>f���6�ۅ|�z�{�E���缡1f�':W�;��@�,6�\J��X�(̅�ܕ�b{d~+�x��Z�m�3~�.GUs����	�f\����|��/YSa���Z�U�e�p����,s�uoƐjPnSEc����\JU�A���й�2�8�X�la$�2Y�SE(�(rB]���z��M���Rve\�Utx�v^Y0biB���>�}�9q�J}�n�;4ye6ؗc5NѮk���ڢI����&�J����,��R�;�V�*L\���܂PЇI�p����N�ЇT�6J��r�xR�:�]ev�r�뢛P���n4��.� ��1x_�+bk^ZGX%�+gK�b�H���6V�Ϗlb�QgP&O� ~�P1����d�?J�	%ŋ,����"��d2!���}[w�C����=Щqd��M%<ͼ��ܤx�����Ht���N8��SS��g�ڋ��̺��ZH�U�rcꗍ�݅ _�đ���U�S��Zֆ����x�݅��Ai�P޹�O��|s'G�q���ѴЇ�"��_���
I��]���C2�aUr�A�Y2	�:i�ϴ�|)@��tԭ��W\h�--�*sh�m�r���>��M|��_���U�2��� x�)��U�$�d2&��(/q�ݯ	nD�^7�b�ݟ0����dQn����]b�����7��J�����D;�6%4��M4���뵤I�J��� t�����0fwD@���7�q��my�CU�=�w���@��-j��m{��-1뗜��X�F3
Y%�	oh�t��b��R�s���Ɯ�������|F�Jq�M�x�{E��p+��X4p8��z�Ԥ�(O�7ybn�N�ε��t�^�?��Zc�7\��P	�q��Z��
k"`��KG�t�싵�Ӭ��c� �_���E�W^ɱrQ�\�4+O证A��O���Aӄ�������'�0���U�1pދ�+hR[χL�㨎�t��2��墷�ժ+�0�tM����{�#�ʖw�=!��gOj} �-&=)�`'������/3��5e����u���昏�D��2�0w���O���"]\�3c/l�a�&�®��cq���B�C,���I�i�%l�����<R�o'���-�~�!���C��'h5ݍ�@cB�"*�ƕ6��Ei.$yB��X�����ݜ\��㏭}_B<c�\ME%�T���y[`9��`���Ib�Qޛ��B��7\��Ru�^i�w��e)�	M}@�0�3�%�7qdZ})2D�.Do<%�_mTį��W�L,�.q��/�q��2ډ��}��"| ��!�z8�9�FKnU�'��xlH2�h1���l��v�0F+�|��7(I�O���=���4DD��\~�	N3e��/"���A��r���lO�4{��]'�;�}��i�����4$?�J8�^2��P����|�8L�����A�
��Y����9�$���Da�P�w5�!��m�57/*P��r����1���o��F�uoa�`̵y��H�%�$%�,�=0c>���E��>�xk]-3��� (hSs����P1�6!����N�>�ҵ����߶���6�}N���+ج�u]Ri���D�o��������BcPcO�.�~��G�5^�1t�Y���)p��YЮ�����+d�|�'��5[l9$J~?)<����\��s���2-�VTQ�ͫ�u[���aH��/ɹ��t��j���AT�N�-n��0)�K�'Eo�e�AN��9���x���`<iW���O���+��;�M9p��s�b��e&��b��é.A�Ø̎�M�4O�&'+�D��d4��0�~���Dߥ ��]��#m��d_�a]�G""_G��\�x��y����{��ٲ'{��*3Y�p�&}L��{p��H�u�����ŉ]4o�-A/��#]5��:�J�oƽG�z�FMp��|�D=T�ń�w[�k0�XY�Û'ćg�@�����x����Q5}m2�<	ٓ��^�;��x��^Bg)-�X����R;��\`9A?Ӣ���Æ��Sh�2�7�_��f �Mh���z�!���B�mD�^"U;P������c�`B�%��L�h�A'岣���V5�	~(Ϩ9Њ�iw����b�T~�[��ʑߤ�u2�����}��K�y���M��B6�L�Q2�{��p�����mGr ��{��	I�׎��E�
�����w� 2��iϓ�aZ�0�L�H>�0�@m/J���צ�b����5�T��}�P��6�<��G��^�Q��Ɯ�L�q�[�='����?�f����P?|
f�2I.��S�L���J3��VXxg�U�iߑ\�p����l�|`v8m�8��AZcAڵ6q�<"i!�(�[_X��hUΖAJ�gj�jN�Sϕh��A?��3q!��<h�k�l����iB+�
�Ub
�}�W�ZK��v�Xdi=P=q�F
��f�l�MYRc�ܾRNzQ$��u�]�>�]$�.��{�3�Z�3�*������e�aMցk�m%}�i��<[i���@��.���0�n����3.�%H�Ûm��E,�CW�;�R�D��ۭf�7 ~��lq�izMy��M�E�R{�{;ngg-1���ų�C�*Xe��,������iȬ^��3H<y���YN���Q�檅�B��i�s�r��iβ�i��Ht��o30�9���^��Su	�){Ni�UR�K��:��z��K{�ߡs
s�!^L�!���aZ�r<oq30�(���Z���ڤ�s2ݬ��`�ԏQ��V{r-���F,Z��ḇNp�z�n�����EV�h��Re:7(c�.\<2��с ���mT�B�,��T�{O�f(��b�y�(#��^���pu1�w�Q� �,���ȥ}�{I����pSO|��Ll�:���1I�2��atM0L���wk��3y���%����� dF��v�ޝ#p��2�f�N��L��24i�vI���Ξ�ŵ��CU�R��:�4�굵�<���_r�s�
}R8Y�r�=�w���љ�Ç��J'�^�ݫ�7�	�CN������@�;(���~A�$�@c��t5����HL� ��gܛ:#Q
���/�/�'Ik �u��j�!ɚ9�5���sd]�9���)�l�~[;��z1��xu�4-�j2�SH#,��7�S�c�kI0�X9R�|�z�7�N�����?>'����UP��޲��4����⤿�V��vi]��]��6M�X/�?&4�Ƹ��17�J{�^���i �_f��d�RSՄ�C=�H�J�TEJ��R��-�����������m�;�@WL�ol�8�P9gAMj�S�A/������{U�9\�V�Z��>�����@mA�3�؋����v��I_T���@�p6*a6V��IQa�#�m.��Y�JP2u��(�A�����|CX�����Ki`�� � ���)(?P��s�?c^�U�u'�M��O�������8�Y����X#Xؼ�dYu΍�QjŮ�0bh^T�wH<j��I��s�F�W�{�d��;)�R����E6�_AP�uA-X�����gi���>���g�Jk��k�������E�,����%"�{/<.��/�ї'"Ӊ��G@v݉���Gá>8��;Ʃ.���k�O��[���^"�����B�}�1b~��"?�M��=[<Ht~Қ�yX�-)>8�.��K��(Ab�tN�P��#���a��M�a�mO�*:��I���u�ĳ� ���0潻)߻J��o��C3�����>I���]�Y�\]�A��?���hX�1w\WD��fU����R�.Wǿ��e 6#�b��|FkϧM�·P�U^�Ű%Y7�RL��}��l�S9� �6#ٜI�.7�GXS<:.lᜬp�^Kn���G5"�����h��8�c��J��V�����6ڿ�I�q�w%�9r��R6$(:�.9��{zᢃf��p�e��g0��n��?�0.�gP�h��q>if'���rz�1ȥ�@F3�Wn�H��R��aGPdv� �m��Z���c�������1v$�wʇC��k�dXj�.D[U�W?��*_�^T[��[���&m�u����b�OHf>�9`h�ҏ*_=j?�r8Pû�,a�\P�����r�p�eB���8�W�����̀���	�=p������i$:|�C����9���r.�D������F6 �3��R�q����м�Mxt�Y�h-uaF�в�5��S��Ǡ4�E�4)?Z��S�&�.���0���#�{�2�[g/�Sz�����9Q���X�!���B�
�.ҍ�\0��H���#���/C�����'����vW����[UV���0�Y64��@v��24Es\h5#��:)� ����b[�	����}o�*p|T
�w~ئRp���̈��"����Z����mn蜋��5�4�9���T�{������Bou݋�W�
J��J#6C&ϕ/ߵ���$팝��PM���J܉;�Ֆ�Nv�� ���!�3v����x����hӨ��N���%����֟q�~�I����0�9	f�.𪯨.��be3��Wȅ�ܙ�^c��@��n���q������A��gv��RZvX
��]�lB��\Q���w�� �a�`Dz/��A7��I�_2+K?/�\Gj���n!�
Q�!�Nr�[m��J>|��%�7�6�H���5^��5b֜��0r-������b����<�e���c������<�(xf�p�3�6x@x�~��ry���<]�M_?K� R����l��W��+�LW���a��Bqݟ�.�^�S=Tq-3�ȡ����.�I���RzCe؟W��W��5|}�Qi>MK{�\�ry��=��tN�ܧ�¡c,�-ي���5'����mb΅�-��Ꜥ���u۶��)���o
ás�Գ��¤�6d,b��Q6\��4g���G��ckde��{���
:Z��q\��X�޳O��Ct����2@^�SG�a{��O�f��&���T{��� 6��ٔ�m��Ęa��DTK���ݖގ�	�0X_>��[+6ȅ��b��-����9��J���j �HML�0�Hyi���[|�O���hw�<<����Ѻ��=����G�hV�8߄�!���E_���Ι�I.�{�O��ُ�6�~��/�U�~>�k�m��t� ̃GM����׌�J�o�U�+W";n�Es����Ke
J��$�&3I�I�	�[��U�{}�E*v�|{&��س$�6�Q�ԏ�WU�T����K��I�
}����&�3�/�]���nJb��:�("~āh��<QP���S?�>�
�{�|H�A���=�vu M|����Y(��O�6[�T-��y(���σ}��z�`٭��ޣgP*�O�ͼ))&�u�Q��Qϵ#�.� Z�� a�o�����m��LUu���32[�7����1�%L��VdJ�NR���vׂ[��>*/M�����ЄТ�Aj��]��*�P}�=7��cx1�UZ+fN�|$ ���RG�ȷ��)X�[��/n��̚��C'�A~��6^E���n��k�kC��;4h��52�{wI����?T�p�	,X�����5D��3�5����X��hG��S���
}�8)ѣ�b%QW2G8%�y�}B�� ��IۄJ��s�r��{;����E�l�/��3��/����;�&ލ��x��s�S��y���@M�.��U����e�y22�3���?��@k� ��k�c� N��x^�#W�x��R�k�L!�G��Ptnt=<����ʤa7���Z"M�m�aQֶD:)b>A�l��W{c���U㑶���!�O��1>u,wv��#~>�U��=��J�x��܅a�_y�+f�5�e���:i�403-�3�+�����v��򱰾n��GN`"�]y%���^Cm�6����S��j^ia�,��=�[�Q��o2���ljq����5
��M�i5�VV���ްO9Mo3���>@�7�Cq��!�k�� ^J�5��T���T;v��!i�ѷ�_u��a�蟪H��Dؤ���F�
�bN����U�&��N����Jhn�JA>v�2q����>�j��.��F1oĞ[:��,F���1C.p?G\D7���&t4V�|2���(+AS�"�s��)-��Q����x�h��i��*"g҃H��9���ve��/����AL[��ٙ�8m�a��Lm��8du�֫t�/�pcz�৤E�*6&m>�>��6h��N&i��E=."�4���a�I�_�Eb�F,���"ۑ���ワ��h$HO��[c!o���'l������E���S�,�ѯaW��-��
�֛~u}�WG����`�t��e��(����ǖ=��b;�Z-���G����|��㯚���R`͍|���E�|{�>�z^+�<�%/����W�q�MlΟa�[�YiǢ1~��y	Z������#����. ո)����|�v�JT��_z�Oy��#�(%�:�oD)����`�߅`���@/L����U��z�8�$��<a��\���&�v�nu
1�Yo���@�ݔ��Ҷ34��8O�]����(�40�<dg)h��!3�	��m+BMGL*͢��R���S78�>���
G�H��W�D�a�^��[	.�{�V��ϩ�s��RcB�[x�s��]]\�2�1N|0�|Q�Y��yo
Sb�8�oGG������Uz|9{*�	m�?"D�8�2�$�i-��bH|@t|E$bL�k	�� m�/B�@Hx�;f�*j�˽���O*j�}3̈́��8��DmBu;��	��G���n#Ef�ۋ��/�`�7֓�6����xm�r��ߩ{��r��%,���c� �#����Z�!r
��"v�;K�<zR���VR[7������7Yw��9�<nj���R��ٳ�!�U矋(ٺ�o�Ӷ���H������.�?;ߣ$7sJ.��Bɻ�cw���X@�VD�IG8���YP[�ppO���g����#:�\,�p1��W7/�MY��F�^��R8����s}C�O1��ŻY�p�O�k�m��}��	��+���#��W���J���(�5s8Q`��@�x#�@����g~Y{R�0�y�����O.��k��Q��[&(-W����v23^1�qش���T=�Ϛ�(W=�Qb������Nt	�B��-5k��hw� ����\e���;���)����!�.�����2)�~oq=[����\
�F�v�L�3��
�`m�$xY�9K��.svߛl^5���**C_$eH8��4S	�_���C=�c��ʩ}�l����F2x�q8����� 2Ptb)do�����_-�\�0Z-G�5��#���;��v�L!#N��W�}����	#q5t'�W@ꁖH@��<�S�Y/{H�`E5�����O�6�1R�9��Z/r�Ϳ �{V�L���)��{�Db:_�tF҅����dC�:�����e� �G�����{SBDǶB=:�l^��T����J�Y�8r�I)Q�*ѳ�r���E���s�?e�\	�6�`<;S�^'E��B���m�\���E������C�0	s}�/k�W\�<���OZ�_�¯l}�siZj[$����Z@+s�Im������k䗭���S�� Kձ������D_���1���	>�MUI�wp�sk��w�"��\�c����<�16� �7�f��PC�}{��I��t,��Ha*��+t�A&���|:KO����_Nd��U�WZ�#�R���G\^�O��K2��]o��3�S[2��O�������LP��O�:�(ī� ���`��:K��M.k U�:˻2,�s�s����}^��I���$J�8���L��,㠻�xД-������-��`�Gɢ�]�75���NÒF&7�!i�ʢ]��^�q���U�1l�c�m��B�L �S����2�*��F�ͼ�:��$�����}��ez�񇁘j�[�å��^�$��K?X������U^g����vcR��ǋ�"��>���+TH���D��G�(��f��bwiHu�+�E�s����=��#���`������BL|��)��e����d�]�>ۼpK�>���n%��d&�&:�:�+d�@�Ya����<��_/�D�&p��w�s.#�����Ӝ�T)�v��}���we��5��k�I���4��G�Y�OR6}�QlئOX~����ln@d]��o���اVOp��qa�0��C��b�Rꀲ��?���`���mE�S�zU��;.��p>14�iFM%��ma�������B�kǮzx�WK!��pz�~d"�1z���r�Vg���,�#?�j�C�Q��? ��ܽ�i
�C��JV����]�3.W�_?�����~7�u��Q�/N�L_(�O��/�.&(��9$0D�����;�K��X�jvW\n�ظ����T ��\����m�P�����HŊ�Ť|V\en���?8������L�H�E��Rg�I��{��`�N��qE��z' $W�M�?rӸ�S��o�H�uK+T;��!S�9�T���Ց�úDh2��?�{�a�e��
C(ս�f��*�i��u3�P�ȩC�û��ys�3�3�r���H�GL(٨��z�/~���]Te�K��y�(g	:b�JR�
3��3��qe;�;<[�n��������j�,�m[��[u즕!b&�i�F��t�A}�m�~���jq�#��a
��Pu�D$�F�	�!؊/����y|AK��K@Pm2�?!���D������ʴ�Aa�Oj��>
l�a�5��w�lE��p���GUb8�+�b�9�ND����Iڇ<7�i�'YN�o�?�(�l6}���5�|��ՊT��Z��Y�'���CZ�:���s�2�9/���XgFբӂKW��ńy(@-,�;аY�&�==��!�8/�sEK��J*L����*��<��
�	gg+�$<:K��:稃u�hf��ID۟Dyo]�S{�wP�f{�P�r���3;F�*�����'��,l\#e(J&�*5zI�:�U]h��d��B�f�u�這R�,�Y���kh3`NI��O�]�)L��U$Ŝ�ek�,�W�]��y�p^��A�W�����A-Z�:H�"/�=V�����R[���m` ���Gߵ�Qn��Z���'���u?�H��%���#kE^�|�v�駈����V8����� pWK�\N^8̛�'�+>�s�6ː����$������~ �OޝE�<��i�JJ��?�ʜ��V�k�D�	S\��Ou9�����?k@�1;/��^^�r S��s�h�Q�[_3o!�@v�`��6����P�7f�ዌ�,f����I�U#���_��2�85f-����>�y$��6�0Y�� ��\����n^�S���l#A��F\P�A�G�H�H!!�*'=/�߸^r`g��\	���ܹ�[��ߢB��]�v^��^�bN^h�,�w^<Fp��v|����lm��[f�6�q�oԑ"���8sPe�8/�Iʑ������R��������@R8���1<#5z�j4x����˷�"���w����#�����s�m����
*�6����Ad�E8�і^;�F��Eoj�W��Y�/�RK����iBHK<�O�u�t�ZP�PDC>X�16Vu�~P�2�j�4��A 9�;\F��NLgL� Opp\�W��~���8�H�@�A/e�	�V�k�0��I������/�wi��]�\�� V��{�{�5W_�g8,b�E�H.���_}��Ɵo>_`3��N�/�E��u!|a�6�K�s2�h�Z�	4��qA&�T�ډ�d�!�ʀ���/d�9��IT�U�L�Rh���w����z�zT�@O�PN5���7@/j��"�(����'���U��ԁf�v��"2�$�%l�F,��g�Jt�B������ԞB��̮Ur 2@���(��!l�G9�i([��L��{{2��L˥�G�Ij��K�X�}6҆`(�<����G��ȓI� Y��*����#�^gxQ�n#�U7t� ��*���c-S��v1����؋�E� �w�(����+�Y���5�t�de��hU� ��,��/�i�$鍷RBֳF�9��'kfk��?R�tr��V6�vl�b��XWE\��i����sИ��PG�C��8{�x��,f��V���g
�.oTm�b�G}[��!�x~���[ٹߧ$l��-`lU5oY[2^\*bFʈ���֋�
�c�K#�lP8�C�P��^��6{�'H�_r��4}��IF�������E%�l��a>�p��]��^��������~����K((d/�+)F܎�9�U��tr�;5��e+���`e��"`Y�ǅcϒd�\kU�&����%�iB�yh��\�:{.���+�i��w��,(VD�����^[��Y�|��md����b���0CJR,1���"_J����Oc�(��T��Y�����B��xԡ4����a$�#b8�mR4,3[��hL�����ő�F�������ʕ�XO��S��*�ȼ��xU����!Ъۤq����o�u"���ps�����(�^��7 �����mv8N䊚���f�հ�S�:��iU����y��I-d��'	��4�/b���z+����q*6�!y�C���^��S�[j1�t�m����c����wEc�w�#98?��z�����W��p�-A���,�G��9H��0��ʱ���{��q�L���ď��լ�>"�n�38������%2�C䇮���/���T�m����C��j�'�j)[����I�j�^�k��s_�AuJ}�8��B�{�����<ߖ�[�.�j��x�6��W�fk�~h?�ͲA{�*�ʕ��t�ę�4dhd��er¢�Ѥ�(�ZT�]�R���ǧ�g�Κ��D�7+�i+,oF��%��i�?���:�e�/��:����j��%�#��0�bq�x�x�(�K� jC����hCG˽��mG!tg�\ gd�������Ly�����;�6G�[�h��d���3.�ܘ�ug�������L.?PV����]�m��U�<��Z�B=ie^�p���;��R3xυ:�^�C�3Y.����+f&����L��D�*�����ޱ;ӥ��yQr�'nT�+� H���`=
wɪ�W4�����1o���(� ���>H�1���!M��4��I�1�
����yf�8�kY_޴(�ʹ�5��L�&;@��"�	�N��,�1���1$��6T� �^+[�t�X#r�;�<�O�$3Xy*�mr(��J����� �n�,]���½�fK��SD��>
-j?-4L>#I
>[����z�*\��1r�<���9�Ğڜ�
4��8 �wIBqT�Ү*�奰YF��XQ�	bF���5�0r/��Iل)C��l�9'�i���j	'Y�/sa^ YP�A;���˹mtLU"/�}���龧�5�|�����AS0��}Mk��MH�@&�"�l�(��ͪ�M�z�]\ W���_��=�(j����r� �K����@��x8���r�(��
�\p4.ƫ��,�����mT���@��fVN�`=����$~-�{E*���?Ƞ�N�f��D���REF����~c�"&���=dw��خ�%.�{X4�=�V�.���/�����mJ�����Z�a��)��\�E�
�Q���ֺ��^AV`��Um+\G�VT$d�Q���y��άbx[uG2�%�HȆl���7���/����i/���8t���8���4G�^{'���W��Bt	�7�^��LT#a=2�@"�\�]�� �b|S��E�/մ�A��o%���,a�͒3�/�ї�N%F8[1��m��W���=ީ%���&1��������Fԣ�Ĺ�ju��Ɲhi��$Ñ�>�[,��D{�X`������w�WC���+2F�Q_�	��dqb<�p��@rb���Z]�^2�����ƄL�#n"2H�v���eW�mF���lzɚ��R����U	��%��$E�Z�����X$rNˠ�ӕ�f�
��Yv��$�3�b��S�������J�A��XU�Fs���/����I�2�~��	�/cӨ�3�i9!Q���%�����C���hrƀ���&�J����%/�c���
TGN�sN#�D"-�$N�;��Th �D�L���|���/j�f]��m1�#�vIN�C�}��p����-�[<CD��v����Z���Ky�$�a�0V�ڽ�ٴFW���'��������
��!5D��ȶ*�1Q���d��e�@կH��$�#�k��PQ��[�v9�N/��tt�5�e��� ή�;��9���ƪ���7�f�Ƕ���G�@^���{�f��16��t�o-����������̂�L���9@-��S 2��k�T9�b��1�;"&?�ߖ���1�	�gUB�F���$V`Am�)~�!/�EpD�t�~�>ʶZ!Ga8���v���t��ZJ_1纋U�|����i�~��Xx nR�N��ת�}��|�H�f��v�����pf��K���4>�W���YRh��f&;ȱ=�>W2�0DÛ	g6+�0�Q7k8�YH+f0�22D��z�҆�fӬ�ثz�Hy.̓j���k)χ���{w?5s��I����	�v����!���ٮ[�����C��M�R�7;@�0�"|�3��7���RC"�@��xer�>�M���n�AW��K��ɝ�^V��=��s{�{��w�1���5>d��^�hG�}��љ�,GG�V�;JE��Q�<�O���u�W�B���A��kP"1��;]�̯�*~Dl@d�lVfm�:Vz�FK�o�>�Y�����ׯ��ݖH�q�ߘ����Dc��里K=N&zˁ�KMK9�����O�q(lo���~��eT�v�_��2-4,[r��^��/��N�;�^�>�2v�kJ��:HY����$gA��9e�����6E�1�be�/�B}�F����'8i�]{H����
�#���S7�h�L}}�7P� �B�ׁi�v�^|W+n�w�h�T�Edn(QH���.���h4�\/�� ��w�rh�:����5��+�(T�l�ԯ%L(�����ș���!��P�i>�F��cط��("�/5Q��M�1,v���ҝ*�$d GM�^^YٞD/r+����s���9��+��xڴ��o{�[	ͩM��/H��/CyE���kA-O`o��Ray9r
Zz=*s�ldI)����Ŧ}���[��sd�`�Ų2���$77+%�٤_B�O���2���0<�<�#����{A�G�A(����<a�z�O�Q<7}���f�rKʿ,�o}?t�yL�d9R�ǖJ�(h�D��H�U�����IO�n%]����h����;�Ǐ��+4YCe�_D
��93��2���t��ްq�9���0�x����F��!�NET�Za��گ|oO�vOK��Y����S�5?�jH.�!bx�_&Ug��iP����wr�)zOf4VߥZ�8||�k;�:��yJ�xՅ ޒ��
3Y2#�p�\�gn
%Ib�k�����[���+{��ַy�X�Gg�cL�����D�C��'��d��4ڮxY��rԘU6�D���#4�����4[�3�k$������H��{!�3��C].��x\�Q.�Wƶ-H�͋�Ͻ��aS�.�F#�'�%"��-*�ƿk�E�h�U�v%.'4T٫q��l�窘h���7�����x��Jd��!LH+%�&v�"=u���x#��E��@�p6X�c_�_?��!�����*�����|��$��td ��7M|��t��������H���I��	+Qn�g��y���:_wN�3�ٓL"��z ����&���sΠycӶ�GRL��s\t�m�����B�� c`�i˘ N�pz�.��}Peg����QtVK���A0�Ի\�J᏿9<Rd�b�T��;��('&����dJ��-Q�XI�������������\��j���!w+q:��q�)�� �8v�������jr;U?�g�n�ys��'�cD{"��3V6�e5�jE��"j�Y��O'}]>1�5j
W*sK�����Oz��A�b�r�L{[2S����S,�i�\A��C�C���4:|�(�/F�_:D��#ۂ��W��:��s��9 �;�Զyi����V���A�f��>i����%�F"���<p�R��8'۠� ��&�t�E9�+q�e�0n�H��B����V��(�a���}R'^a7�G�buC9�g] V�a�K�r[Q�;	�7?�VrF�aa%�hD�%D��X�~�+�p�Oap0#G�����$@>$�e�L'mRIU��pv�X���-����e��d��������h�	���<=IS��?Z���47��i^�+��������q�RBg��eSPa(~���@�!�#�ۻ3(��yh�)�h��K�$��b�ZI?��;~�H��K�%:��ϷV���#��ڋ�협�[ݜ�,*�������m��x����c���2��c�p���M�D�n��(���¤����sβ�g��Oe�d�<��4�L�ەx���H �%�j/\i����f�u�Ԯ?M�������9�Bo�:2��Z�>�:9���?7);Zd�BuG�$
��H�7�o|�e)���t���m����ŋ��U�y �0�ՃA���s��xk���8��Z�b�O띱vT$	'�P�봾��N3�;�ejp~�
R���  Æ���n��,�hmb�Y��0���W|��^h��D��[��
�:���2�Ҙ�c�cw�r�J�?��O<��NJCp�#l��6=+��F�ǹ��A�x�A;-����c���ZM�lM6lG��X1�싷��w��WH'%[�T�k�H�J���@<�L>�zR4P�J�����:9���1L'��)�ǅ=��1`��jU,��F�Xr�<��O�>�ci�j�3)�!�8��s�"r5�H\P��3U�r��}������-Ľ�JQ����8v<Z-N�= �!��d�b�h�P�];��9z���!���&�H�8� �'I��C�0S꼃69Nt��#��D�ZKSU0ر`��v�vy��8�!�v���큋9T�Yڕp!��u��.�����(��eD�0J��|i�`t���ef���Kd�K/P
��٧s�Q�`]�l������A6H<t�IL���g�fx��-��L����� hJ��~.fS&��/�:�urylw�3��q�8©�+/*�i7}q�ޞ_d�o�)1s��m!z)ͤ�����PT�غ�����>���L��U�U"�?lG��BskS�c�0���֌埆�� �@R�jm�$t�����*$���8�m:�լ؀��[��V��Sz�c0�lV7k)4 z3����u��苐�,�:A����"8iw����Q�5�r��5k����G%A�� �)Sw#�|.T\-�$E�Oz��8a� C~�Y��q���.Q'�ȽB�в�VH֑z�{����(4���u�5�����"����T8��*��ډ��>� ��OQˌ��jҌ)̧�9�x� ���a �z�J�Q ���;ҟ��ԛ��\�)W�����v�Y�}�}���(���l�@n�Q-q��]!����� ˨ֿ�A�̃O�\�Ub:.=�=�wC�����)�)��_/��c	}Ő�i�(�W���vfJ/"�XWR%������:����.i�b��mDr�����)kZ���[�1?2�<ǚ�E𝸓Q�1��;�8�
�M����G�����?���<�-�
�?�`��DP��!��=�"����|4n� Ȓ+��B�WR�'B�S�m��>�+�8�E"Q���Na��q6��s�'FI��r�5s��=��e�8	�4��7�A4S�!�������e�~Z#Jk�1s��F����2�4��g�c�����&�oa�o�2/�+1�����<���+ט]Y�-�����V={}p����)}�?~��j��~⡣օ�d-�S��>��32)��N�.���(���*�*���s@N���?sd=�?�MV�����e�L���X�J�ܿ�Лjt����Ծ�v���|��f�Tc�#�@��,>eO�Ȉ&��,BH=���	��t/�|�Րέ����jcNv=%�I� nV�����➄��F��i.���~+
��[��ΐ�ʘ�<���d�x�W�H<F���'��h�7%/�҅�E��BQ�9�%���
���]D��x�7(ם�Aa�:�tr�()0尮>���+���0��v<%K6�x�L��X�f�ͣFZ��`m��H��X�j���Iր�2�3����=j^T<<t$L�	8s���P��M���P���S��*�sF�K2��|�il*�5��k�����3W/ոَ�zT��WC���Q������Fk��T�5S#��^�����8�@a�@Y9�a��(����t
̞A��7T�|�2S�}���>	�M�*���m���9/�[(_�Zij���*x �����rM�k��"8��JOF�e�n���8��-	W],-:hmu�\�NG��w��a���}5w��@+SF��������������x~q* ?NB'����O��ѽ]�_�N�`H�-c���X�_�C|L�*�끗���!�I�8����`u#�޸>�P�n/�k�R��{V\���R��mz���ThӦ=�b}"�'Mj�cs�N :?�-s�IN�r������n�=K/�~���%����X��(Uj���
��:ص	p���^[�KQ��X�vb�,�2��W�}�k�>m���<H����4e�o���k"��)i~Dd���)�C�2ٵHՅ5n�!$��3���"�Q�C!����ͭlZdU���c:y�w)������tO�;�R�LpW�ʧ�)�� R�:ܯ6tP]|k��`@e���6+��<FA�� 闠@�Ө��z��O_v��~���\�jъWA��i�+w�M�]c��Z�k� xS��˛ֿ�BQ
'��	AMVb�ֵ����M~~�����.����~9{��M����)����U�جk�I5�O��m/k)B��֠��e)��+[�&@%)��B8��r��w��كI��7��e<�F
���L�ل/� x{�l�h�+���)v�'<��y�����Cn���5���s��^�,�.+�U=��gC'�x������Dp�ʋ#�}��j�6��Cz�3�*�
s�}��Ii�٥0������a��q���d4uŵ ���͵t����L�l���	�Z�؆���vpSM�/��u����2L����FY�LD.�˖�� G׫�;��]�ѕ���"��V(�����S�jbd��N`=����
��I����F����`�nC�``�f�0���1Z�I-��
c��Y��h��
k��s͢�����#�{|�/��ð���5�f!��?௏�P �G!�����\��+�7�l�[�����!����z�}���p���.������5U ����<�D�P���֠h�g����1l~{���d�ܜ���^&w�Q�)�/�I�1	�#t?�b1D|��z^C� +��"Tδ9.��-�
?�3\q����.��?����-w��)|���^#���Y�H{�M�����n��9�SE26 ��>�h�ԧO �A6��d�(�oj%�J�{�+�vm �AKp}���M-��m��HO��˼�F_s�[�e��L�]Yѷ-l��<ބ�J`YwäW�O�T�x��q�%�����2�P�e�*c�&F1��&��P�!�i�OĈJ����Z�$ZTamDi&;䂺߯��W�_b��W3!�	��B`�7��-�\LBZZ�G�sҗ�M�@i;�@�k7�96��q�+� ��Z�Á��8�Tѹ8 er��GN���D��bD��_�Qn�~{�(8������5s��p��$ٟ���䲁�5�5Ob^u>�.�N�Ov�r&E���h6�H~�3�ے�b�`�y{�d���g�wن7Q��������gIKM�\�K���'��<��G42Rb�<&��̠�NoA��T�Cj�����A8s��`28��*G��K�
FJV+Ի`����򕈓2dT��g�J��RE�5P.Z���4o_��[S�H괗FI���ۋ�#n��Y��<:5$l�>�A�|{�K�ae�vJ�8���w�G	8q�����Ǿ�}ؠ�29g&���"������#yLy�D��Oe�T�6����>-`?)t�c��sSX��|'����I$'E����|�ԍ0�[G=���_m�TI� ���[������x��s�=sp�d�a��0?g���l�M�ƚ�G1�9��*���G|x�a�n}���晉�d�4B�n ���q�b���*��M���Hz-Y�/�5��NU~+�n�|	�v֗_�]͜�1�LG�^�SGS�j�ž��2H;k�V�v�4�Q��� *�ǌ��)т�(ة14��ǥ�z�Ʌ����w�����9�06��?_��/�vg�.�*d�W�� ���^`�1Z��@��g��+���M< �#�
Ʀp���Q44x�i�)�[��G��}~���T
}̫�0���H��6�"�t�������1�
���$���o.M\�����-PA&YNjU��V�Z�}Ά�+���*�K9nIj��Ff:��i���>���d�[�d�b��p[Fҧ���+���Գ��XD^T�� o�g0�=������k+#�u�6�q��.���G�{ϧ w�^pw�=l���#5� uS�Wu�qp�N�4S6J��u��ɓ�ɍ�i�B��s2�ۙ�D����LgA%�-!��X@4"K�o�%�/��y�J����7N�@�={2����P��k��/U~0�	�8�p)�%����K��$���������T7Ҏ�~��8
�����^����{�wNZ����l�Z�8���}L=��]��[���������wx�����WO�y�tى3۷��8ޒ.%a��\�#�nE�D���e±B���52�HN%����\��y�P���Y�ft`&�72��C	b��#u͘�
1C�uj�\�����Ů�-#.3��";HB�rA�h�C�v��qz3пR��K�a˙���c�=ij�:c�5x��F=���L<X��%�$2D��xbE�e�����������$a��,˚;J+��!zϧN����R^T?�M�35�9�}�ɳz�&�w���d9*{��MW�g2���6�B��w���ۄ��i�k6[˗\�R�9�X/�F�1�vG�7�n����Ճ�P���PRK�p��ٗ��~�r�(J�N��`t��:��N�]T�F���;���k���
�T��2:���o8�f��Voʍ%J��@�x�@�Y~������Ϝ����5)�q�J��g�g�Ⱥp|U��Cw�m���d���p��a��Vu3ГP���\�-�pD��0!>)��wUq��grM.�>�X@����J��+Y����>_�K��M���ƭ><�UP0����£���~�j��<"$U��v��0uz�\x~Q��5N��.��f�-ad��ҡEh���!
P�	PDB�0C�E�A�C���h	�	��ML_=#�8����D%��?���Y%���{�\���t�&@$�M������-f|��X�C���u�Q��{F��;�&���㰦��/�(�@��uC����Y��4R:D��M�]����~�p}t½j�-ʀ��I��r��K���RU�m��܅z.�6H�����i�	�����*�b!�$W�-���_ܗ���R�㖷^�ƒ��y�A�A�f�4�l��;@�v�?.�R��Ss.�%d?�B������.��r2��{\������1j�jA�'�^?�J�s���)����� ���Lɐ�8��'Q��0�(�K�sF��v�L}�S5��w���o��+_w4���O���M�e�?�aR
ȱ��_� �d3z��c����a�����Рڬ�D�����Ӹ�1�t��xf�Q%����=��w�!�it�\��<�B76�o���'�Dn��ܳVa��e��>�4��mF�at�B�b1Z5S% I��>���҇��P�Hd&���+�Bmt]�z[ML΍���X�c�Gͅ_�޹�gfgHj:Nh��;�`��,p`U�D>�*Y-������D�
AE������NYq�:���~�=�ЗoF�!���pWb�k\/�3��F4�v�l�TOh	%��U{������j�\��v$�L��z�=B�7�#�; �`u,��.A��ݰ*���	�0�j5]��T��I?��Up/��2�E���<=�[��9')��	� � yh���3 ��VY��Ysl6@����b��b�@��]�T�� #�a��!4VM�Z'|U�ڟi���,B��D׹�q؅��k��i�s� 5
���+�Z��U�A�v?
�
;z艤�/�"Bd�XW����T,��P�ߊ��oN�?�G(���0I�_h*�y}�|P��B�
�2,
w�L�U/��B��V�e�.�d����Q>@H�ɓ��q0_�{6����!k�e~�Y��)�bE�vR�ۿ׆c ����ք�M��4��+�w$DH�/�8�}�����F�]	�(A6�3R���0���w��ف��+��F���W[���#�JcS�Ͽ<=���@�S��H����$ain�ꭏ�M:.-�E��t��2����A,�Ǚ���c���Ɯ��'��E_V%/��zGc�K5.r�>Y\pP��f�&���!*�X����A������>d����J��������ϳ\A�QG\V��嗵|J���Wg�7�8���[�s����/���)Ui���V2�n|��@׫D/�����Q�/��(��9E�e"��B���4�k��L�Eٝ�Y!��ҬV1�Z�X��ˁ0��ɚ�K�K�O��.bk��/��mØ����ܒ޻]�7�|����j�re����|�?SXz�B�V�*$À̈́y�"�>w�:�c��#�>�nQT��A*�gp �>�y)�l��3� �}X=d�P��l��FN�[>�@v��Si�
H~E�"1�D��k���"���0�	�I�Wd�ܨ �lQU���4^�DL���N��qrf̺Od�5"���g�B*V�rX�c�г�Uj����^m�.Կ��32�	㐵�ʉ���?~�"o(�\�j5�	�����sti7���$4 �DX�5s ѷ\Ť0n�O):g8�!uU��*��D���$	<M��a�ܢ�٦�z�����-��u��8�.$#����~�:E��R��J��c?���~2��W>�r��Z����1���,-&A�q�=�po�ɰQ��D݀�&�]�O
�2p\�z[^�H*���'
�C�&�v���۫�Q,���~�6��-�0�o=�W���Y�}%��b�!F�\(�7���=�D+J؍_[+��s�:�����$֮y+Oዌ`�t�nƏ_�IYw�Xd�ZVO���σ�������Y"p	�u�M^�(*T9���jVת�8�(q���~�;�*qr��b4Z)2�_n��T@Ɍw6�Y�ɻa�V%5='�t�'��	~� \�ZS�O�!���5�4M��u�Г������G��'ci"E�m���Βs�f#>T �w���/_E,��^AK��ߠ|L�cQ��(Ck}�Ӿ)UP��M��H���{�����29�oK\��R����=J�N���';9���nb0�`�fi!�o��n1.�$4p����F����Mo�M�wx�Ӝn�mm?KWA��K�OSs��x�������\���M=�����M� �gy��列$���X\��EV�qZT9�G�b�ެ����ґ��ȶ��=�0E9M�U�dN�%8��J��p�s"\і�wLu�����X=4 ����� ������WPNi>�.)�m�����w+��x��V}�?
%��@����}@=ٯ%f�b3X&]�C4�oӨ���.��O{�*m�������~��q^��r+~	��E5[��U�	�D5~�����Je4�c��3�Zn�h��p�\�V�k��,L�)f���su��-�:-��m��/X�3(3k��&6�8��� ��r9�b���8�VS��y|]������)�1߆	����j/@Ʃ{�*� ����Ӫ��+:Pλ2�� ��<*����g�i"��%r_\�� ^�}�ӭR�w�3��	�i��{P8n���i4<wL�����'���Y�LZ=�͕̽/4(�U9�%�,g���]��Ж���(Ob���H��n�b��@�[}�۴�0-��󬁒���x�Cj�05c�!.�`��jy�=qF�P�ë�		i�K��͖��wK��}��1�R)Uu��*"�b�;��f�̍��&�yC��r0M�̺t���D\L0�P��[(I�i����)w��#�m �UUI����N QsK.���G�A�cc�3D��!�������W"=)�v���������dM]���`K%��J),:�V=�n�v�S2��x�^\��0�iA4;9m�)�F�a[H�}�8U�j�xȣO�+�:���Ίล~�zՄZ05`���kWg�=5vP�hC[A. �m��{_d�DSrjx�:�N��h}̌��\��������9�\����i��to�?���(��Y���f��g�����q��q+�q���B������}6���/�iD��	��$5�$Xs1����8<��|�>��X��������
�$@��,Q��u�	d���ɕ��V*~[/�����{�1X���~���Zr,t�AL7��d_d%���>z�)�s*�%	ۄMa��if� 頷���&�����ų޲� 󄊫t�Y:;��[8�m�z���e����Ϻ��m�lgzG�^��B�wCy�|��0>Ƙ���:e�>�g���]'e\�UyT-���ۛ����Z7�sֳ(�P���I��-�DM��W5�߈�[gm#�� ���J��V��ȵZeA�f�-�� �܄`Wi_@��,2�vМ�F�[��r��{K���w�WCb���@��<�Y�B�f>����_$��Cؠ@��A����8h|�#H�?gE�5��J���`�l����'`�;��{1�w@#��8r8��I�eħʦ��ZV�7�U�w0ky�6�R�O�3n�?N�24����"����)�ł�.k����� �C� hZqoy+?�g>s��j�|�@�~=?đ>_u��O�PC��k~��;֫�]Za��EY�?�ס�\�${G��2{��Z����s�F�:J�~���q���$JH�gA�?x�3��ukI�'��N�Q��?��І���K��l� #-獘Ӯ.�.s�I��ü���ѧ�����i$BC��X��B�Y-���������l�w����!U��f�b���eY>���mN�!�L��6$6�����7��Y�ػ�Tcf���a�d�+��̸:5���&D=a��qwk���f�ZN���^h��:�﹥�� @�R]�`�x�p�ަA;h���Pk���|}���UK* I�K�<�U�Gd�Ru����R���|��z�!=�䩲N�����7+�$4���C�U������[��m�޷��`�6˰۟�\���/Y��FK-*�٧�y���8�1F�Ơ�8e�EA	����i�oB�p���(��i9]��@�f�7�(���=)�G�:�iqʢ��<���6���(���p4��9Z�~֛�E$̒AW��'р?!�S��ԫn6p�Ze.�WGd�>��i}�Gn��a�5��]=��O`9��2uH�_h�Y �(���<3���jK@�����A�O��$=T@�m��)&�W�}:p`)�n���(���j�9�:t��7��E��2��=OIs��5`������x,6`���x	�Фa3#�]>�Z詯&�q,rse���3W��y
���x0����S �(��H��؋�h�����641�1&@w�\<.��p�r?����\Jwzt���ѵ&�� ���-��˙2Wr�"����a���A:D~;v��!�Q@D<f�2n6�ӑS��g�����O�8l�v��Ja�k��5�F֝7�;�\� ���e�T����;��c��"0��� vy^�:d7�*r`���Uy��s���O�)�n������ۧ�D�e�l�I�n�x�c�)N��S>Aה!V%��~ �	5���OW��<�-�rs�7�]�����?w-V�U���t���
�n�3;bt�� ��b�7U��,
���{�	󹔅�
�%�cMd�Ъ3�a��\T������I\z�)�����1�!��o�0�SG�J	��]��.�],����@1���^3S��e��$|T�_B�+ �}�Z,I(f$?�O|zԤy̿S�����f7C�f+X����J�Dk���0�E"3� �_������+,	��,�Jv��Jح���*s���&���lN%Ow�a&��|6�?�yvrls(F�G��t_��c�Z�m����.��U�b�q%`���):�T�4�2��~0�%Ec����lBo�)����V`�ā�^%)jes����>� ��
\�P/���FH���]�'>��Eio�oN�,�'�J����8��B�@����m�HD�4Ͷ�)��`](#r�L�韅fUD���B�n��Fv(��<yW͠t}F)�ʔճ\CD�Sh`��6��E#B󣒁O9&��q.znY���������1f�>OE�� ���N.B{����Yc�D��$����Va�N;$0v�^����5��9Q�_����nA,n�v#���D3��&���/�I��o�I��XgT�Ȫ�綪;A2�lF##��|?/���.Z���R��^����Y�K��\�q���rg��pxD���'<�C��c��5�Rr��/�i"9ꛁ������~R|�D<�*�� ��y��b�MaR
 �X2��Q��n�Փ�e�)����Du�4fg9�C�e�`���6قR=�za5�}XW���R�=���m5m)1��h6_'y�#��˙��R���,�toA ��&��xC��K#H�4��[{N�G�L��l��ܺճsߖ���.�&1Dp��3fa#:����D��� m"�������^p�a2�����r� {~���$�j�U,zI� ����Е����)��� ���.�u=z�$s"�(�3�����7
��>A���mz���,�{� �ԉ�Jl�G/�G9�Ś��B ��q�0�� N��>΍�>XmќDV���C���8�����M=��%>�(�g�]�T�U���ܫ��҈�t�/^�k!_E8A�m�J݇|X�L4�P���:�?���$�(k0��ET�ۋپ>�H�5���-��q�&����Iv|"�ugV�=��l~�����r2���w�<��]�	>����H�1����|�]�H���E��c�"��E�zԞ�ꆖ92F��	�M�SZ֖�p�!eԞ\hnP?s���0^�h�����chx8���:q�o�6�
�p5�>u�5�m�;� �b��$���
��d��_��F���l����IY����HRP�j#�w�Mz��9�{�ZP�_�#p��c���O���~��2.jQl�[��\�ٴ~��A3�+Lꇸ1�{o�Ҧj�#!�����_-9�<x�Qb��%RH�O�B���`�b*H��<nC�a"v���3.�� D�#М���r1m���OO�NV?�Kz*�� �'	��uee���Z�UM��8k"�`�wg��a"o>Nc8n?���8��=�a�@ֆ�
��)cf$a�������s7ˠhuA+R_a4�L9Y'XG�o�U�����=���u��<�����h6H(�HVw��p������h2�y�{�TIMtvh����Z
�P�N�g2�|��%��7�6�ښ��l*c��y���`^�<���J��� v��\%#W��J6�N׭s��_��"!��M�Z`�g^��Rv�֘(���v�3J�Q9x��ޅEK�n��՘p���@
+���a��"PP(��! �fYaO��:9�ߦ9CIQ茎_�~*%t�9�  5��l��k9dv�{�Q� �о����o����Wл"�OD���E��,�h�B�k7U�~٦?��n�wl;��1A���� _�n�Z�?�b#m]�I=��j��߃GQL������rk�1�bU�x�7���s�2�h�)&������n�KC%�l{�x�!9s�~�2��ի��ʄ�B;�<���RY��m��\�[Q��)������.c@��k>o7�}���[��>��׉�c�6����t�( ���|&��vW0�.�9Zd��Ap�/���鉸�W�%��ly6jK��Jcg���آ���6�W����ֻ���<m�y�h�#x��t[���3dY��g�C=�D�9���\R�3������M/��ҁ��v��������̄���Q6F�T-<_����~���l�Á!����~�L��ıv��[�3f�T����X���u�ޭлg��E�Fmg�Œ��Xc*�.����5�Bk;��[�b�5xi��:�@^��w�T����_���򡔊h=��
�0�i�`FAQ�sQ[`U�-֦W�M��?d�Վ$F�b��s=O���2edʸ�\zR7�^&?ò� ��ܼ.B� �;���Ο|3�ظ�19�,�7t<�C���fr�r0s:p�_:��'�����lzu�A8~.��%�:���~�Z��!��3G��EbB��\�4K�Z��<Z�A��+�㪙���.�����N?$�c%�*�{�M#��3��,�X��y����g��w��*� �!J?��SnS���@H��Ο�@1<� �2��*ȿL��Y* Y|�P���p�G��IR��g8]cb���M �a�R��O��LJ�%�yx��\��A�Y}F� ��� �ƽ�.*�5��I��D�M����ʟ�MZ�=��Ԁxv,Uv(<��n���S�k��[�S�v8�L}QRT8�%��b�4�سW��/��_� 8�N&�C�P���N\=�D/L�н"�n���!/$�r^�~��p�
5А���?3�tv��g��>2С�*�C�K	�E�E�<y���y��:��]e�VYs�;C���k���
��e�9�������h�kt�T�U��e��	���6�|��A�o�S��Tc�0$`i_�����mC\COƻ��M������/���h�5�7�-AE��O�,^FP��B��(I%N� ��X�ч��9_:�F�	������-�~�SX)�>L�ͦWx�v�ݥ�:#1'}�D:�����4�ߡ����S�`����[�#ТY����[Tؽ���V�+�f��u�j���yv
��*LT}w&'��^��f��h��g�D��w��#����E��j�k0�`2�����Z>K�:�F����/��X���ro�|�8y�/����C�|:�G*�k����k��잒\�kd�C-�m�h-�D͉��2dw.PE�4�����T��Ԛ��N��&��(F�?5Ik襢�z�b|��-�A�W'k����R�S����GX�����2 K<P��jH�a"��~W��o�kHn~��:7Jj'�4,PdV�)����~�e�-��UU��c����[1��a)�1�2"�f2�2����2F[*P�G�AKEt j�9(R��\�����_s#����Ft�v�Q���ң&xTD�S���[�^^�3c.�r.s�Ʀt�Ac�����M>��f��%�$|�R�LN�_a$�FX������*���I<�^d�cؾ���u����-���ݜ�JT�ŗ�s��Z�7In�¹�,p�4�u=�v׆{�dzk��
,}����_�0��"B����-�jS���4޾�Q���&)ܜ�`�'��x����k�͡�Q�Jߛ�WmT 7��V&X|��u<�6�y�j-h�i�(� _,z8x��4Tϧ�	�ʝR�%���>���+��'����T�oU������S�F�A���4	vf�%�=��
X߬����
=,\�#&�XMЙ8�g����J��?l�ݽ�|��w�}��YΉ��b��Un;D��k9�g��t5b��w9���Z���$��q�Qs�-JX�$�iA!H��U]:zdqf"�ۛr�S�"�6bBJ�⡇���W�j�0�o�
e�����нs�c�@��ի^-'��vM#��K˼���]�h*�:�B_a�[����X�X����Φ�	�q� f,s\$ن�+1��YN8M�(k�h~��Uߘ�� UC�JRT���22`֝�4��&-�n�1�T���!���E=���2'�@���)��׿0��=R��4d�q�e;��c]b�y֓s�\o��_r��b��=L������1�,4��[Zh*���Y����|%��ԁ�C �����s�,R�>y!��K�/;�K�?�ه1vS�������(\�n��'�+h)�p!PhE�bM%�՜���v9#� i3���@!�XWu4����o��L���>�S����m#t���U	ԋ�
r�-ع>����IU�	v���5X�6��nD��mP����z��(�y~�Z9���� w��.:DL�H�-Y��WQ�>7���jEc��M�I0���S'��E��Ȼ���Q^A�`r�\�i
g��z��� Y�ޒ����*h^��2��|a�Qi� `Y��<*@(�H�m�9���&�,�ٓl�������9�-��'_��q�[#-SEs;����Hy�;h)˓"*L�΅#��A:"U�_�Cr�5n$��Ml�B� ʅ{{D���KPb�t���|�6K3],�Dx���k3hk>'07�`�C�Qֱ��Z'6�$Ev{�Q��T�V����G�~>��D�<�<&�T]����G�}����?�y �{�ُ���� Ol��f���F��;������'��b�R1K�@NJ�U�؟�n忾���Zyo 5{1M,k9�����:J�X�>T�T�h"8��q]��0��<�֛&t�sx>�1Y��}6^�;R���8Vu]�B�7�|$K�/���c��T!��Ǝ�����f�u0L��fȃ��LGZjK��_~ �B��3��x�"3��l��N�=�[�?EkCA�S��,L8<�:')ξ�̩@�!�gi*�gh�ג�x H`�#H�($�%�%K0�mzL�Z�B`sLW���X�~���z+�p%R�G׋b4-��![��ʕ�$��-��tӣ�H�l�~�rH���2L�UѸ�,����~�ي���uC�R���0X=@	鏴۩�`�?|��[�Ɉ�3=�WJ��^�O;YAs�Q[U�$��M�v�n����~�y}���!���qw�v��;�sr�u����f�-bjh�"s6L_FC��N�	�����k��F[tb塗��x������3��	�8�yZ�ܭȖ��feT�KZ%*NrDF*'B����*�`o�k��'�[��#v��ϑ)6��)��P�s�؉�^�8B@�ɤ��h"H����gBknnR�mi��<ԕQ$�d�Z�P�6�Q�H�	�0�0��z"���}V����*݌��b�w����9`��N� o�] ^Z����lt"f_z�2�3�:�m'q���<�&��f��+�>MCeJ��<P���Eda�� /����������{�@6;���a���	�)v|���-�]�����D�3ɿ�k5Q�������Ix�B�Z���l�R2��9c���4=��lc�n����W�OI����
G����-��$������,��궾j3Wvx���\m5NQ���`{��˦�JrHH���������4���xK���Z�M��u�ׄ�%�@���ͺO��2�V&}��!_
����v*�4���3��}&�����;��~�'�\��syruz��nU*TG�SW7!h��h��">���Z�l�,Q�^��Ư��!JuF��[}�y,����KgЧ��~0e�������SNZ�~<�E@t�c�	�X�$�q�z6�t#{�ج�Y(�;� ���t���i27_�4�a��b��_�ȀN˻H#n����wh"i8�Z������W7�h�fU�?Pj?��'�Ή������F�=�{O/�6QbT���*
��UBh�Nc����Y_ YW�5����q�qG�|�w+�8�;��W�_���A&� Pp�P�����(��l��g�:Q��#i���V��"/x�ߡ�=�f�7�Ln���(�I�qZ�0R�>z+)�7I?��r;D�a��$e��b?�������!��d�.]o:Z�wҷ7���g�h�Ow�_/ߴ�`�����%���g�1s�A��#�����5�8i���.���W��k�k�x���\�P���j��}a���T��S	���g{�zo\�}�yr�B7��G�� ���}�h��f�E�a�{����搷#Vڟ��;4��8`Nvo����y^ǉ�d5;G��w���k*���z <C����b��(lJ��pѧ �ދr�i��[zJ�@�����KY�OB)�+�A~�~.c��􏔺z�Ԑ�?a�+M
��,��vC�}�TN�H�AQ����Z�-cIf�C���/�V:@�w����c2�q)QlYҦ�����l�"�� jL�^Z��J���+� ��YBϪN�R�n6�L�Lʪ��J�g#��qA�9໮D�#����lA�_I�%Ƅ,ь�T�S����͏-�<R�YA6����v�|d����r��ȬB�܈��%w�ݩ���C�
9���P^����'�B��:XW^�n��=�Z$���K�]��LQ��}��*���o/C��3$V�!���~��9�9׾��/�u7���/yCM�S��_�_�0�S'��F��yo�S�F��HZmg/���u?��a�:0߃g��d��pVZcR�Brq�U.�����g�g��!�q���k��#8⑅�V�}�f�6�WV��u�!\��������I�d��;�^��r�;4��i��l���y		��/�H�u�֓G΋]��6��Z�\�;j��TrSB�/W�)! s�ڍ髌��ZZ���4~�)�7и>nX�g'K������T�0j3����딧������xNn���������@��&ڒ��J<�'"L�Ym�C�q�k�m8�	�����Xoz&��XӉ�(���-���Wj|�ST,m��PZx�t'W��U֩.��������k�W����6��ړR�P�zsp"��m�|��l]�!�f�<P'�RXI�:ֹ|̱���z%��S��*��U�;�<}�1h�$=ފ����ߚ�I��-�*�hե��n�:���~z���I�	�+�U۷��i��\�G!���M�S��|Ĳq[#��P�8�1��}��8	�V�p�o	�1���TRu˥���*�,��B��H����g��[��Ț�˻,͍l}:�w �,
k�n�X��fȻ{'��;������x��RM �����z��*J�0w� /چ�̰�ō��]z	0��(q	夾O�e h�l�sNq����_2^��DRX�8��w�	?g0�|��jd���Igr��Zӱb?
�dx�e~3��L���Y����E�`�p�3,g:ҽc&���ԗ��Ȧ���m��&,��j�V��tyϴ�(/�������fѲ[�`�ȇo�6��0� �����ԓ"�ٺ�Mm�!z0��j�����\*a�YH>D�k�R9wU���1@E��@jz�`�J6��ьc$]�� >�F��@�m�����fhyM�cKg�L��~g������M�π"�hc��ˈ��b��9�*�c��F�{���+��Z�7�+�6�X�D����*��{,͒��l�w��%�瘁SQ ���CY�(i�Dw� /Yh�P��^�t��Õ��I��C���ƿ��ރH3�.id�O�M��9�JG�D��n��,����]`d>a�.q�ӧQ�m��f�3T�ב��\�VĪ��\�Z�Ha�5���w�q��KZ5ha���(�'%Ţ�u�/��;�� 
@��&A"׀i�|���?ha��}ݎ��N����c��zg�r�Pߝu�sUT�Ya��Q<.�B�;6��"�^|���f`���|ow�jxh
�<�2�q#i����pYE�(���s�)�'}v0�A�k�NǓ�=+x2Ѩ��3�8G�9 L�\G>Ր�t)�T25�&�iH>�}b-";��%���)��Wz榭2�c\�����P�Ձ'�������Kq���x���������3kn��CH���v�G��z8����s}����N� o��=g2fj�)��['ƍ�z��ֳ�3Z@y����}h�t[o3��>��-p]p�z�CJTH�*��] ��xv���{��v(���ִ4*#T3�oO�aI���P$BثP@��)��u\�v��+h�So��Ӝ%a7�B	�Xis2�a��&Jw���)#�5��sW��y\ܩ����ɛf�ɴ�,��z�p>�j��[���LYg�'�������H�ph*���K��,�&�b!� �1�)%1��x�Y�8dO�X�p$�%�1#Y��yWt%+r������	ONXu�ĸ֝c�^��S�2�����hL ?I���KU�"�Y�o>��?XmQ��<g�oI͛D~/\�Rm��YTxݤ�XK����:� w�F�J5��Dc&P����Ο�y�8)���nnX7Y]}�{�'N%#ԝZ��v�+� 4�(T�*��5��4��_Zw��o�[����|��g����wN�ा���S�NGd�M��ӣ��9<��m�K�7/M�=�N�1���gU�
P���(�q�S��Y���{$�{"\ X�q��$���5ĸ�@�!�카i��-�����oʇj���*z�n�����f[)w�X2�����T��������iF�����N{ϖ��iS-
�@�!��F�2�$��)�>y�xx�Ӝ�"T����mvH��V ΋�o���a�_	�L �I�)�E'����OW���O�i�iȬr������_��{��;3�����(�{�F7I��e.(�죃�N?��#� ��f���j�[F�z�����g���,Ofn��r��Kɴ���F���.�J	���-��Uh/�j`m��ߑ��:��bD�\�U+=	��8}��{�&�:��BA�:_����d�NU���f�e�,4	(�"&�H����d:�)�a�v�c	�o�T�W2�Ș�?P<���
��<� �T�$̺K��1��ߨ�5
=%���[7I�)k��I_���@aY��<�m#B��:G��& ȉ�+o��9�T�`��Dξ,�;����7���q�%�z58�s��������^�9���יXX*�L�V�G_��i[�)ķnҡ5�tR$���}yn>��@�ot�z����TL�`�j��՜��QM�8��1Ow�?oA��������̯��p�h��#�h���T������*��'q�39�F�~ζ���8��yw�M�ܘ�)��1�`�l0��� ����b���<Y$��h"�hU�ku��.3mue% �ħQi�H9����Y&���p'���BC�ّ���`0�oBV>bN��6��p����:�.1\Ýl3��)�k�fU ͍��*m��2�`��_`�V1�ӑ�O�*
&�>܀A��4<1ׅ'�'�Q�{�0�,1B^1S'��k.� ��T�t�)	��Į �����h��!>��Mk�j�)���1Ҙ��M�h�+�"��2Z�� ��_8�*G�j[��^�)c�Z��ۚ�!��Q�Sb�͍��u�A��ļ2�[������t���'������Z���ڽ5���&�l��	v�b$+(�],&h9w/����`���T��b���03eM""��}S���Un�N�H��üI3hn�A#�t�Bo�۫�x1���L�����V�O��<;v�b���!�|2���4[b�$���5�HsX��n:_���=�b��v^�[��k�M���j���G�3�s&\�
���'�-s����/vv�E21�œȈ d��/���3����|�I�̼�{CO1��ӍUe{�rՎ��0���z9�!�_�s��pە1��A�\�6k9��K�d$`f���� 5H�2+Hn(�HN�BPχr���`�Ԭ�*��):�9�q�2����݇��7�o4?�K",�gvFF��0��S+�ɻ����⻎��l~k &��	4U�o*�(Q�/��Z�N:�[zv�O�Θ��v���=ݹwn���Y8-Q�|R�y�Y�|�t	��}��<Ų�9B#A�~(P�>���51M��^���	���԰��'jDbh0פ/_\�w�|��lh�uK�"4��L�[���$��*���@M�8?;pg�}���yL�P1D�3�K��0s�D+�*�8]j�=�q55鱔�k����FSz·�����]�J�h��iU� �5O�q/��o\3]��N�>���w�qY�bF7�J����& �*�g�0���8��� L�|�b:4�#w-ܝ-k�pv�o�f��P�	��˟J���8��uS?R�lI���GS��gU��)I/<��,F����s�It�Y$ ��
s�rc4�"[֗�����K�f5��,a����q��ǽ��op��%ZVt��	jM���<'aӼP-9Ba�=�/�V{qr�1s��em�lس��twb� �@M�#ͧ����������_�Z*Z(ƽn�^�1���)��~m��E��XGx�>E���K���aWC��)�zG�Y��#ɚ3l]~����T��Ud�>>��E��<	��o�B����}�\Mv�������#=5ߦUK0V!������Q��{�u���_M�L�%y�#YI��"��������n��	�`�8 p��S���[�,�SS!���̽qQ���&��)h$R�0�*?em�R���4��}�V��W��m��H�YB�����h�*c�ì���f�� 
Q�q,��-����v��=�[U�*>^��(�� *���(*y����rEт��K���8���e�s� ���(���/��n^���'5&ⳣ�_Cw���ʅk�\xD��"@�-�v��k���T哜��E�*��^��-p� �	gh��YA��)��}�"N�QޥK=���S@���B6$r����k$`�5������˳E���Z�d�-������J�����q���j@�P%�+��1��]�hz����U��`���!�4~�F�1.n�6%�.�zu�1�n3]KF
�������і� L~ LAy?�d4�q�R�bA)������n���SB6�p<��R�J�9S9���N���ç]>E�qWa$C�Z�"B�;Yyݙ Їc��d~tO�
����L;�70��#���t�|4��p�'�F?:�Q*� b`�`��~�.aMI�h^�7��ZBR���)�&�9��M�	��<���8� 	���)��������O�3$6_��.��#L�,G8Z��W��s�m��]���B�ZL�����s�l�����im7_�k�^+��Xƌ>���w-:�a��a��Ѫ��� !â	U���R�ܒڼ�$���b���,%[�'W�7�j@��йRj���㐁�j�c Elx�'#Zc���yU��텭�d+6a6�Q��@8��"�Šz�}��f-��N�l�D�d���H�Ls��dCN�uF�A<ό3�$ �C���6H�s��M�,�e¡ 7��Bn_���y՘�go����氠���\ ��� S��L�׷��ڏ���{q��j�\K��m˹R��ү%WL���c������Zy���0�8Ji�Y�胟l���
���l�U�
���&�h��I�������!��Y��`�esu�F-W��G����(����**�cA�M��+՝��i�e���#/`�Uߒ,[o�$Oj���B�����;J t���7!����NV@���^IlƤ�Q0,�^vm�32�a�<J�Pm�jn��sg3�)bQ�$ꇙ;#��im/B�w���K���!Z��R���u��H|"�v��傘|W~ٕa5wr����B`<�t��x�v���ŧǘ~)����#�n�ƇaG��Ps�rڈD\� ��I�ID�K�8�wz;w���˷�J ����l�g�rt���H?��^�yMc,�ޅ�2�3VyP�U���F�_�ʊ��{�d���T�F�h��|+�u$Ӓ�	P��\%VU<+�Xdl	��3?��p5�Mu�O'�z��W�/u���E]�0><��=j��E�wIN����p�S�`�S��Vhw=-&C6hWA���\x���7��A&�� _�8�pm��#��`NT�58�p>r�nκ��8S��|yj��F�
��u@x�x�����(�{���?s�{�����S���q��A�����K�VT^`o�:(qJy�q8�gt
����]�]nF�<d�̧7gI8a��Q���=�_n#�P�T|xM�~広�ɮ�PsA�o.*E���?��Ԅ\��ʉ�wФ������{�7]	��M����Y
Ͼ+�?D��gĽYm2f+!�4�������R���~��"�wcZa9�m/|��S�'?{��4mvu�%u�&��9��&|x��1��xڊ�E���g�+[�B����X�W�H���/�F�p���%��P�f��
ʿ ��e��c�����L�M*+�*f����6V'��O���[���C�P!�[��D�����a]����GRPROגנs;�-���`V��Dd ��#������e��R?[T��`Ӎ]��[�+1�B#�!$s��o�������`�,l8�)�n^�������%V�/�0� BL��V��f�]��p���s�;ƪC~� |a�VȈ2�P���~vpR�
��i�� �=V��s>վ�X�ټ�^�.�J�(ƅW6|9$�޻���ρל��cN�wSFa��׳Z�R�(�k�?�S�~P��_k��i�WS��L�q�K��sN�����;q������M�a{��Cy��s��H���!=���Ҡר��ʋ/�:1�!U�K�j��8�����J�uBz��-�a/](@޴A��ݽY;���SҰ�����A��2
->������~�[
6��7χ������;+X�RF�K�yI�<� �@c�>�/�&3.K��R��`����z*��D��r����HM��9靧UsZ5']E�=~���6��ε��e��jo`E߅8�L6����zX�0rj����?���=>ɽ7�������7�/S8rXL����/�S3@FBOǎW��M�H�M0�4����6�7�P�+TmX�KFSVȆ��=��ZA��EhX\r���X�)�,MJ`�����Aw��Gx�;ت
=��
̬~�|����n=jk�p���]z9Z�	����0��?��h���_+��UKR��N_��Q�3h�˪��O�e�AOUv|�=��3�Ԫ�b9��L�1�kԉu<�kً��N�EߊS�W{���Nr*:��[fX�8�����m��Z.u��~�/.�c��xt�\W[~��Pc%����(BV6Iu�څJ	a�VE�zy��x�$�E9��J����%����<��{�ۺ�rզ�%�l��7>
C-i�{j��"(�G��Xd��	��~@o�$�h�I�po~f#����)����B���W˂��I�:��+�Ɠw3(�d�"bg�Rǳ�d�pyo��U��g>��в?[v1�'a�s��j=CfE�b��ut���~��j���u4��|h�H����A17*����<�է�K4�n��BM����{@���v��ttk�dm��@<
6�T/+ч��:gs��	_�IG�uN�8,����W)�ȹ43�2�L�%�0��('�-�2��Y���r0�6]��a�
Ml8׶��z�(���� Dș,��L(�"ףj�1�WC��az��`&�'!������a�L��,D�ϖ�PX/�P��m��u9��!�^�2����tOȃO?�Xa�����h`s+޶l��WX�<Y����P��cL�
�Zzq������s��2��ţ���ୌT�:��b���@�*����Hh鰃�͒��6�gƤ�q���8��dC�Όn(��%�R^t���m$`<�D!\�H.݂Ǻ&gs^J������Q-�	t�+�`5t��:;����U���W�4m/�nS�6�'�uq��m��{s*"�,��UrB}v���~���Mm�(����x�Ϻ`��wh�7��C��[��f����rLƶ�U�6a�'D'�R�T��չ'f�a�����>��J�H`�(yF�z��D�9hY�fa5�*'��*�)̤I&q��#�K�s,�@��0'����"bn{k��6��̑���>��׭.��g9�`�P�C��h{����(��؜d��IYc	ٱjD�kԆ�=�Cc0�{q�fDY�[��J�~Q�.�/z�-4>u�{��)՛�xM��������Oi]��Y�4 �3�bh����ؔ�8���Dᆉ4��<T[|e���飌��ȥl!�X�	����ͷ��U_Vr���׎w������;6��|�i��X���;ɢ5F�y�pR�N;Ӱ��NE��n����<���">?�u��(W���	���p�0&��49�K�S��)bN>�.��C��4\���C	���ؽ�y�]��P�Oz%�\��e.� T�9O9d6�����n������)USe�h�'�J�0�N����w��cf��8%:�y/���X�`�'8����2�ZY��ʕjUP�+��2=�СY靆�Q�������b�G_�<t�ַj�J~wޑc�8�{���Y��f蛡�ɉH�v�Ӱг�0=�@eS.����<�n~֘�ǯ�4Fb2_1�x�>|�v�Rʤʏ��Z�L�1텀N/��'��lXz$�
}�~�ƈM�R�_�{J�UCU䡘҄OۉsM�[�6t�M��K�f���+܏�jN8$��-������~�E8�6���3sbʹ�@i����x�"��K��^���&���v�VO&����~��3n��1W��R�gI�)G���-p'�	�W�xd�F��.4)��ҽ	�ې��	�Iт��c�O|q9�ӽ|�����\AF
F�	8u޶G5������Y���e<0��y^IKw\�1��@�R�'S2�p3�\��r&p<�7�)O�ӆ:r"]~���8[	<o��E��
����w�u�R��uC<N���S0{���74�A�_�����I�d̂L�6#���y�^����/�$�׉��(�}++��,�������$߰hb��_��R���������Y���>�h�̌�`}L��t[|
ɳD��&�l�q�q�E�k9���*@s,�f�w,t��7'�'Z���ֻ5Yb�� I��>c2,���m�&��u�mf[J�����I֨#��A��x;^6^O�b�<�c{�P�5��I;{?��M�Z���ɐ�2~`8u֪���t��%�׉5*]��v���%w���K������\��|T����3�}*w�������tlpq׆�
� ü}��r�Ђ��T���3M�B��M,��)�JD�G��σ���n�\�������@0տ��J!F�v��#4�;?������T�*ŋ ?&tSV �X�v�vFiU/��z�;|�;�����"iB����EYM�c*�g���tmW��#�>�Lx���v�J{���s諮id�Ï�I��A��UL~Q�Q���Q(eю�{���=�{��{�|���b^�`�1��xh����6w�;r�~+����L�_��!�߼�"����R:�hB�^r�|^&d�&����hJ�y����"�jucm7z��p��U4�E4�I�5�����n�a���ǫeE�q#u��+�&���Q���H@��u�$>�\�/Yٞ	�Y>�i*?��N�꛶&�Lx�~ ��0�#�	��Q���.l��F��%��i��ہ瘾��Ƽ�M��@�Q"S���*rFyQ:�x=�і�,��c�LH>?tp�,�,�K�)}����ra���2�����:�;����8���r�S)9?Oq�}�����A1L�]D9�K�/x��B1\?^"2�`�T�4^�E!&�]e�C$W�n�s8��
_["$%=�$������b��#L?7�q�z��o�:�$����x|��`�J�9-��&-¯���YKS�|�샫��o\Ǵsl���z��>w9�N�a|w��ϕ������x��-�����Y��ޓ=�)C��Cئ���eZ9��\��<���EH�K;�YL�����pEߍ�"����p4��|�a"}L��(r��W� K���޻�u&$�.���	�!R������� �X�)6�2c���p�uߜ'/[����S�&hu�� �E������D�	+tb}$z�N&�@�����(����8�����?�N�2'��Gĥ��HawI;,��k����baP�зmD�yG�1�|ay5K�^De;��	Uo�L�'���{/��oI����<lY�9�~,��on��Q0���R�����y|E:�)��������N��#Z�3�.'K�@\��.
|[ �򓳊Bh���.��{8�>o&�ǬжaR`%𼗔,��8t CPI�@���p��`�q�'E���	-��|���j{.0���Z��X5\��,�r�U�&���L�HT}� �F��xx)w����y����s�"����F��ρ���6�Cbi���'h�G5�-C���N\ym�����F��������|�:�M��P�[6$�lsI�z7�y�D]Qb:�G���&R��*Ir���ߢ����6�Q��8ś��m�I������s�h���@Ohp*�K5-3n<���n檱n9�����oW\���pf^O�f��fl�v��#śRf�0VF��	���Սf�U�B=���#�NI��}���t�1�\*�o�����&\�֦j�X���&�L!�V'��+\�4�T�͝<=�+�f���������V��ў��0�����o~@צJb��f���Zsѳ���c���L�:����.H�	��rB+3�a�(n^�,���DL�YS)�F	ʃ��>�D�	���f�H?�O�=/��6�T[W`�%F[,:u���۹�`u��\b�b��eq-���'�,Uq3�P�q�b����hq_�x6��ޞ��Y��K��Z��mM:�(�|r�&��`�5���)�ӬTv/ODܥ�#�]���ˉ9���R$�ѷԣ�M��n՝�����-�i�W��xN
�h���;��N>75��oXe�U�aQ5�I{�L��dS���{�D�	M�~�hͧ6L�zd<mU暁��TP�L@J0SM*(���u���K�>����f���zfX���	�ꉖ���H��w�9y
���+zt�w�ƶ�Oid8���\$}C�U���q�Ȝ$DS�kp�Kq��[�>Gov�lP�rb=�\K��d��(i�������*_h�vLڦ}:�%h��~6�ObvĮ�Q�L��X��4q��a��j��ɵ�ft�{���V����h	��"�;v})V9i��A�Sg�P�����@^�U'�0��HɊ?�l�t���q����l�U��oW�tΜ�A=��~U��S���*�@�[.Y��|�d�dOJ����`G(�3>��d�m!l�W�B�p��bF�!̞����v��'�o�N�C����E9c�z��Y�K`J!��uF򓜷�dedxΗ�F7Ķ_��v�����$�L��&Z;.p�����D&{���"�����_3����!g-F{ G������m��[s ��p��.C�}������C�m^���R��d<��0�m�@a�!��t���s�Az��;�%�]>�2����Σ�1,���K'��zXG��37킬�V ���'xa��ӵ��,t���T���l����'ח%�Z���-p�H���%�y{����2�5���F!�>9}:UAw�8���t��0Uޠ�u�}�֞:m����7��Gx"�Z�T�^�!/M3�� /<�װ��e�1ޭaeI(�}b��tB�(`��;����W�!"�:�o'_;����[f�k�������I�a#f�.G.�[Aj�ui鏕 vh��ĶV
<���"�D���NSAj����<�+[����|�%#ʒ�!>r:��'�Z�����	�����7�7��\�i5�3-0}$��w��Z������:!CN����z��tSA��7u��Tqb��^A���4MY�%e�q�e��;�Sb�?p
�B�e�Uw��-�v C�n�q����C��i��	ᆩ�i�V�� �y��#|)�ZN�<��f�rh�ȧ�tH��M��NH���E��Ί�e��0��	��7��8�w'�_��A2�ZD��(��m�{km�FϾ��1i��y��M?�}����:��7ُ�:0iSi/�����vT�kN���3�<��[dqBF҇��2by����-[M�B׬*Y�*`Z� r�{,ﮆ�e�1���Ts��Ya:}�#�m�?�����d{�Vv�t{Ȇ�O��U/WA���${T��2[��h�{>���t��% ���������n����\,L/�����-m�N-�N�ㄤW�B{��u^M$�{T�[��u+y9�R$%p����r;��?�_�XS>�d&7d9���s�^��X!�7��d���k�m�T?h���$B���q�Xg���Ts.Z�x=?HyV[�Z�L���[�x�8���P��q��.ւ���BW�/��H���/�$kY�*���[���a���cs�������pw�)?!y���`����U`bl�N����V�k|��)<o`[~���«ѹ�"��Μߍy�����VsY-�1(�=Q����Ȋ��87rf�g<�Vţ��K�6o������eTf�F&��G7�}*���3��?#�/��Y�\��Ƒ�.r@�/p�Q^��K�+��2�Ƙ@��&�֏4e�k��a&�	�b��<z�27�w������QS0��k����1�f�8'cc�z����h=��RZ�l{�sE����'BO�<z�K���Cr�s/,�~�a�H������V�Ʋgl�n�����o@��	�hۣz����;{�W�?�c��ui=��%�j�eɖ4��'^9�?^
.g���Qnq������䐖/�2cRa�w�b�m��mN`����&�5�$��{���g70˚�����Le��~Qa86�;�U�0b�/�B|��P�y�G�mb�sz���j�*��Z�3����ނt>s����e���DGt���o������ҏ�0�G��(_�V~Ɠ�5�>x_1E�	���E��}�YY���ɉ���-�l[珣�P�-Y���-���]�`�������Ф�b���������+�Y�v�VU\���蹧'��X��8��f��ב�uR Զ��-�y�ʳтjs!���R�G�ywP��6Rz��Q�.L}�C@�M@����dz�y���&tp�:�k���%�C�v�_�BK-�ڙ��~a��a5-k���+��⺺�:m�����_B�d�����h �����z�8�BףNYiE[T��%�{�jZ�ix,��	T����"���W��1�1� �+a9f&����4�)12�"=��ظ�X��� F��-!��8d+{2��@�~��{��q��5K�ׯ'H��T��F�+U����Č;\�3a�?��Q��.��+d���O��D3_�j�@�2��X#���Cz���HC s�3=�.�?�%)��������M�]YI�k5�׾���WH���h�o�b=�-��� � �΃��������y6s3�W�^C[QfOq�<]���A�o�>���+߭/��p��19����"Ǎ�h00�	۾:&ژ!N�\d�Ypd���8̸~��F0 �����||���5�ڏ��E$ P��^x1�G�[�x�L��a�WeTҥ����$�d|4'S��դyyI �#�~Ըm��L���G�I@�݆��]1A"�w�O9��k���1Y����Hh8��RJU���1��"�=�,Qm	x�s�*�2����i��ݭqKo}�Z��O�Z�9��_5�G��o�3'=�� 
<�c����=��� �˚�����Coxk��E�~�F���S�˟�^ X%�	�"���8~��߰	y(!J휿��UV�G�eg��p�Z�#�Ϋ��>�h�:�	�2�¶��� �}LDK0wt⬚D���h�-C�d���@��k$"�����$T�1>�,v�$�	��]�&�3���JcdĢ�ä-��bO�J����Ϫ�	lcFk���ڜ��6�pW��Eٛ���Q|�+n( �E`�m�[�c:��x�X�r��ߒ�a�SUh��/Q�͜�|��r����ξ1�2١�\�<���F,�;��~�^H|�D��#>m��H�Cݣf�q�D7rzES���m�ZL��JQ��+5a&�3���PЗ�'�]�/�ITo��W)��B ��M�&-��`�)f#�ξi��Vgλ!�:�x��#^�T4%t�5+܃v�3|�$�맞��'Ad���To�Z�̿�}Z�e��@u,T�Sc̄���6�!�I��V��#.��1�Ϣ��ih�ִ�O��j�1;�d���@��*�!߱U����BD���x�2kY�������Q�����fm�E_*)%�>K܈ ��T���ӂמ+S{)�6�2֥x�t�Es�h�D^�H�6�c3>�N1\��w�G0��:7�9��B��HФ���.�H���J��:�t���õd���
p~�;�G�PN��v0�y�ꯟ��@t��_[#У�H:p;g"�6a����p�R��]ײ?9����`��:��^��&�J�I8~�D��?9����:�H(�4w3=�����$8K8���Շ���:z��vs�6oM�����K�����
|pCJE�9�h�C�ɱz�s5%r͇��:f��a�N&�yWPB�~�C�%b���Z���`C���%3���5�!��Nme�w�Ą�A�H�ޓ>��Y-fj�Y{��e!�8\R�ͺQh޴EUg'%9�;�k��Sd��Ȓ�[|�^��(k�|շb���EB)QG�m�z_!�&c6m�0.��	6�=��420�w�~������ܱ`q{\�v�+�������럚�d�~S��?�����?�W��L����$��� "A/tw����!w	^��|M�nvJv�̈��2Y� �6` ������
%�eWV3>M�3�l�>\�Zp�rx2����J"G��fԧa!kI#�s�_�d8����KEM�W�8�s�lA��Xq������y"�fmlU �È�H�H�;)������DB�E�?�����G0��6�\�z�-��b1k�>g��!XΩȨ��Mvfj�b�f�t�Z��88�g3�&��,�r5��>�;��~��l��Rľv���v`"�xv?�;TS-	�q;h|$�B[���l�f�e嫸��C��8��2l��qo��^�HlIwz���_I�3����BY��%n��w{���0r�؃��������[T��2��0�1��a9�XP˙�+�k15��"�(0��g�QZP�[ĥ��_m�Z�	��� z4ʈ��S>l7�N�\��0y3*��"��op�x���~'QO��G�zdT���QuR�����dU��ؓ��P�~V�I�m￉?���h%�H��`{|��.��-
��դ2�ʉ@��A�t��3U����_�6R5��jt�Y��6��î:Qp�E����y��d��Z>�RO�?�a�B��^`�27�V�i�%�HU�bP���*��y
4�
��	���)�Meg�+�������D`���ZG����C������:x��\>f��CՈh����CHb}I��ב^�#�A���ce��6�����;��g��Y����N�����F�E&�f��4kR���nK�=$��䕔y׊Ȝ˞A��ߢ�Y�o�ӵ�[����ſEy�;�bY4��%ݽ�P�ͮ]�^�����n�P˹�
�l���@�gᏧΐ���<�Phh�������j/͡���ݮ{%>W�ٳU�@�������� q���
�J�.�Hd��@F�x��X�Q�I��4���I.pw:��؍��j8���b��{���\H��������Y��]�5��V͢h����R��}�"Npήy(��L
�l(��ȳ�k4`XO �÷l�I@)+�L�ۂ;|�P�<��e��h&�I����GÀ��fX���4v�PJl糖�QLү+��ʏ��M��:iX�i$h��\e�Ttl6�+}K��h�5s5"?��%S�����j��l<��c$i6m������Id��j��N|Q5�a��t�D�mҼ�"����EF`&M�z����3@i���Aͽ��ߥ��I�>����KRNs� ��@P�ߦ�fS7��|��z�}��s@�3��e ���F��df�^
)��I^v�d�xVMvb��1�8	&�L����������Nz`�f�5��UH=�$bd�&Sj����'mڛaz�9V� >��uD���}���-[���������p��g` c�+�H�c`}���!ϙϣ"��q%��B⼵B,k����Q������;�g��P=�����z���b?��Q�VSXZ�����p�(YK����Ō���(������Ά3��xkcc"h+�7���z���C%�z��5�4�a���b�%��o{��&��#~R���A ^ ��®�a�����ª���o_XJ~Mr
�t��'���Y��'v4�n��Dӻi>�[�f�wjDĘ�ع�T驮��j���Q^�bߟwzȔ����R���$#r�4�>�hC{�]C�t1������vq�p��*R����c.)|x����U;��$�:��o]5vu���V��A�j���j�,w�U���J�2 b#R��˫9�̽�q�	0e4�oo��#����1J�9��:������4�1�����C*�!r*;+ջ�����Z�w��nߜ���7I++(7���w�� �,�b�[��04�s�q�1l�O�M�����g�M���~�L�<�=4�-��b/Ħ0H��*�y"����n��>���������������0�K��ȧG��1N�m�Uw��q�e2 m�7?ӀZ[�̙�O�ȴs;�����/���Q�O
F��(�¯�Q�/�Yz�ס������0�A/�Og�Y�pC���ƛ��I��J�w	�MA�	M.��8>0�+l!u1[P�y~5�@���#�Ro=|���7c��v��uS�*U��5���b
 S#o�����r^�Ӧe���<]�}�e��$\90��+��`���#��v#Z/�|ݢ? ���:.&�I�,�'������@�yP���-X3U=/��z9����$f:��IC��)(�X)� ������`�f�e�����P�;��Qro�# ���P�	m�C�k��Y,�$��Ծ�3���؍g�Q���^�� ��暷�~2�n��ш��D�s�]�s����i������gj-N�G���	hy8=�m�������r[�U3��R���\$cRS��ޠ՜ٌ��_Fh�1���D�7��2@a��c�xtDqAE#�r�N8���oH��k�/#�K�o�r:�%G���oZ��.b�4�L�9߹2�t���I!`W��&c�s�;�RqҖ@�xS��^�{�ԬpZ����,	
	�g�p���e܍}�YW&�'&D]oȝ�H܈��Ged��$�V.�
�P�ķh�nM�?ѓT޵*����R�Vh�Ƚ�k�l!���_�`$jM�
M�O�r��x��<%��1�li���zR٬~͚j�姀D�FS��+TI�V�
0����\Q�����Y�]e�����Њ²y�zW9Z���_�rʛK}�M�e��`��A��D	7��Ep�j"�ے�����q��E�4�����'o�lLX�3"���\H~�ID��_���'Ry'��.
Ir��.ih3�`]0�r��<�%sn���9"�"�0eQ��k�8�o>�%{�.XoQi����W�d��rt��<\�@*��ش��)�+�A��
��0�?�uș���5��B�K�i���C�Z,��Ȕ=A���1�D�dzMz|Hy�@�?��0N���zǹ�+w6-�>Cᇗ���V%rQ�Φ�����bl�P.��������������N�d`�1���x�ee�o[H�h�������{bk+�	����E��:�}��֔򑛛����ꇁ���:M1���p��iM[����)ngu�n�r~��0�d���h����Kt��(�N�WZ��6-���w�D��ډV+�����|��L����^��� �t���j�����c�b������Ug�ŭ0����A�u��������D��x7,�dgZ����g>����␫r��;�����rL���9��e�z��YY��1%�~�V;���o�`S�����v�-&��,˱ᨬQ,h��R|�Э
�����y��y`J�Y��Lͬ�,�m���	DI�'��~�|�#w����H^јo��CzzAZi�>Ç6	����r��[F�x�!A��uJ����)K~�ԹM$'ۓ-�o�ln�̌3Z��I�2�F��3̵mb��5�'����{�(�
1�Ws"ǹ'�����U+5-o!��3e����t�B���~���2�e��|&���QK�'�z���V/�ea�������K���'���t�)�ft�«�DYz�v���������kF땐�?��=(�6�E؅Dv#�>�xE���#s��(�	3� �ڱ�4r'z��n� �A&�3����H=�A���?�����W��3����!���W��3+ZR C�j��X7n��n���`�"���^��z`�+�,��#�B�ô���N1���V�v�ӯ�7�h�:t�Z�����_J�}<�����D�:�Ç��N!����5���~a��s�+zЊC���R LS�c��5>-9q}��(�8�O쇷_=��<�1r2�Z��A �?4�X�4Ԅc�LQ0L�b?�R5�9:^8I�.��/�Z~���F)���h�G���4�)��B
�SD���믤"-���n�y�0c�܌�W�%��*,~фx����7���o"5mHh�����O�C��b�zg|��@�+gJ�]�l(2��sp�W��i�q��],�g��o��^(�KY�`�����������b-K�`i�-Je>%�M&l��4�Ƭ�d��a�«F����1��)�Y/~�`(w'25OԈ�Q��e�!ڛG�u�5_�4iO�sR�u�4��L�"�y�����Xf��@�DF*�2�l㢝@m'Ι �h�P���!^q���)�̪<|z)��Q+����q�r=s�ڲ�o�c��'7�p�	y����P#���	\��ώ����>�T��-$��gfú5������z����-��A�7h$������ڣ�˜�r��=���s��X�H,0e�����y�A�@ĒN��D��^��E����	�DYdw�rT7e[�F$|��!ɌA£���J{i?����2���w|����tp�W��66ҵ\z���ö����7g��������A���wT%,�º���v�`�����Bܽ�i��$���	����� 삠ݯ����IO�	��� nEk�d�r?�l�:��m��ƽ���K��u}�25�F�~.�}Z	���)"}]<����ܦv���zw	bJ82r�����4���G�?��טMB��j�0|�C!���Lm�o��UMY[,���"cY*���֊�'�
@�
�J����z��_��PK�j�~8jy�X
�G�udH�����{�R
c=��kXr4zJ�8\"ޔc}K�&EΏ�/d;�.F��b$	b*��z���ģ�rT6�S���y��&��!�ˤ+�=��ɂ+���{���S���i�q�)S&k���������������q�0���.k:\�����`�EX?z?3�m�����^�Q�+��7�����Nx���N�Pӆ�h*��4��l[1w"����-����W�9��+��z�&!�}���4�XV$���׿�Ŵ�69_�.�ɳN	��X
�F�]�jgj�P<l���(����`��mo��-T��Q�U���l��	^��_:�KJ��h}Epc4�aҝ�l��o��JKjH�1�0C�:�@wR`A�lV৏�O|wn�7������]0$o͎m&�t)��@E����9�>�f�Ԓ}�	h//���NC��v\	���;EOw��,��~"
��r%2�d5i�"cE��8/�&��8A����ּB���u�}�x�<ŋg�PI��I��]�z<��R��!�M��,�y���&|^I������1�5���Z��y�q�)�$�zY\/h� ���^>��C�(ײ%V���<.E��W����n3C���B�b���j��l-E�0j����,u�RZS�	P��־݈�2�I�%AB�Y�a{`赊vm�dyk��z<��Q� X�3C��Nk8��2�7�]�_�o�~��S۝���'I����I:�h&<2��4�	D�a�ځ��fΤ.��x��
�Ŗ<�r�����F���	��"p����>#b\�����RUċ/���A�X���}Z����r�\��U��S���T���W ��+�:VJ)5 ~c�N�O��&���1:��L�^r)[_Bl.n�ͫY&�3>���yq[yQr�.�4��w��g����B��XRo\��ݺ0�)D�R�Z0�Y�BD���)2�{���ԩ?���F���>I�솾��~y��=� U�����Ȱ���$g�s���o�jקD#yg��z�.C�s���BS����n&W��Xy7vA����A�j.�7�]�\t�{_����7xK������"A ���ï�s�J��g��yxqɹ�v�3|�Y�(y2����ːCN��p����i�3���`T�2(kk�t�'h��,$����H��sȠ8i���_�0)	�eG�=&�Z�K2��Z:�(�"�%��� �^F�'��d\����ڄ���t[?w����)�ZC��r:n�����0-�Ż6����LX�vtX|\��>ڬ+y$����K���ퟒ)����ϊ=Z�9��[9|�sv�ד��Ss" 'רϐ�݈AN����n�����0��߄߉L���.��ؔ�V�*�r�$RJ�Ɗ���9i�2|����Ļ.��n �!%�f��0�3�rq�%[B��X	���A/@��ǩ��.��G^2�؅v[�O���6�?�� ��Z��Y.�0��Wok��Z!��B�a�����e>��4�?�"�<��%����~O{j�C�h��:0g�a�Dx�C�y͡�]�Y70��U7�k������A��^By���@�`j\��4Q�ͬ��a������?p��o�2d�� 
�
��i��SQHoKz�kj�{���q��4n4f2�y�AI&W>�[��Zr	�5^Ē������\����o�����*ڑܿBb1���x���6ģ
�B����������	Zs�� �
�$��4I}U��{Y��rq-�Bw*[*`Šh��!s �M*�`n� ��ز&l��"2~�;=�\�����.�6�ΰ�W��+^�m��?����t6�ScP5]�H�����F�:�l&�ʫزf
�1�q�MWݤ�N�6���\�oq�T���㼈��Ϫ��#F�r������L� q�tP{2�2G�*ƾ�.a����/i`����;V��|��11�M(S<����2��Q�'i���S}��-'Ńo�g8��b�0q���b�.?�Nx[UE>g�BtdyY%�L`Y�l�Zf�	�����e�*�v� 0l��� ��8y��st�z.D��@����T��uh��6�s+�5�&2�J�����b���YV�v�(��4��K���yT�?��pV�)�B�B�Fr�k:���.A�K^�o5�
ɍ�@�l2����>V�Q��e�����P���T'X���L���5�w�0��
�������L��C'DW�4�fX��)�01��Bm@���-��ݗ�:l��F�����p��������)��Е��#0��걚��U�Eǥ�a}�P���Z��H�E�B|��b^�Ar-�b�sW��[��H_8-��D��!�'Ͳ��9���V��iG����f�щ{j$��n�$�t�QQɿᙜH�{�Kű_,�`����o�����lP[vO�m`��;hPY��?���O��;�����£���gPOw��P�aqK����hWQz�k�#ۯٔxok�;�N�ڋ l���J�����e�+�[#��}��p*�*�wb�߅LuTOۚ�VWbHΆ�Vm^�&���Z.��ns^�W���h��9��z={��ά��8�8��< ���j[\Ǜ��i5��Y�� ��{X��e'퀘k@��;["%VHYA��=��{k�<+&C7+�i���>ˑ�DU�;$qF�⌷�W�g�����L��	D	P�o�)AF��k50��� 8����#�<@k]Fl�� �	�4|	�m��I����@Y��S��o�@Y!^�ie�/�YY�PN��ԕ�2�Y�3�'�~v����n�Շ��k�V�,$�?5��!���ZۑOgg�`��U��$���6�F�x|�~t�u�v�-�|A�*�Y��f����������gW����D<>X���Hc��ƪ�tz�F>
ŏ�������A�YP��."��#`jPu�S軳���duX�į�7�)�n� mXi,9'��:�6%e�M�"+�Q�$�/t�g�Vj}�&硭ВR&�-vCko+�4b�l���}��Rfr�9�a��X�
0H��A�V-�2�d� a*�i���y>�r��h�0Q�XB%�6���5*w��@kS xV!�� k5!�P�:���<��f{�~=�8���K_T��n��vQ9
`��N~5*�Lr�1���ۻ(��%)��:&p
)�x�/�FC����!��f��ZBu���
��>3��+�vV���+X=.�n2�cq����|�ʧ}@��(� x�����׶"c.�6����8AN�5�Y�"Z��'�Ǡmm"%���*#~��7�,���ɲM�T;*J�&��nIcZ�^=m��,��N������jU��!��$'S�c�i�,e���푧K�ƺ����Ѕ/؞/��T�[+k�/�5�x�7���;ԫ	R�8i\0]�����D�^똴.���Q2�J��T��Ø��ܜ����r��8 ���U���N��2�1𾹷��ENv��--c��U�c���� K���,)���)I�����J{�<��	O�b7�6�B�	�KH��'lcg�����
2O����Я��*��g5�5z�[9I$3�����Dt��I����LH�3�E�\Ws+��9���+M��<L��#��-�آ�5� ��F��:���\q��7>k�l���C��FJw.��T��̫p��;��5n�ħ	A��y��ҁ�_��3..ۥw��L&�?;�w�T(.^"sG��#��{�D�o�U�s֚
,8�������3�(F-ȭ��	��`\P
U\m|�a7���`�Xths�� �'�5�2�@t�Lq�|~��2+�~ٰ��'��7X#��<soW7/���?!S���Z�/BD[e�Cb7��{GmNQ;-��;����#97v|��Ku�]e��dEӰ=!JGzc��]&��mשq&G&�lW@��h(���U�����Ù~����J�1�PM�*X�Io��Ґ>7���(�6$뭂��`Z�)�4$M���/��Od��C��G:}|T�4Zg��P�4���I,��;+��퀰2�v�V۠�\�u�J&�3�i٣�s�>�\�`�g~я�[�iͱ��]��Ҥ�X����dIhHp��z$����}����?2�D�󀠊:��E��I��l9=3�w�Z���y�f�-a�p�B|m��U>����z��K�Fs����8��W�{��KdB�ӯ��aKF����k���Ԍ+ٙq�������,|�'���錁�;���V���wɑ@-�j��Y�c=��"�I2z��3!��@��fME;�c�}U̕dt����Lm�t�D��\��rdJ�>��q��&���?��3zD�<���d�
���z���T��j�Q��Iz�CV�*7N�_�Z���d�	ׂ���A�w<����"V�+X龎I,��L,JaC)���[��e�Ǳ�R]����X�ɔ&�*����Cpw2��C4�<*Q�N^�c0�� �U�;����9��cة����XZ��=�"`L�)�In�_��<*2)�f�L
�S�P�Wm%��k�Xü��\�":��SU��6��p�H�?���(�W0���K_|�ڬte�8������fx����Aq{���sgu	4�ۼ*�')-0��#�P~]��S}���>b�͂�Q'�e����(#�O4�ɪb�hU��ڳ;�Ʃ��Q�w�C�f���T`�e*�ǭ#s1{3�=Ěk��0�_$>�J�U��[�ezA�T�h�����:�䑿�x.��8��,�:�I�\��Wh8�Gm�z�r�:n;��14�X��n�*!�;��"p���g�D�rΟ}:��/�@ti���Z��#h*��[�C��Wmq�`������kWѲd�W^�W!s>	��}�oz�}��`��]�Y�P�2�HtHm��1�c[�ï�>���<P�C�O&�0˙�U'ca�3���h���j~^]�j��)�g@�d�"�ǚ@M���.�T�k��l�͜ $���Nr��%#�a���G4���X�֠��;���E�2���;�,x)u6A�-|]����X�L�]��}I�Q��q��}xH>y�o��[�b�+ê�����i�5p�o�%������#����Y��������+=	���'>M��Ҷ04(�k3^[��>�鴰f�I�	&0����f�鹼����e�/�4��N���Ɨ���7&H}<ҽp[fr���-����YޒN	�p���?ɕ+�`��JMՠ����n��3�q��Cד��@���n2�=�����հ�m���WK�2x�"y+���j)��0vGN'
À�h�3x=�y�M�W`k^G��ԋ��nS�AI`ShT2V�i~kA��%����T`M�t,�V+��4�4�>�}���WJ^jxu-�ms"��J)jA�4E8��`.�����2!�hw����X�÷�T�B3�T4��xʎv�����V�9�!:wITm�!�wD��6+��dN�W_��H���o�11-�.���-��9��|]̵�6 Uk2�g��0�`�^K�hI�l��3���1���T+-����N���H%��U����UM�E}�i'�}"�ֻ����������|��3�P��"�G�	��9Ep��I������_+�r�~��}��h\>�s uS������l��c.�3���mu,��X1�T9���+�Q��Ճ��R�&��+(�T���M\�E���_�4�4�����Q�	�,�y�;�[��ڒC>`����!�Q-�#����w�|�
����T>S�S� (�c.D_�Ƥ���+�MG��i��Ɉ������B�j�W��%���VJ�aJ,;�e bѴ�f����f�&BC����ۿ��R��X��r���{�?���=�`��9�2_�T�"d�m���8dY n8j�B�py�橅�/ ��<~k�p,��<�� ?�rY;�[�����|�����5�Q�][qdv�P�=����k�+F �KhS�Qڒ%����lɁ�h��wɃpl��5*��Тq�2I�q���R'��g�Ҥv�nSP���8|\�O���J�bй���ר��Zp�,�R���Ut	���i{d�Z_TW���MW�r���N���\Z����_��h)h����j���}� "{*G����:<5�f�=w��M�h)E_�W�̷淑��6��!]#<ZOj�؂.�p�gO��9�>��EW�0qd��]vSA��� r��0�w�\᮴���V���;��!�]��
����ng�)�RAI٬�i�o4�P���ٷ��7�?��� 
)����F8���i�I���!�:�P�2�ui��6���B��i�[�y&ܢ�n믇�,_�~?AbC�ghDu�'Gy�/���A���q>-�;Þ�]k�����d�t:��'�&�y)+�j����:��w������<i}�����qږ��ҳ�$���<w�\��<��?�`���I�u>�l	�5{f����N�iӰi��|�����Ȯ<�N�b�0��v�ZN1,Zv'��|�J-ܯ������5��B�����MC�)���S{�2����!�u�DY��$'���L�#�����CaN�	�7 Geboj�uƽ�+��·�*��m8�{���ų0��4�빹e��K$���iꚿ.��7{�f=�����z�q ;+ʟ�O~�t�[�"xJ@�bR���x�L�;3����6U�>�t�5�U����A�2�o� ��3+󺒵Y;̉u��^���S
�f�?)\ش���|1�l�ibXqj���G�*�~�����U����_�q9@�{�M��������#oc�8&�0��W���fg+K(�YYCV!��\ *(	K�~`���η;�ϱy\����,�gv��c�a�(�P�j=�M�L�D��5��i��ݷG�J"�藌#��V�+ �u��t��I���"��^�]�9��t�>j�M6��|�.+G�M�IS�FZ����BӚP�J�f4����"^�{�]�� ���X����4#8w�A����Vr���a��Y���\��(힇	�y!��纡$Nɭ���i�y���#�%�*����qEo��
�$��Gµ?G$F��魬,�i��K!B�����	H����׶�����p����U�S��,�����Tz��[&P�sm��Q�����I��̓�~ �)=~���L\�E\�Q ��_�B����dq�Ei4�N�x�[�&ٙ�+�H3�^Qu�#d5�#����+��EƲ&��p�>K$75����K��$�05r=�d��b���U�v��'R���k�g������r��N�������a����(�����
lask6�Q�u����%��N��{�}b�*�Q���`k6��<>�7�abG���%�wl	y��yLlK2pn6Y�i�[3*�S�����#� �W[��I(�ɵ4�����c�Cn��5M�3�<�s�� �� \��������v2�6+P/q�WaK���	 ����
f~X��FS��>�ܐ�_=�F�`�������--�=�c�A�kK[m��ߖz`��_�G����������ӈI)���x� ^3�`W��Y��Z{��6��z��1�t[f���S	=7R[j���5�)"�_���-}Ø4�k�'���p�a{�zSo_s@��'@��p�hQ7꘶�`ܟ��>�b'M�@�x������A���9�בg��轱k�]�&,T��&Բ����+�#W�T�\��k���9��T3��i�O&8�D��J�{'M���@�y� �|R�a|X���cnZ���<��f�� ��,�_l!�����Q�������Lm"����:��6� ��#�-��C��*� ��仛�,��͎OZ��0�9�,��L2�Wξ���6��ȥ5�9!����W��$#����mB����u�Y�0����(۟�v��︘G����1m~f���!(`�4��)D��&"E�D~����6F �	YE)A^	��`5�J_kC5��t��V���q�y~���e�e�Hr��f�vG-/���}�5L�H���⻞�� P �1O\��d^ �Yk�j<3<F�q��]gG�7m��W�m� ��R���G�{洞����¹��L��Ҏ�8��҆�?�Ms� ���p:��u��6���0�{��U�[R:���j���(���pѠxfs(��}O���	���T�J�����a�/�10�rf��0,A��6���\ڂ�iǛ����L/>b����"��^{�`��A��a�������)��+/|1p�󝶩	��2YX�^2�j�(ѣA�X��ۤ<�&��r#~DW�{�-Jğ�h�OcIl����ҩ�NgK�[M�#Z���a*����FbpY��W�Jؽ�ɍF҆����l-�A��u�:;���P�8�D��^�4�p@�Ҁ�dz7��:�����58!����P`>���C)�u\w�5Z�
�*�S�R��?��W>-�,΁���s�L|���|d�J��P���""u�
/��48з�U4J�5R�נ��ɧ���W%���ґ�ǹ����b8�C;���� ��3�Ұ�w��FH0���]J�VϺ��8"����e,Q� ��	�]����'�i��4���e��;}��GL�w�6�	�N�����1X�:;=E�@�g�	�F���VLӐΒ��F;V8T9{��n���e�͸�̷Yƺd��84�P=L�מ挹 ��\��CI�_�]j:�[;��v=⮉� Cic�D��>jh%jR���8��0�0��|�&.�G�q�nq��ev��1� �ȁk' ]��|�c(n
��W�������{�,�'���*^Z�������}�=����_1>�Z�t�C�U@R�c5_v���C�,5��|�^����Mpz�����m����I!t��U�i��=e�1#^f��Hڴ-p��z�ؾ�:X�8��^ut�=��N���I�+�eBz%$��G��ӛ���[m�lqN��,�`鉋N�[���'���۟���k]��ʹ��q�ՙ�c/n��^l�'����E����ixQk s�%:Ms�Ӡ#�,�bN�4T�p[Jkv&���� x����'s�.���{l
��L��
�C$��{X�a���'��- h�ׇmN�-�;B\��Ω0h�H�g�y��0^\�.ݿ���}a�����)��
Ѵ �dI�4 fL���h�W�+���>O��Wr�Rx�W�a�5t��n�MM�����X�<%���2~:;;�����;ߢ,��+�O5�9�i���9 �V�KT��{8@zx��sW���l��җ��������C�v#2�q7T������,[`����WM�Y8�I����XQop��\�1|��17"��DNasr��J� &��oؕy��ț���4�m�@�:���@ڦ���%l<�n��D�p*:(3���Z�iTE|�B)R�[�P���:@�jm�ۑ���ߍDw,�)�j��7R������i�BvU+�'���~���X�4�2�8�)�Q7`3����
�>nU���%1o�l��������d�zk����Q��'�Z��CPY�2&i�,�-���挖ԟz�����]X^��MQ;k?����2;Y߂YLP��ъ/�`�q�2���hqi�
�|g1�{F�ǖTy}X��J�Oh`��y=�e�T�>ryJ�������ӵ�q@��hB�k�w��>��5TS�����jQu:��V>�����b�w���:�5"�j ��K����}*KM8 t���d��IwU��#�#s�;�u¤�E�X�㬒鞿�� 3�(!����r�5������J�˪���p���J�qzۨۄsxɶL����Y�p�p���+,�d]& qn�)�N�'Q��1SIV��5�� B��fD���#���w?>+��	_���ͳu�m�?
>��3>��߉Tڤ��r�1��G�kh�Iv�G_/�����}����L�g��G놇D+^�!��*(�"1G
��������Aͯu'�p��-F��o�76ZbC�:�l&����Y@x�L��i6-��Idf�Q'�����F���$:N��m��9)e��#fb��+�<rۭO�	"�;��ḏ�� ��?G��BR��/�PЏPYL�^	&�0P�#�0�ތ��b�Φ:#ơ����@GA��?=���v���856�=�@���)˸��&��P��`k\����;R���T���}���'�
֥�w�$x����$�&�>l^h�Y�=4�}?��OE���d�j����^�v �?��s�զ�T>�+<��B�Y��l��]�lU�gk�머�t^���/<�y'�"3�*���D~��[������V����@�`ek���R[��ْ�5D��62�����?R�,�_(�c���ֽ|K{���	/�ỉ	��"AL���
v�a$�cGf��b5����G�(�Q���x�wQ�m�?��9|ZH��\�o�!�W[���nV��� ̈4�(O�P�j��r����۩�vw��LD㠌��?��.*�PP%%��x@���h*�oUZ`|�!�mح��,$^.=���m�b�/�2b����h�^)������w��G�X�\= 0����(�>���������X�R���f�k8�6!T�LE�f�/��#��1���%�HE�{X��0�ɅZPW=�&���z�@����9��`�HFF�����7��'-_>�V��;���S���e�W����󯊄e=a�/���&U�,̂Ͷ�)rr��p�5��`� \����g7d��,�5�~�7�td���ي� f�~lz��"�K�j=u�v�nZ%�Γq�8���+�	Y���kŪ�	Z���w|���q=��}K�\�� [�;�(�'F�"x����J��H�r��fZÿ3��� Y�NV���k��0����E�	�ߘ��4��}-ӧ����s�e���+�C��{a�|�($_�͖G�5yk�>���bZ�����?Շw[�=�nP�z��p@�c:WK<8THbp��y�;�Z��|�sȋ��ָ���V�R�	��eG䁧��Lx��}�A/iWf�F|����N�p	���u�C�F�Wõ�j����A���Z�Bq�`�i��⧚�hM�)d��&v����a�5���x���Tk�d��yE刷XT�[r��_��y@�cx`�CB�i�)��XDi̞�����4s��-���\(�����-B)��'����gDo�싥1B��@uk�J��Ļܮw$y�;�>�0{���0zD�q���??��:K��h���"S�� ���+N6L��g k4'0�=�;C���(��)m�r�y�d�J��>lZ?�z�V0���TIU�1��Z�����F�ޛE���f8=ˉX=(�lnlĆ�=����hv�����<��m3XԽ:���΃>�K�!��Y.:*����\�r�%3lA?p����sj�.ٿ���U����7��v�ٴYGZ�=l�>V�
�8U�ʹܟ�ar�$�BG�ޔ�6�Ǧ�Ood�g0|���� N�Nzm��9��9�-2�Q$�_���f���e=쵚�����A�����c���� x_�  ��Oxa����,��	���%�����k�l�{.����g��\�Yb5J��ȑ���n����}��߽�ɑbV\�P�uP�=���!c+95���F�&.tD+�F\�x-?@�j�H:ӧ����dU3�5�Ή�ؔ�uw���&�C2�~��w��_O�=Ճ�HHX�ܒk����at���nc9�GM���W�X���W���~+=>��4���=�uE�l|/9��*Z��E>i����wPg�>���K~TR���B�2���<-�ȭ��p{�^f��Mfa��P�A�������~M>3I?�R)�s��6%��XطХ]�N[�Ы��@��S۠;��3��9��t&��`����*�ؐ�us�檀qwvP�,@�ފk!ً���������+0>�H��	���=��m�+�<ũ�:�є�|`#�� 5�(j@��|B�D|�NǶog�6mº_�6ja,�P�r`vU�c�`���Qv�<5|��@�*8U�Z#Ű��|��?�2*��o�q$b���.��x�ݶ�dIY�J�K��qc�?]�͕-3D2b�83m�%ض�-�hO�(w��@2�*0���/�N
�QGcf���3���3��R����y>�ډm����'w���_@��b
(�������F%$WV9�
 �����髗��_�ǟ�Ԗ�ތ��*?R�zrV��z9������]�h4(��� J�<r��w�J	�}Hk�F2�M
��V��\��0����=߷Kw�$�q~�"}@g7G[ٶ}8}Y��mi��l��M�����>V��}w'8
$��Ǒ�> tpٗ���QDmP�&w�1>p	�o��-,�ܘ�o��M�W��5iK�B9�L��v�r��A�ԧ�>9X��^\�5��q�@ʾ3��h&o�,I��(X���X0�^N8���W��-rW�7�}��I;������#�B�D^����'@W�U#�`B�+x�ZG�r�}�,r��������5fgD���)�Qq��$D��w$ng�p�[D��$$��8�ZB�L��пb��zφ+�˹cz��rw23��Q�#��~9���[��~0iS�ח�gG�Y�)נǌ� +�o��)�EC���2�*#�n�@�4��6��EM�v�x�����#X�����M0v�T�zԹBL�����u�����k?�����E�i~f�VD�f����^�Li��W)����) �w�����ߺ�c���yU>�lm�{v(�}���,WNO����\�����p���1��nxż���Ǐ5�Ii��A�I��2^ �vo�e��op%��QtH��q'pC��<"'{�0A�=4W�:�-�bS&�j}:��T�e�/�)叆O8�t"�8�
�$�ђ��ꢽ!9ȃ��vg���Ut8=�	.��0��0�8�I�
�7��Z�Zq\�����B6$߫m�X�Yɦc�J1�����X�=��
F�8�}nBq�~wQk��b ���?�i1VA�RГ���٠7�"/��T����o
Ӻ��r�����q��f"g[��ʻ.����^�X�TfQ�jֻ�&{�[R�&#Uz��i!�x��T��{x)0Ӭ�Fx�n��"Ħ�� ?2O�6�f�
����Zs��EF	b^	7���C���ts�¤�:��w������;�$����Nc�9�0765Okv�Ga�r
�?½u�(�zuϰ.B�iV2�돯߮b����3�r��p�P�i��uB���K\"�	��K:1�}����&,gB�a��p����
���F|[T9����l3�}K�}֪���s��~* �1��>z��֗U���g� TX9+���`DM�xW��KP]_;�'�t��
���L19��_�Y���� h�4GxceQ���9ӾW�bJ3����i^X�K"���?|�����R0�h���j����t�:���NfZ�ˀ��o�2�݂=��L-;�f������cR2U�e�Č�*W<��2cV9�E�8�A ��(�b�JU��"�T~�3]�`��-U<B�i��'b�cx#��-֐�l�����B̬��o�X�WXPr{�}�0^�C�L����z��O&���%�q<���,|�vR��[�~��1^��c����h�t#H�Ʉy�v��[��kAjF��q�p=�nuf&[�,!/g�*X�/�h�u<�>��%���UyM�3���n_�8�C���څ<;2z�	��o?�`f͓|bt>�1w�'�(��eA>�S�����j)r��g�����V]T[�(EW`?�()� l�r���-��)ZL�&��u�!�
���BL�N��88�w����ѧG%��I��銩 ���0ky������6�B�l�s44��7�Ya�gh�2�\���PD5Ʃ�>���.�Ｖx�h����z���5�Nr"�[R����bsf!�~������UZQ|�B�s3�1��F�A��c%��5��㜅���G�Ih��xT��n�+^�?�O'���̉��xҠ]�����!� �j*/�Z��UHǧ&���"3L��T{��ȭV�
W�v�V;/1����TLZj��Q�'5�_j<�ܜa%$�h�3G:]���r����1{�f��aLc$Ѣ�����C�d��8Y LF`m���[5s���QAmF��f���zMa~@��n�v�{X���(���Rދ�y4���N�8�a:V�m�۱ZM��k�2�����}
�ǠСW�a�2���}�X�9���2���l��. ���4�k��v�<��L:�+���b�� ��f_"�Pr 
n$z02�:c�_�]���x:E��+_n��7|�D&�5�����!�"���]{����)���r6^�V"8�0@��FhЊ6���r!_M$"����v��\���J!�K��:|B�D��N�g���جa�t\FB��[|����-D!%c��nP-k4c!H�ͿƦe��'���a��q�F�3p�$�0�H���FL�+}L������_�l#B���3���*�U�����`l?�Wڋ�N�e�b~���Ñ��P l#�q׾����:g&�	ě����F�Ң=D�'�a��~��v�$U�2��m�oɗB{ŃwB��daS}��W�H���T�h#�Ǫ��9Z
JO�9&�Q������HK����t9�����|�Pa�鰠A̼�e�"�W���H��̀��Mw6Ş��g~��`�G7�`K�	#:�X����� *�.e��Q$┺��g��1�?Sb�Q{�uXx��ǿ��{)�ߌ>�x9�q�mߖX[��N]��R!P�b�(���f��������n�DR��tE.xľOy���c�zsC�ɧ,��}�o��Pk=�0FIή�(��}u/*���U�_��ՁhehI[!��(u�*��מ�sb�=ܞ��Q��˧���Y�q��������m���?�=ZSF&A�c�I�7�+%PR�u,Y_�
q�i ��V�̆s��/�br���Wb-`��Z���77��i�S��Z���5�+@ݭ�'Ʈ���h-y����R[����{c��v����{=���# �8
���i�����(�jOZ2�M�"��-&a��E��˅�g.���m��H�����B���B��2��G>/���t���g>�Mx]�aÒh���+š�(�v0�\�`�d�j*4�8N��� 5"	wD���#&Ow�-t�cET��6ɥCRV)�Y����ù�$��W���ق���ҩ=7�=��gEri�+Ai�g�[��U��!Df�xZ1j��\�wW�'�QJ#M_-��7
9S�����7�"��c0%�x���ן ��0���Ȃ����ݤq�9��`�J��`������O��Sa	Sn@NK�~��w!��2jf'R�c3b�����5�v!�]���}��s��ŦwQق!�f�*���g4/�*���s:�7�+�L�ǯLU�K2�5� �3
��!#��_o'�b�8)t���i���P��_laFT�Tځ5����r=FfCw��˥��@�V����@W�Ό8p��T��>$۝q��b�(�r��'x��xT�Iy2����#�d��}cj!�a����a�A�}�7��7܂?�3��Wήϣh�l�i�٩�$�XP��;S�9C:�X6��i��Lt���
�)=��9�9\��%W��2����W�>{�c_ԙ���S��_l �Rw���"I�Ч^����
?e�X��U|\��:q�T�P�9�}�j�i�x���ף�B�N���f̘,nd�ǚ��p��KG����>I39? ���̡��|Z�Y���֟-�FG$��(wƟq��-�^'��X����> �S���^r\Y��yX�i<iȤ:{x0����j"��Q�p#������>�_Ν�m� n��$'�s�(�N�]��Pۏ� ji�lI)��6��VN[�y��k�in��aH8)�eO���ON��xԓ�Jnĕ�.�+��B� QzZ�T��$<��Zd�q�+����4�/n+b�/��L[�B�T����p^[�Iᢚ��H��:�bn<@?a���^���%�^��QjM�f��]k"��J���m�{(":��,y�:��Zz
���O9@ RjE];��J=����J�r��эʁΦ����=�y�!{�^\�vr�Se]t���9��ͭ�L��\�Hb����[�����yf"��u�j�x�����z��2�Q����B�/�sB
�b�G�o>E��J�	u^��"zG����rG)�ƚ�y�g�Yi�_���+'_]W
u�����t�*`��/����"��e��0X۵0c�M�?�h�T�c&4`��G�` @�\���6�f��9�׎ �d�}�L��|±Y��5O��ayM+�v�~���J~(�i�2��̃�4(zv�Ն���a�R�
M��_���=[�����>�K���{\I 't ��5l� ���D_�p�K//e��X>�lyk��YV�E�ޞ�̙-�F���d�Y�& =󹿃�������ºN�󤮕| ���Nđ ��W�zZ�w�^�a+8����H���jD���� ��}Ԯ��VC�c$����<�U�Z,S����<��_�h��鹳��.`Q�Z�8P�/�R�l�����G ׬ 
�[�c{���_��ADh���I|�at`���:�o����7T�e���\����1�l�u����f�_5LMtt�����js��>Y �{(�7�[ܑ�,��"���M_��}�UnK���A�%U�j<��Y\�
����j����fR�"~:KfE'
�/�������=��C{3y�! ������>���Q�
������@|&�E��1�J�$fñj#aǬ�����[�b�o�B�2�J��3�<�����0�XFa��o@���O�u
�	��L�M�m�����`E��+P�Mė�?��:xRA�:n���
ˢ��o9ޖ5;*	�r��A�(���aFզ����Bn�P� J@�<��A�B0
_����k\�F�/%���\ӆc����S��?I�>ה]��l\8���"�)�V�@M�p�r�M{fg\�I�r<�o�+�1���������}'�kϴ��,�]�B�Ё��uW�ËH�>'���vD�^o�%�̡��C5��v2"n�P9�릧��Pw��R�����#i(�����Y��׆X�b����Ich�Y����p��o��O�&q��Ӈ����.kM�`�3�Іn����T6�E��P5w?u�y7Bj>'.�Nc���wΦ_���	��5HDO��wE���C�U,�T�䩟t((;d�>@ ����Y�8�&{�G:Z��w�Z���=����it�:�'92ח�	UK�������n�fwb�1�P��X2�V�%�=+���h����M�����x��V�SW�VsA\`�o��І^����-&.ܰܔ>%��?GW�;�7Lt�ުS��gl�sU����`��Nu�F�̧��E��#e舲:��ѾD�#��c\�<&�o]D�c�j^/�x�	O��u��(�E �]Ay���Q|�kpc�?���OL����C�A��׮^	���؋��鲨Zɫ2��h:��׭!�mv���d�HE��j�N�Hb��#�Ʌ�\D�n�P��g�l½�Cg1�wz�}�Nہ"_^9ғҗ�m�ލ�5��݃�"n���$b55��=�O
ʦ��
ޓ��5�M�h��Cq�g0�n�
���aP�j�q�
�,M���X�Ñ�g�u��t�Ɋ�#&ǑS���=��`,�w2R�РE�aJ\�Az1M9��+mU��cmO�%�g8�ݛ"D��y�\���/�������:�j�|�Jޖ��ȕ�I�K7*�v7U&+�v��_iZ�/վ��.Xg9R�C*��_�tп�4]��`�nC@����f�H�}.��p)�������t���5DZ)��y��<�eG�|�A�W��"��*Dg&�h+�RR�W�0�Ѓ����R�W��)��`u�n�zmn���F�5ElG��9���A%	E�	f+�Nh��<e���
d�M�G=&ܺ�F$u��4]�t��XG1�������̀`w�'�DjEA�u����k9� ��f���v[+%�>⪶
��t-1i|
m�2������s+����k*��������]��@>���k v��Tǃ�n?�I�a���X�V�B���ߊ�a|s^����&��5ܶ�����[|� Ĥ7�?x���~nW��@78�����ƍ��j��w�Y��cg��b,�R���x����$ò���m��Au��̔sxB�ۅ����� ��p����xqu���Ŏ�Cv���I�����<m�??��6`5���iS�V�t�a�w�`�ɝ #-ЪMv]x���ӿˍ�6n�(J/y�e�!�ȼ3��ǵH��Z�Iᳪ������Q0��G��	[�#x�b�l�?U2�t."\�"�ZE����۰���BF�m�4qd���j� :�*m��@%�Q��&&�-��SZa��q]��q9lc<�ST���#�5D�e�1~x�7�X�p�e�34~lSu��*cU� �������5�a�c�Q�Th3�ʒ�k}�?q��i�Gs�b:�#�q�S�k3-
股^(3f�V����aK"��t�ܸ��b�#�5�G���Y���mx��g�<�ؼJ"C%��NG�A��_�\@N�a} ��M ��ʹy��%:�l���ve���3vr~�p[�\a��q���AJ8hm�E��M��p�e�|�Y��)�|Wؤ����:s�Z!թ�BQ����'���73̶�y�Yf��_�,��X���8�x�l�#3�rP�� 6��q���{�3<$:�m�4�����ZW��������
��ځ=.�R1�$��t�
��J<-f�BcfW�=/%�«���z�8�z}��%�d��6x�C��Mm�_a	��;:��}��QyMA�C��q�\�$9w�u��1�A�!��,����Ҁa��(wi����E����`W�!zn�Tȗ�qf(�x�%@8�0:�K� �C�9)��7����^xU[���o#o^E�4K0��Q�W|��W�L%�m��:��+lΜ���-���W�b@|�W�ﺄ;�����F?��[
��K��r�gg�_�\Z���o1%�� 0HYa\�,��4���Qd1��GA�!o�Xc�����ĶO��G��5s�U)�G�B�5��QA#T��SV�I�p׿�4&'���@�Q�],��(�
�{�2�5�&���̞���K��G�Q���~3KT?Ӵ&��S\���(��d��z
��ԝ�s
(S��س�]����lk��5~]}yٕ���j)'�舏����d�'7�k8���t��&L��Ѩ�	��T�o5��-܁�}���}
p:���v�a�=�8�'�]��er���;[/�ݪB��mƩ��d"<�|�U��bG�C��
����nϞ�K&I�\]����1�Y�- M���
C
��,ư���+�����K/�����*'-3��S�����N$�@��0J�t��?QQ �.dѵZɠ(���<�USp�Fjz��(���SZ{M��ڨ��g�lʱ�����;��s���46'�L���/\t q��L�}Fy�^O���K>UJ`C��Ezc(0T�14R�y=Z*}E#$�uM�h��)��(k��k�� tf�ڤ�r�6��f8��~-h������|�������/�P.�U~��|Y�5m� e:���9��i�ڟ���Q�	A�Hq/����u!©�YE�̗rި�(i^*6����5"��4V�𜷖�\NA�傌��
���E��N]t�g��MVio�m�ޙ���bE��v�MF���_�xユ�n;�W��`tƌ�캼m8uW��'���J��(C;��õK����i@�5Lv�j������A���NNF�䃏�r�v8��mp+l�Ԃ�b`%P��{�]M�ZV4�0�D��T�>�H������8�އH�6��P�y�S��C�N=�:j؍ȽW��������	 2եU��;�1�_������vN{ץ����YZZ�� ��F�j�2��-K�'t�h�>�v�lI񌛏���E3+ @�-RnN���ġC��{��O�>*M���OE�Ӑ�V��e�������z�@�O��ષӀp��#a|%>uET�z%kdͦ1�h)e}2�M4�M����A7u�����mY�YDN,��o��nrݷ�����=&&�H=�����3+6��Gĩ$��aZOe�}t4�}a�?&>��N�%@u�{ͲY�'�W
��'K��z���V���%^"�u�����Y*�rC�j����eJ�Gbɇ�5�P5�d@��"�;a�����J�:ϣ��`�6�Q�-����~jN�,�I9����xY��d���x>�b|�_�#��.����¢e�~�~!��d�ozj�(5Ϯ�0����fȊ��Å�׮f'��e��(SB~\�������h8ҳ{St ]��#�_�Uks�q�Ǝw��2�?ld ���2�|zP���-A.�N�j3�C���6��;��"7Z��xׅ69��ٳ�RE�od�[g��:!Z���v`i=�rRav;���O���Zq�@G2B}�G{�x�r�:�^{ƻ�"�9�j��<�C%��P|��L7T���.��
��_��ֻv	5h-����BD��bl	M�%i�l�Es8�=���X��2�ʡUbhx�A�­g��~��DBB��3DbiƐc����Y*��-�k7]F(�=�9���!k����k�q�{��Ɠ6ҳ���d��qA�D�q��1�:k�q�e~�/���%$��ą�&�1�w��R��$G����Z1j6g;_ǯ�}��L�E�V��}K�Qp����@�q=cm����Ʉd��T�Tz�7�)�d�>f��H���)����q�=��%Z�# �	qlk�J��v��.9k6�l�_x��Sp6����b^4�<=9�7�ׄ�� � x�O!��CH�0���r�?��L�ٸ浵�=2�>�3�� 1Y��K���>ϑ@�T�2���V���=��{'�n�u�E�,"�^�o��+�,���A��Ã���A�#���ĪЃ��� \��U�:��t�V��7u	��o��a��+F�Zl`�1���lR�Q~Jf��`�Y{�ge�����9-�n���g*�:1�BIs�2̲V혁+��͟��o�.�*�VC���f��[=Ϣ�� 8�L�A��^{��?�xE7���:^z�����)�o_�:��Io��h����dG;9��)#��c��a����W�IN�0y��V(?�
�;~n�C��7�����ڬ�&L�^��Os���	O�_�==U��ڷ���@*�WQ��8��vz��W�Β�/jm�6��ܺ�jeU�=dV@"�4iR�^sBQ�^y��I�*C!�Ή�(�E��ZW���v�OF�i�ΰ0��H�g��[�ֳ�T �',�ev��L���1���j�sV)����`{C���z�M��I��z+lM�\CzJ{�F����:q�B��Wv3פ�"����&���^�$39�zi�����Ћ��d�+K�z��a�B�@�ځc�O\Kw&}Z�����lc��j�)0��%���~����6�c����笶T�uB�e�����Ǉ�Q0�iz/,'�{�\�
5�z�_6F�����s?8�X1�zzs��ZD�8�3:���2U̣T.bC�򎨨��P�s"��Tݚˠ��
T���U8CU8Ƹ�i)8�V�f��%�sm�����=���W]4p�y�y5� \��A,�8��	p|���n^>�rb���z�L��m<��Rõ�ٶ�|j��W�Y�n�V���"&��.�r�G�ǎ���r�ދ��:1R�x8U���"����vr��>Ú��Rl�٦�1��-,�=k��� �&��ˀ�<��n�tP���<���LsɅb /��� .�/E��z���u5Sj��zO|�� r�PhG��+�0f����BP�$!a~�bU���|~��ALچY�c����4IR��oo��H�0��otQkK��f-�{�\c(�.L�Ͼ��4���5RN��;%�w��;����q�ײv��� ����R��u�5�30��|�.�1(�:�{�)�3��f�`��T�K�
��^�=R;Ĵ�����oS!��U�㈭E�6�%I��i�^������	vKVS���F7�BL$��t�W�%�4�	�d=UbJ�z�*��YT��]���Lj��i��b+��sꉿf�wH�O����*XXw8��C����gCք��T�_$��|��KߍS�=���3f��C�wV����H80H�QA?�8�/�;~����-P)�j^�����J|>T�g�)���0ⲇ�������~":�������n�1���,�[f�=�з�E���Ù�mvf�N�����A�~N(%E����x���S���+�c��x���d٢���ɭ�T�|&05LD|X�ڃ����y�[&eFyp���m���K�n�SJ��T29��=�@��5Q�x����AC:��~:8���p��S���WzmH�QW��.���`x+����V u)� T� 0��s�3��}¶␋C3�3e-Ӥd8��H���&�u�㞋�/��E1Y7�4[i�ZH��"@0"�.7��|�ҧ��>ª)�4R��H:_��D�8��8c���cf:"v뾽F����F�*A�z��(',�m'�u�o+/�O[c�gOH���4�HW8��m.��u��=���y�R w��+gmHO_:�&4ϝ�G���J2͖�J,��%����{�|�q�ٛ�0ֺ�8���><�pE�b��i�,�qP:�g�z1)�
�%4͒k�p�m.��x�P7�"���lz�\A��gOl�*빻��Dp�T+� [fp�ޤ$����P�M�(5Z��u͑:A_���Г� �Y�E���v���2N���;�,F����_�������g��; �$R)�+�Gј��>�)s�a:4�iй�U��C�d�r���w��o����J�|�G�}��0�CP��h���{�Z5��%5|;��O?vՖ���E��:�?�^a��� t��?�;���AU�%.$�&ڴ#h��"�p�Tn�e������D@�e�)Տ���R�3/�[��>� �?��ɓ������|�C�\bW���Q٨��[D0�f _��â��Jl��o�Hx\P��%��"�[�̕a봯���+6�"Ն+|q�7%J�(��K�����h}IG�&�ZM�4�J0Ԗ�v��X���k��g���7i����50��p5Ø�㼘�W�f�Y6�?��#�|I��
�"2$'d%��!
�m�6�2��* v�4E(��t$n"T��.����zTGW�[Yu���u�&��)v�#\4�?�����9ЈQ���[(�{L�8�$��J��겵˄c�b�����o�����C]�Ƨ��']�<N��~�X�����x�~L�H���E�0�
�n�]�N�>*rv��E��8��>4��Pg����AN��q'n?�u1�����#�6�~n�2>�CA۲O"~zfx�n���8��|}1[R�����@�A�jt��HE�)��L�!�{�4Y�o��`p�8��Z��_\ޘ�R@�D�ŀ��B���+�D	jI��g]��m.�HWXǱ{<j(pE�8��Aܠ�XUr1��؇��m��Rу���W��G��3�z"\\c-��J�d�S���x�"mi�`���HWWtN�/"�$�w�x�H����:�J4B��I��Q�j	80\>U�B%ѐ��Gս�j��%�)�E�b�٭�YJP꤯�����^6+=�؉@c�M��a�]��9��*�������6�7�� e���!�Y�:���m�*�UV_f�:�ُ�Xj�;V畕�[j��$@�B?k8���f�b��B�������0���-���6n?.����W9p����t�9\a�gg�ʷ�ׁ������/}�>4EA�B�V|W��S������ͯ�i�}������Q���4�JMf$V¹�O��<$�#fU��a��}�K-�kg��Y�s?�v��YVWп{m�X�� ���Ot����m�Ö���%/��Г9�,�ɳm�}��C��!�.�#�;b������B�v$��HC��׺��gۅV�0�2��[�Ǿ�Il�<�߯݆Ui��bmQ��x�G��Ŀ1��2bg���ů�������������Y.�	ƀH�����.xP
�O�ިh:�K@+ wO�g\"=��iD�w��gI��3��x%Q��j�V�3㢽qq�-�:U�)h}�ߤ[WL}��	���O��p�p�5��e�88��(�Һ��A�N6�CM�逛��j_ ��q��C64����+�F�?gX��*x�.����(�ؒ���.�)�Z �zi���v�ޑ�G�c4�	�E����ш��H�8�~��Y��K� ����T�2��"וg{�!�k �E����z@��������,qp��;�Zj؜����	��*47�k��c;a�U�T��-H�	l�-��L�U�{���̳��{����icq��s b`j����3���*�%�vh8UH�}���1j�b�r�����zk5��&�e4u�&��;<0�H���(��(��¯���q�����r�n�wہ)3�S:p��t���II����J�(���+`n2�9��P�I��3�JΡt{�Aצk�D��GW�����8a��QAQ�L������wN �N⫽�8d�S(-����0n�9.�n����/B�I��*���Ïz����M]���QG�D]�#��M�w`�"Ӭ�z᧦�|����/o4&�l���>-@~�V�����밴��+m;%%��8�i[����~��_�R�e�j��b\�΍}��a�t�ڎ���mb�֤�|´߷\�P,����"��7xDf�g���DLZ3��:a�gl��ڇ!@�ۏ���R*��X����fKriK^io�) {(f��̿�.��ճ�{�����[	3����ӠDD�C��ɿ����Yڤ���������0�>ޕ���zp�H�zP�_���dUFѷ���������(�_%KW��7V�)6�XNu�y>�UV��$�G ժ|l��(�-E��խc����dɠ4�RI'���+�J���	'ٕ����V������3^D�U���S��[X�8v�I��D׆(��P�	M�FwV��%������,4�`�$E';� ���M7�3���F"����/*�Ůhe[L��;��ԭ4I2�� p�
����a@,o|��j+-���J���ye0�Ѱmq�.�aI(}%�������68���kA�+�q�*�P>\�,��P�P�}H�AZ�k�p����0so�{�o8�m�&p����9%�B��4ց'֭`��b�;�ya��(�\0>sK�l�c&H�E����
#�
u�?/I�n��Z ��啰K^��l�T���Z���������K�m�ω*Ā)� 	B�v:!��Gn����SUl�"vG��G���*�'�a*�XF�3���l �FN|�C��>�Zz��>�0���@�Pڋ��=ld��N��W/�dJl	��xK�ejRN��hn�F۪|��K��Y�=�$>7��vD�����Xx�x�@��^�0j�G�K�oo#j�R�)�*�M��Ft9T���}d�Bjdu�8���z�I�Y�J�͊,�����.ĥ� �݂?�v�{���S��<���mN��f<d�����bF�Ax�՛����0�#�%��}�9=U^�6�v�Ś,�D�Qf��`���L5�!&��T�a&�A����K~�@��(.���+���K@|�Rcq,t��f�x�x��mt��B��g��O�IM����Q~�@��a��D�x3'KD�&����~�ƻU����d'�X�V%/��8y�� |2J7\iԛ(��h�p�;�Z��T�m��)���v��<F�ڶe��S�ji��9�H��-Έ����o�u�v�����ן����R�-���P7�:��U^�F.�s�s�-MwX�y#C��UF�{��D����RwBla��9f����2)��U^���ɛ�e0!�����W�,{���jm�u	ʽ�z	ƾ�nz�����}T� ��N�m��Qv��,({����ʝ,��h�����N���Q���v�X�z�֡����V]&+z陽�i�����lű۲�s��&79o�MV�>�Pن���?�(�!6Ό>��u߈��aGq_s8�ݢ�n�$�J�w%��N��$+�M�[ة-
u1��gQ�Y.��g= E�L�h�������ߦ���~Mq�ܣ)��*�'�7�z�zq�s�$�j��]�[)u�k��9�e�==H>�l;S�A�V/��t�y�%d[q I�5��mQ��k	�^�9�����
��hT������޺�GY����L�*�2�}S��n�S5v�m�a���%��i��K@6a�t<�`d������8�l��@7���G7?g�b���n�TܨP��{ ��J�ɨ�6�œz�����*ZG�R5c:'d�9��M�jE�9g��|����V����Az���M�;+gǐ��<��\w]5�+#�M�\ )e�@{�c�ʸaB7#!����^#&8����@�I?R{�.�aL�S�1Mi�5}d9u�1����%��FZ�)��^��%M�U(�	�3< s�i�ܖ!m��� k��}��ep�[�H�S�҉pz|G��Fڢ��w�{��Ţ��5B��'ѿ�|[�h{13d��2+%�3*˜+�����R�>Ů�-?-8K?�P�?����O�{s7���'�lz��P'Q�9@3�������L�Sj��W����\�1���$���wt:l��%Ⱦͮ9x��-g7�`������@��>hמ�������V�!L����`��1��ݔ�	���C��s�<iPB�:l(��ׄ��T�2Z�X}��q�a������Ve�{$S�(T���U�9��i$8ﻴ�<�}:2��m�բ�̸"}}N�R1���51¨Y�CP���Ge��/B�G��^�Qu#�W2���5���H^�0��:���&�.�����kM�~�+,e)�K�UB��i��U�ќ��%��x�
=��Ż�
��i?RT��19��Pu��u��gw����&D�BK��TV��s܏���Ad/�C,���c�e�́�GmXu"��t��}V����f�+t,����ƉͧW�����n(�YIsY�1j��J�.׾��o��w�:j�ډ��p�L1BTu��*�\�:8ҹ�n4w��MAg��u�iGχ�7�(�t`~�Yb?�p�<̓�%4*���4�́IYb�C^�덫�@�r��S�@��6SG��[��|�� ����(�}�՝N��F�kJ�`,%7b�d�Λ7�ӧ�N\O�Ŵ/��TID�hFO�M]�����\MWm=����4>��?!('�[Ns��ͯ���p�; ���>�����7�{��b��b�g�?!������]H�*�؃����y����9��ԂhB:~��Te�֒��:����'�RL�#���d{q;�'a���e�Nv��D��7�NØI�,7��Η-ҀK��ܞ���D�:!��;Ccz{��6��cPϗi�X78��@��UB�ZA`���W�����3l<2r�S|m�ޫ�,�����K��t&z���/��nC�=e�^̗6)*�m�G�`^�[:�c���HYW��Tg�����;�#я�S����|u[�jLqTe��g�j5qC��Sh�m��b�_�HM���S��my���#�*dE�:Ų�:0�7��\���Z8��QF����#N��b5�I�-�R_T;�:�Z �B2�T����i?�S_J���DA�Mo�{�嶛S��vR��D�.�4�\�����B>� �T�I�aKQa�P�u4�>-E���^G��ͲU7�Y6,�QK�ș!�}U��L�jaJy�� ��Ri��@7+vg�`=�xaΦ��/�c��V�������N�����Gܸ,���"�ξ���`2JP���i��IN��m��Q�@���#���&�=%$8�(x��m����W�7�}�'��9bֽ�iʯJ�b��ma.�P��N�'��`�>�]7�v���c9T�M�/O�g�j�|��P�
�4h��1m��ߎk�S�m�#3(�B]#A=��W/�*�x<�M%�-K(�6M,y��͕�s��&zCj�����Kҙ��%��W����s��w ���S�͹�l˺.+Z�[��Ӈ�'�������{�h�B|F�g��C��f�c_-M8�r�ǀ1�/��s��&��\bn�Φ1��Τ���v׸H�zsd��v�pQ[Rv%�z[IG����z��E蹂)y����}��c
����� ���R�B^�=�������	��g������Y��/_-��f�]]�ܽs�܃MMs��󓎝%�$^;����x[b3���9��?0ե�2����o�(^6�q�;���3Rj�C����@�)�.J(�u�%�t��o4$E��y��	���̞��#���T�.�b��b�rw���	N�@�t�E�&�[�*�wW�?��wu�ц"w�SL�x���6��J�T��
l~ޚ�����9:a"E6b�眿�����Y��
���ɯ|-�ֆ����j�I�G4�s
��\\źPnЙ=Lc!'��zG��=T[��m�)z_��%�`m48��ns[T$�<)#.!��L�6&8)�M�(`�{�Lw��&+9_P<9�?%��J�v�JY�-��7굪2$D�߀8i�(�E\J��܉���}~�k����TR�O(q*�ݫ�)�>�� e6��s]�S)H����\�a�uR��5��&#�^��A~Nk@��W����
�NU�V��ż�!�l���ܦ�vV�h���o��xV=R�^b.����;�-��ڒbҺz�u�mϣ�^�4��$���ŵ�v�dߎy�'�K�dY[S����&j�wmE�@�Sl�@���k��x�$`��UD.P�^^�/R�YTè�1���;���v���Ыŷ!D>%9�&*�nAsiu,9X�Uo���_�[1��M�������*7d8�PO�8mq��˲h�ѿ4�0�x���^Y�<�ZQ�e�q��U�Ht���X`�Q����r�5���P��2`hg��6M�k���y���o�Q+F��	�.�`A!'a�l5���J�D�6v�Et�.��]wu>�6���'�Rh�Z�g��~�:��qCm�� Dw����#�I@ʼ�fh��C��_�^��eHep�b-����7��s_�ϟDJڔ4����muX٪�@��po�fbR��|<�W���/z����|m��ӟ%��s�h��Uh%1��ui$�g4t�ݡ-�*aD�H,���-n��{�.�2s�65��86�9�_(��֥��`	����@F\�_�/LWÐȳAx�b�\5j��~�~p��c]���Oߐ�E�ȋTE�<��&�/P -K0�bl��i������[���*$z�'����b3t�;�������;7��`̿��V��ܞ �G��scf��|�ܳVa�oW�ZX�O��a�i��(�� /Dt�3�e�v��Wa���u`C����~�y���P�[j�IInj��ј9�'�ΐ������R� �M`�������TT�/�D:Q�lb� ?��n�P�`�ذ�@'E�|WE�P�j��9�=�^�}:U�e�,���-�Dw�\��sր-�G��Bv%(m�1uc�X�7<��|#�6�4�V�m�{W\"�RJ�-�5��Z̮��%�E��ʥL�|Z�P�il���
��k������'�	)b�%���uo��C`�B%*���5�W�-��&�� JYK2�A����},�[;��'ޢH�o��~�ve���Bx����ͩ���7��:�r�R�n�7�������텻��D�]���C$�=f��
�yPRJ����7	�mҨF�2����^GY-���_�fj�-B t��W�r�1�m�T=�Cy'U��N��� J�nʕ�:Mx�Ӈ�n�c�\U�ۿ�%L*V�-�k���8��[�8V��a�S;���K�[�?=F���� &�K����V�c:GG�:�����[ŌW�e>�b��\��-���3��u�"�Rh�u�]�k<��hਞ;�ڳ'�,/1}�����Z��<;k��%��
����!m�?bE�vgvU����h9�-ct���W̝Z�!s{��֔��M�	�J�ԡ!�3 ��Ӕ���X쩉��`�lT���o��$	�*�Bh��V$�r�ҵ���IT��0[.�iA�>��>�<sB��.��Ʃ�k_��|&��̀��t���>��҉��ҁ%��N� @�������m3�7$h59:`C��Bߦ�b�������9Zz9���f��",�N[������Q��4�*Xr�\�O:��ڟHf�)�dk�A"�"���4̸)��;�B��K�'��t��Q*vH�����%V��6>��e���ܨ�ֿ�t�=t�@��p�a�:ף����|X r�dj�W�@N2�s����Y���U5g;1�*�*i^t��`��;#�k�����c���XQ�.��[ǆNj�v6�EgS�ggT�k���2��j�%s׻��)����g/�%W��S��S��<Jр��s_/q��8YU�-�	 �Wm0�	oU�C����H�*Dj֊�8� �1���V$`�~$t�-���7ErkӨCiZ�rMxg����B�X����'WKmƈ��[P�k,"i~��4D"�*���0[�ƪ��p��~��~o����=J�R	-gCH��(�����"�$U���t�U�;�[@|�ùR�G�=�m'?�:�5�� �X�A&L�y�5�vH�$��t�Yi��X��FHC��&BeK�g�;�|�ӕ�mY�w�Jk	k\�cX���܎�p��0 �� �(�d���L�X}"�6��pM2lII_���
�D�����şt�ժ3pه(�	)4��%H��m���f򫷝S	��wm�THt�J���]6H����h�k���U�q��2�ι�_��E�t��b��n�pn3;x����p�>O4�!'=	9�ɲ�r����.��[�����l"��r�&x��g���J�����J�i�$���-��i� [�N��OY|q+%L��� nA�,�N��:a��E�O���ü����W�<�Ē���� y���+<�.��������U~e���� Yޮ
7�d��E���OY^C��\�B�jDBY�n{�t����g�J�+=�� ��ful�6js�^��h�NMlv��K�l�0�d�5ƕ��̕�4�bN.R���OG��7�Keܔ��x�"�yA�e����d[���s���7�1G����%
�5�?:q_V*���7� ��#���h�R���� ��-4����T%t9�E�ז�=K��}~������� �J7o�5��n6$#R�ǋ6�R�R�.X�lm�,C�x��g�i�(���s�d��e&Au��{5���e�,�v���XI~^�/����&c��*�S��a�KԀj8?;��ř��MV��y�?�a��oTF��)j8|���n��~�ax�p�>vKCT��6��G�6��iN
?�Óe����v��'�0X�"�2��E���L�lD���=�an�t(���֚π��A��|2e^35������;[�������#Z\l�\$�ˣ_i�G��m�q��幄#�k!Dnp�r��$J�8=ٻ��\�2�Ȯ �u��X/�����FB���)\���$ݙ��)DUM	�K:v�z��ծ,����q������3����q��8_`����'������{&��%�N�$�s #��8K��\vqĎ�+��St��\�^ӗ�B��:ٶ�i2���|�*�8I�i�:�HnE�f������3�6�G٭{D��.#�h'1�'8����R$�����*�1rēF�R���Fh�>���2����w_Pϩ��]�xC���+�̀���=��Ҳ�γ��6A��oG������~����m_�`c�R����(
�T B:�L%N~�6}�;\
�����G��
���5��t��=�>O�Dh�@���m�v>65�Sݭ����B�.�׊�R��"L�S�s6�ء+��ZF�~����?��~�=���2*��AMڠ*���niU��}��W�W�	�39J"\�ߏF�x��]#�U8?��55�{�kI�3܏���BE��!��l$�yN���(lD���c�
wōa��4v�73�k�+j�oA�`��Z~y����v���������jD��g��<�Y�7�ࢄ��i=1�
tp�#���G�������2I]^�����LCp��'�6)�6�o<��"�0�|.LMnvm��`��@��4i<]0���e�f2�\>����o��ϴc�*>~����e���8���ˤ6���h�]�#�{��I$�6�Vd{�3a��8?쀪��\j_[�����R�]���C� {�Ж���S����ZL�z� ,���v,[� ��?}���L�~�[�l���Hs��N�5�ƏV�����A�^ۨ���-��d�S�r\�[4t�W����ɕ��\0�w�;�Q��c{���f*Y���MK���8���z�REAL'����F���,���/��Jb��H�6;YҠ�$P�/�qG�'m��K?�2�eʚ�ϔk0�""e�M{��B�q����:�z�:�&�7�_��d�*�J�2�n�tE޽��J�lmT1a�K!���#c�l�%D�|���R[�ݸcjx	O��܂٢�iVq���B�c��5OcQn�J"�:��668��,��lɄ偽��r@� R��iz���c}$�) ����%��5��i�
��tq�2a�(��@�Aܥ�Pݠ�����݄i @;5z���;ٶ7IW����r!N(ot�R���7��r�m��4҃6-�x��Y��͢�6!�Դ�i�$�� w��P�3��m����R �ӷbd�$�k���Ա%����"�f��(�x����;m��� i�n@�!7ƠSީ�hL�{�L�]z<�*�����r<oh�b��]�~��F�6A	�wu��U�> ,���X��3�Q8�O�-����T}���nk��ϛ �����K�
��	]rKf��5fؓm�)�/1�3�`��ĄzK�J*�p��g���1�o0���3���#�� >��va��n�)()��>��N%����� ���F�y?3E�j����5�*>h�F� ��)������2�G�ԑ�N[m$0'�����o/�J�Ķf��蟨O�����ܕ]܎�r���vH��������<#p�-��)_v��(,Wn9�T(:��P�O��y6��v�/Ji|�UL|͌r;W�`��[��i����y�tpp�]g��j�z/�r���<dOpw��}�����ҳ& ��*:�<?L����ɼv}�e������2�MA����������֓&� �����N��_٬`%Ѥ��ŀ��E{�vy]LМ��TFjR�N�Ƥc�L�O U~��Cq�=�e�9l��)���ż���%N��"����0��Y��D�0�p�:���,B���Sn���h�i��|���$������癉��yP�n� ��R�l庄�>�qxm���D�f��P����m]l�w`Y-Xx�|��x��+�f~��G���] :���~���U��T�8 Lt�l�/,��+)�v܂kִ�EA��/Չ�⧪��֛'��'[}	7�Q���-HH/W������>F��K�&CY�D�,VU�ψ�HZpS��'��Ě����2�� E�,��&>��N�d;����Tw �D�I�[ÊNb�dKa�&�W? ��IZ}�/"
�-�m�
�f���[��,I9�,�>z��↫]d���	Pb&zm6�^�u�]ZN�d���,rl�J�ѧ�JlZ��(�����^�|� ��`lѐ.�͂Ɩ�%$��XHyy�������N��"���=$D��9�{o�~�����X���uGwt��+��s6<:��+	z-�v�X� ]��ʃ%�>b��bd�y�i��G;+	�)���cqs��89��ə�ͪ��H�+�;C>�sZ�B�@&�)U�hEC�T����q0s	Ж{��6��]���3�NH	K�����Q�=���XA����	�U�z��0(n]%��d$�$j���͑B�o���F�1�"15�8u\��^b��wC������.����f�����u�Z$w���\�;f!?v7C��F,ۀ��ꏟx���!2�3o�-�N\�=�M��"�C����'c
r/c�~�Л*,�c�[[9����+�@]2�[t��N=�� �=>�p'�' H��G[����pS[e�w���m���	Nor˔�(��5����}����t/d��CF/��<�5�T7r������hoN�|�ǒ	��v����	X��igu�����������LG����j�8��ڠ��6,���~��K�7Ж��Fl��)��[�Fx �>���j�^�ƂL������<�[�\^��I(�b�
(��v��F�Ք��<�h��\)�O�l�A��X3]�DS�#/T���Y�ٖ�.B2��7>�ǮIxU<�h�hw�-[�*�Z� ��p`�"�P�����=������2�h���/��sk�������3U�}Yԫ眽��)UT�?�l�H�a1V�}��vE���٫^NGO���a��a�j��J}j�C�I�K�����띊�������4��^9y�ɯ*U\�f?��}f���2��Q�_����_'(���O,Q��Z�yg=Q��CY��Д��t貢�Jl8��wI�|�!��9+��]��Ǹ	t=�:��l-��5�{�H#t;�|�������#S�NP���:����t�Z-5F���i��M����Nnnԫ$2���� !�iXk�榖9YM`X'��w��i�SޠZ\��̡Ս�^�+��d?���YS����ZyC�1(ǖ�}O�aX�Sl݁>��j���u5_�aWFۙ8�6�(�lG��[��!�C{`g����9�"�UA­�5+x3\?J�]Z㠙�p�P��w봞�E^1)���t�2�d��3v���T�G��
JI�v:"�#"�Y�#)=a��¤��u}�v�l��B�*�C!�����q��Or��o���	�xc��p��4�#9��y*����z�=>rHC��)�5���a�Q��^���H;B�0d|^L8��Ww�R��fh��?���'Ln霞y CBJ�X��g�b�S��p2u�:��==�Բ���uк)���ϡ]O�K���a7���u��9�����/~����^���-=�pn<���2ESݵi�O^�䚗���d����I̜)��v�xጃ���d�k�:lu��Rж�?��-�o�\{w�ӌ8� ~B�ՎAŃ�$�᧻�+�,�`*�v"�!uf�>�J�Sh̎8�_m�C�����'�T��>��������(t�KHc�I��bGא�en}C�bN2ew;d9�،g�V7�ߝ�<�Bڑw�8�s��.���w��}��^=��9�R~+�ߛmڲ�|��pp�����D���x{�����)��u҉('IX�XxY�4+��	G�D�5�P��}z��A��Ew�r]��*u�9�1x4�I�1�A��e_��}��I�s��D8].�٭@�'&�> V��AЏyF�9;�7�r����C;���t-mʨn8�0���*�dg�Zd�1��!�&|�NL�V�-����LݸEd2�f	;J�8'(	̚�^�ҏ���2�j�-�K�\����N
t���=� E�����@�R��p��]������|t#zt�!��yPRJ�:�`7z/�}�|��Gm�W�>K�o ܃&��9o�$����QK��~��N�:Hc�ۉ0Sz��+O_�tJN�Q�^Eͻ�(@��4I��>GXy�,��GP��/B=\�����6��!E�AҖ����Um)��9��#!�/�j�e�{�$�1=��Cq�<-�*Wy���Ukb�+*�(��!�˸&T���.^���<��xd'2G�$CY�!(��K�a�N�
V��H��b�5�߳)s&E��sz8VD jH�lE�<wH�m<���)��t;j�=��uK&����tN1ܓ
ŕ����{��&W�5
^!}����!�0N��EbE�g��"�&K�&��kR�=l�
�����%3׃�~�$2beyE:�����n�I������Z	C7��]x�;�)��.��r��CVM�������IM
U6�4�T�]D,�*��֮lR`�7�<����k^�7��\n�QH�')@ӧ�*�4��Y`n����㇈�z�^�~�
n�[�f̜�_�is/��$�1	 ��hLA�:t�KbC�g��5M"6F�h�?k�b�YmhJ�o��Lߔp�����5)[D�������7����
p���gC"D�H���v�Q>0 w��i;S�-KC���6��6����2W~��ㄠ�y��%J��6U u�_�[v?Tf�??��)��(�ۃ�W�6��>q���a�˂:j_vσ�+a½����CI`�v���d�Q��(w��y'�4ʒ����#�ؒ����:V�������`�^^
k�f�`U��Vz߀�8uʟ�Ѩ�0zmSY�Cp��r�Z�Z��!!�g�]IJ�.�?�چ�W"a ���E�?�cq\jƲ�Vr�K�/�br��W|]Y�SrRxU����^r�y)r���fi�/.�/�T���%@w���rA2 }>�;Zеq/͇9g�K#k�VM����V%�Rc�ز8���S���U������IQ���r�_Џ9g�i�B��`�Zi3蒢�jIX��*��[#�i�LD�`��h�4r��H��Ӭ���;ۿ�!��Kn�Kشӆ��{ܻ�3q{)r�����

!V9q��#�rZ@G6*�B�v�%��j�3�K�P�ay��A�㯝=]�>���BH�u�#\dv��4I�r�c�t�KZ&d꥜ӲO�����A�۫˘4���=!���pT���DD��'�uuy�98���A�)2೨�Ȼ�ŋ�I�(��BVrM��w��{P>Rꋤk���4 ��N������Mض�`��ʽ5T���-)�/�ב�5z:�&f=Dg-��y�j�LV����8�����#sqՊݟ0�S�g:@�{}!�.A��v7�����צ��\�
��B!UL�zDs}���vIz�{r�dp%�^��kQ����k"ڕPߋD C��}��{����D?�w���vn��u�LEX����$ep���R��#%b]9�14gz��-W��P��lc	�L��ռ�6DV���ؤoiΤu<�>0\���ۍ\�ņ��_�yj��YO��.���ݕ�2�٩%t�8��c�xҚ-ܔ�22-�i��$/�r���]����3�{�bf���	A`��9�$����Gq-��f屔�!N޳3�����ax@i8=ꝩ5���-��ӭ��H��q�yr�dJ����t�[���^Sh_�i+G����.�
O��������v��R�W���!���"��&����7H`�+wh�O4a�&��� cڑ_��e||½��������u�{̆��$�|������b��/�� �9��0e��������L|��1c��I�HL�L�n ��Y ����0Pѵ-Zx��3��8��CLkn8:�0W�ty��{[��i���8�`PΦ��3�����fe��Ҽn�J���Ѭ��������$�E�Z���8S��
�j��Xk6�ܒ&�s��]Ih���y��M>�^#[IO��T^N�Z��z�=��)Pʀ��!�`�Z�DC?��c��su��RS`�vԸ}�u��U����]ꐂ9��o��|����w5�31�f��e�Z���"�[Y=��������t�H��J(D�!d9�+�$��~��`�iXP\F�IXL�<�=^��+�����I�cWӆ&ˢL��������E 
��`J�
}ˏy���Q03��ڊEo1QLJ�l�	.�VE_������Z�H�T��֎JR�"�C�"0"&Z�ݙ�
��aj�*�B���G��p}����{�9�¨���BG:O�5*(��Xm@�;���
:�-ë�\�e*�u�z�C�jJ��hѯ��c�Ȃff���'&�6����&���Rሎ�e^1(��\����.��Вj��*g`�˖�-.����W��v�饓K���(�b1[�!��VdV��N���~:�p�
�$�
�8�þ@j�-���>b�*��K"�pC�G���n�o�O_��t�H�u�4�s���Uә�o�쏕�����M���~_ʦ̌�T.~BW@��sƹ$��!v��=�~���ă1��t$U�ӆ^�q��t�b.�.�>�ghM��K_B݃���э?"%�K�<V�PAaS��)����b\�Ls�'��XZL�<�T�J^���y��'R����0���e�1�Rp��nHHrC�(�A��0ѿ�p����[�mP�|�ܰ��YU�lW}Q��(�%1�4�Ċ ��Z�4�����cmO�p��A	R�Z' �#ufW'�n�m{�{0pZ��`�/�xRK{���ܶ�~�h���}�`�;7����&�p��c�G�i(�ch�1-F�t�L�X (C�ٟ$z,ԓg���9��x^�of�bP@n~Kp��S���=�6���"��h�)-�m�P�{X�N:U(�t5���)��q$� m3�ۺTJ;�Ԙ)��BG5(��Q e�Vv ��|���!� ֎#�Œ������e{�v"��!�-�C�m� �/l�D%��2�D]v�L yDx���1�v�l75�W�����N<o��3�?�0�[&^9�� �E_��s�����5�x�~����WW�6���CL�d�i��5�_��쾤���O��_�n�Z�����#����w5�6��4Z� �-OK��wve��E߷~R�˝�nE��τ�W��-ɵp��� {�e�9�M��($�%�bh��)@�^I���� m�	�a�L�^ K����6��a�o�^��S��+j�hlRe�>�$sHQ%0L��ܿ��E^�TMP���a���3�����!Pӯ`vo�ſ�/{�� g�x�&u�6�d��@��Uh0S'M@Y[M�;!�ߎ
|z
�y�yq��_k+]���ֻ��W�T�r�����f���Y��E>m�$��Β4E2����i�g���)��抆3�8٪}�����h��n�}v1�۾��U�r}�cv[t]a�4,Ǎ��S.�T�́��4�r��l���$?�!��Ab�	�Y�[�y]�T�4J8�]�6��v�|�����J�	Ȼ2���HS���:L` �37x��@�����rjX��wc�{�ne�{w)%pr����T�Y�N���J�}�-��׉b�����?舻�#�O�O��8DBv��9��̯)�Fh��3q��B����d�I��L���YےƋ)�������1Z'X\���4u)c�d�y�Gp�Ғ&IVn����:��#a�b�3����:�C�~lx�D�]¤�RGV:�k}�>e�
��V-�h�@�ۡ��S�,/�!ҁնBi��~�X?Mނ�(���{}3��FO6��TR���OR��/Ŏ!��'�]O��d����Zܪ������Y�m� ���{8"5������P�����촖Xu6a���r�3&��,k���>d�re@��;ى���߆:a�T������y����T�w�!�=���c��!D�"�Ȭ~^�thN?�;f�;�D!P\�«xF�;��P�$��K8"�ñ�Eu�Xd.�Pn
�g��N�Z�+�d*��`��\�*�����_t�5#�=���"H�z��v�/m��Ʈ�tx��9c�!L���5Yy�6�.���>����>����C�1���_�G[+$f�Pm�ɕ_*Pk�3B�wI�vc����m?4f�Bh�U�`�' �^�@-�YH�������q}��(��K�V�j�z���h����E�ݥ��S�7��{q���c6Ji/X�u�%A-uifU�p����/�u��8�zrH�x��8�d�{�b����<o+�bϤ���ٮ;��ձ!�*r!��ҕh��ma�u�&���O��&v'	g�;Ī>S  _����VJ��|���3��KF��Ec�HԖ��w�=�����d�fz��1���>��U�ׄ����/$)��tQ�{v����֓3���Ӧf���"�^�6��:���Q��=��Z5�� �7�]��s*�O���/�
��d�4�\It�_��V�w� ��ɛz�]�E�h6'�Q	�y��e�����l�h�(T]`�eXzw��?燣ҳ^�k�X����B:5��	UO�<q��9�]�� ��|*�x�T_Ը��6]�y�IL�y����F�O����4�=DT;aA\��������54���p�O�تA!�|�=u�,�v縘�-������j�V�c���j5��	ߟ�G�#���*FҐ��Г8o�ν�����^�lo_M�sɤ ��_e����6�o�
f�z�q���1���p����)��.���?��X�{_��f���Hl�w��࢐�����h��ǚ�Ju��h��_��3���9z��S�\D�V�v���Y�K'^Tѯ�Z@XV��m��lr�D�ӊ�7���H��ԛ���T��|�Iʮl$8���ɣ�$�j2pZ���	��/�<�.'�"�̴�S/)���7?�6� ����ն#o{y�vψI�5I�(�����G�~Z[�:	��@d?jvm�[�~��� zJ��'��X��y�c%ke컱�{�_P�������
�/�h�b��c�b[��_!	F*+�r}��Y�A�}D�m���.�������wOG�0�P�h-aL�
�%�4b��@igB�����]��h�4]폰8Ir��.A�&��r�o/,8��j����L��b���eʐ�����33^�a���4���Zx6΁U�&�.}�M'��J���'E��a���U�1Y�5.�������V|�Wng5j�� �Z@ظ#>���D�}?v
���&Mmb�1��O����3H���U��G�����?r�X��.5��2u�"�հ�7(^��?ǂ��{Dd�J�7vm����a�m㟾��*T�a=b����K*0�'<,�@��0���ɘ��+�0%e��n3�>M�1%��;<I�ꍘ�?���MJ�v�;wY :�R�Т��|�@�80u��>͋DD��߀A����� �V�[�m4�4�/�+���6ǘ����="��J�=%�5����sƜ�]#]�d3d�?�d���wH���(Y�R���"K]Ò��������3"�|{�[�fWV�?����e���H�A@c^��	rH�pgn�,���c췩@���NC�\ ��Ԧq4#M����<�Fʾ�C�.�8��L��O����*��	�bv=���������7�i�j�F�_z������itGbVl@K�P��ܲ��!�J�y�!�֒�P�Ur���R�s���xs2Oė��1��W��(���%ҩ�+iO�g0f4��f�G�u���X`����#s�.�X�۔�^O�@���_���ͣ�ؐC]���9�p�؟O_��N.�0���&B!�|�i���"6K����!mY7��E�`�g�;���<�8Jɚ�0��+	[��*z[d4xI��±d�'�:�rO�ɣ/��a�]��K���8C� _���w�A�
I��Uo �0i��>��"j��^qPc�J��SX]���H������rb�_g�VN�~��e�d��誓#r�2��=���b �v��s_����[9Ot���Ҳ}�?�̢��(�VD��ۘE���q�30�2�D'���7h�ݢ��sw���_�!�J�{I����!�Y����o{��j�l3��1�x�r$��ش���XW�?
�R�v�x�p����FF�����R�/ܔEq%������-lr����D�X
�<$Io ���$�~	��~Oxs7)z�6 �לoVϽ ��AE<�� \��aK$�Ŧ��8_�P.�#��X��m���T��'�t���5R2��z&+s��+��CJ��+Ã9��l�YA�m2	�qi]�}~�-U�#���98�'�yf2�:�u/Mq@��s�yq �7�v�xS�lN�M�?�'�PB{�{o���s�!��^'nhOdKpF�5�*~��˖r�L\?���l���2�BI��ό��t�1��ٰ�70t�z�z�J����T:�AC�i��3���+��r�IhQg�{����� ]��X�=����O!d�CyC�"K�F�Q�-�&}��]�aQ�$�?���%~��呴dV��˃�HXݭ\1��:��a�GY:��3δw�bI�-K?j�� !�WMo{�[/�7)�^�G$�����2{����"=\���1�^ٞs�M�du�f!A�D\?'Wx`�I ��[���@��-��6�	��4�L�8:"�qtF?�� D��m�p��;�Tb�%^�G4PԦGSSǄ�5�s���5O/���-���~���S�57�ɍ �U*:�q��MY�%���S��#��� ��L��[t��i\��^��.���e7����	����	u�g� �����^bZc`�쪎{u������M'��[�zgž�?��O����D��.�ӻ+H�J�س�Eb�����tےQZ\���	�Z�C�����*�#�E�gJ�1Ќ��|n>2c�q�) ,,b"bf*D3��Ғ}��O�ڡ��3�ƫ�ب*H˧���^���h����Ks�m�=��Dqߜ����j��8�<�k����f��Sfã�7��'��J�U��ӂ	m�7dQ:���*�/.�X�W�XK<)ڰ7�YM���d"hg��jI[���"\P?A�]�l����X��5�M���vd�b�w\,����>�.�K܀~;�,���*;ٍ��Dq����|H�+-��/R��H-\cjU����@�˘�a�9�ƑA����ݍw�]J_E��\&O��L8�!�����!���[���ն��y�������H2��F������ê^�˯��=Q'Ι�q��B�`ȋ�U�o�n,}A�Ap��x�{�XnT|�v�|o>�/��ɭ��N��}e�2J��	׈W-��S�|��g�g�Ctn=3����Z���z3p�g���v���Y��9N��Ӛ����r�5�J�����v~�R�Tm�W���Ō�&��g�X#�mg.����A��=w�gM�Aq�*�q���2I�3l���04��_��݉� �����7�m�]=���O���M΃��t��;w�t�z��\^|�P`1���O]���»�������һv*��t��h�6�z��<k�q!���<�ؕؖJ�	6dX�ݙdG*C����$	���E��<կ���/v�\�5�k�3��!uݨ�>�gG`�Z�eF�~��[X��3Ƒ�o/-���m��U,�a��d9p)<��X��=.wH�l��D�W7DΡwꁚO.^R����R���l��1ꍸs��� յ���b��^�B��^\-J¸G���j3��c(��&��)X �6�`I+=���2�
�Ѻ%靖�N���S{��v~ �%������s��^3�)�e�`ӷ;FcR4N� ����Ȼ����<��G�)����8�3B.��� v�c��갟\�E�taĨg�'��y�n�����VJ�Ԃ�����b'��.e�o�%ku��;��#�3D,4�7�1���;�C��WA�gy㳤X&� ��/�Sf>���3�2����C,{ �Hh-�&�;C{�5x�������4�'��!|
�_&:4����� �,*�N��D!"��2��E�E|7�0U9/�0��ݮp�E��[�#�Լ� *KM:N�⧓P&C�+І��g�#Ѥ[��߄<aC�xQ��3�m��l�z��g����BjHǅ]Jef�$i���4d~����0��1r��2��=޳縷��le9J�I�hfx+2���	Zͱ�h)|�kF�vd��E>R5<gN��W\�K� E6��F]�:��J�m=2�~���x�%eʍ˟�e�)����C�� 7V�K??f��2m���C�D��iσ��X�u��$EH�$�l�3^�=rp�ҏ"�����u<eϪ���(�=��~���f���Q.B���MD�z̭ZF�y@�3?$��7���#|%s%Lw#���U �������@�y/&ze��\�C�p87�-?��(���#�j4�X���ӥ�y�d��x	�1�^�ʀ�Ա:9�?�u�yv8��
���8���B[^Z� ����p�T�D�"0F�*���)���-,,���f�g����{w`��eER �h��N�o�F��@	<*�o8Uh �l��2i����pAV��� iu����{�5l�:*��߄����ѓ��àwg�*Z�݅)י�q|V���'�9�V�V��3 CP�Z��篂/�M��V����$=+�����_ri�
���|,�O����Xs�r8Q9t�}��B�g��vD�eE��VRN�*|h�^ȏ�=�Jz\ʡ���D�E�.���2�
�Q�Cۃo�Y�K1ݺ�l?ȝ�.9�|�,ރ���y���"5N� ��nHb�r��+l7s`���T�O�;�D(G6�ܞ���O,�c�KO��D�5�ڷ���8�e_韱��<"3c�5nux�P@����~7��!D�C�G�&�Q11� #�P�Sř��zh�NnY�Ү;Fk���z$x�>0S捥�� �23��%?�j%ua��
j+ccץXun�*��s�lF��`���[d�Z�6�w?ui��B�*^�Ppl&���{'��O��D3����I��eޒ��F���<p��+�f��p�ǹ�� r�zn+��j�vgd� �\0�CŅR�Q�\��Ìٕ�|O�.�R�5L 1z��?�.�E�M��}f��k�HӮ�b�k]���s"g����6
ڐ�鯨w���蘈���zj1�҇فX���刀�/��$��H˭�ͥ5�:���h4� �$�e��_��?*r�W;P�A��T��x�)ն��U{~��[%���[�a<����s +�C�-9-<�oR.����I����p
6�n��7����8�\����k���Js�d-H�pu��V-/�T���M�~쯃q������3ȇ�.��p���&YȄ8]׼��ڬ��z��'���F��f���}�^�m��	L��)�L���D��_�>�޾�LG�M ���5nL�o%��H� �m��կγ�k�E驊q>*��s�NV�S��sB:h;Ӽ��DT�ܳ�TG���eM_���� �@9�剈�Y��2�f��G��]���{��k���?>[:\�cD�~���:�,`]��4�IH���&*��Y!w샧=�p�
]��sMn�:�3|�[$t�D��S����D[�4L67S��+@0\A6����"�O��{F h�ބ-�&���+��nɧ��4����5���ʔ�C�gm��1=5Xi��P�R��� ��UR�6�@���r��Nzc���]������j>���;����%:��+��A[�R���Zx&���u��>����a����M̾ ���(����3�������Ld�*�A�dV������LfV���K,�I��mg���D �6��yOn�޿�CԜf^�]���B?��;���Vd'_H@��+%u�K5�ܳ��;8� �ͷb���ӲfS��Q�/�M���d����UQ�,i+b��)i��ǀ	9�� [&�E���¤�X5%VE?��:S���.�E�FRN�X��6pc6�Z̲���4����~��Y3�볿'�������#���7�I�㯂�������(RV㭄������>j6�K�02�}�X��(�T/~r��%�$�S�N��v�e;�}���ͽ�x^�t@pbtāϲF�.jh���?Cv����%�Ǩ7��Aq���`79�N^�Ă�����S��̔_6r��ߌd���5�u쉉�'
����;�[��+=�J,O%dap�K���o��8����/���s(?����!�[I"N�$7��zR���i.m�St%��-lY�Ln�R{P`7?��:�T�P4����5�̤ǳ;  )��P0g�*� �n�S��C��Lra�،�ABcK�Y$p[~w�1�ߣ^�e�EZ�zb�y�zg��d�a[�\G�%\�9W��u����9�x��=W�|�B��ψ����ﵞ�Vb.�^��,@�E��qk�������Ơ�c O	�LSNs��n�:���S��U�t��#2,P�|w�=��f|��Xv�"T�c������z��8 �聠�GO͵Hߏ Nj}I n�ħ�km����NK�פ-��9/��6FFӹ���� �� ��{����U?�GJN��\��"!⥊n�
�������I�����œZx��E�RR�'�kd+�f`_S��"��9�:6�ɐU�M��M�){閴Tb�/��%���\�)����m����e8K��I#3R	��j~K0��|���N��
��'AƁ��[��Q����t��;�[�sOKXN:˯l�c4����4@t�/��6�ϩ�}��N�P���楦@�k�4U4E���c)��%�@��-i��/���2A/�Q�%l�hP�@�G�������p������ͤ��(k?2�����������`�rM�P+��|��5Kz4�g�S��N���-�n����tfc���s��H�3qv\�|�Jb�6���a���*�ר��O%�5lD5!>!k���ܷnά�{J��C������_O��J�F�k\5	G�L�	L�ɏ��� �1�"�3�.XbA�H�D ����^��SH�>�|���	���#��P|~@P�)2�h��Tȏ�)UXtrfy�roL�!X ��Z%&o��l�F#䴃��3�.����A���N�_��ֆ�;�-(���,Ǐ'5�|O���f���w�����sB~7-|�9b�2�D7bA������ׄb��|�opCU?;,Ɗ4M�b����\M�g�Wt�݄��x�)�Z�������'[#��tZΆ��ayI>���l�g[�@�u��4�9'̟�O�����)6�����d�,g�������ݦ���-n:CgA��.�f�tY������''�U�P$RL4��ؐcg�����O�{���pQ<X�QzD'���qˊ�:�?���\��+"+�.@P�T~u����@e>�y�Ɛ-ؘ"����>Ó��I�b".H����#�\G�ħN��3R)��7 RY$Ldik�J���s^�:������S��ks/�'��!kb-�&�k��ڭ*�)Mɕj���ֲ��xm��י��[']�[�[	�
h���&���i �����5�ɠ�}�eh > �s���I13��[��aA��U&��0P����	�����n��2`�#e��FL_q��e�"�����1bz�B�X7��p��U%ơ�q��4կ�O��6l�<��J�e�[��q���J�ۂ����(��Qu�Ai+��~^���U��ga��<v�o-�� >�C��^��>Ir��`��	�wr�n�'iId�=9��U0OYJ������L׽���4�6<ԉ�<Aˀ�?���~[����"�Ş¬�5v+�=�"��t�{:�//�rm�<\��[Q�d��Y�	�>�շ�2�����3H���n��|c�R'��$L��u4i >�-��@���i����s?EV�u.ޙt�RLV�?�NM�O�4�HX0�59�!c-���:�؄��
���^M_#s&S��,Ĕ�瘨Ԡ��m�������_|�1�fr��^ȌDbCJ�Y��{}j��ٺYT��c�8�Z�&�w��rh���O����:$��IM�z�EO ���bO�3j�EI9�<�h���;��R��#;�Xѩ��+��M�7�ɶZ"�q&Ч�J�r�/|�PL� �O'o
��!��)��PP��ɠZ`���?�I=��9�b��{��;�˛$�pk{[D�|�����ܒc�)��ƍ����u0ړ�s�|դ��T�~y^��g)Q@���U��L%�ґ	{�=<��p5#K0�o��3P�U5��v%G7OGV֤���M�9#�ŵ��"����zN�㩇!�*ep���R˞�t�G$�k�y_��F�ns]�Y6]�_�z�Y�$�#�k61��c��D��Y��3Z0`l@��aͽi�J4C��7���6ug���#�b���n��^!4��KAGo=���BV�-����aOi��������H�^@�I*��u��F�]��Q����2�"�^�3U��a�9N�	j�F������`X�U��c�C��-s��Q�X�/��ʄ0�R��-�F���D�cA?��3�\~��:����A�Б���/����<�M�Zg*m^یr��*�\�bJ��ӻu�m����L��.��(t�`̔g�D1��;�Y߳+:"ju��i�7�y ��2M��ܡ���ò
�'k}u����
��؉�( 5/Q{S�z$�c����1� �܂�����r�D����Դ��TH:�(��C�_�ӧ�`��F#�8�C�@�Q*.WLn��MӔ�|�'Ǹa�>+���B�ɤ@�ҏ�6y{�!9n�@�"`�˧�;��ۼR��B��v։ͥ#/��ϝ3^�k�g�U��i����5\����}�G����"CI�͌Yʻ�QA�ڗ��fH�l�5_���� �̈́����P:c�����!b�6:l����D���TQ��@Z��t�Q�_P�7�����QoPޞ�==]~�����V4�2�Ӟ�0o��`C��c>��c�t�}�����.X�j4�D�s;)���K)z'��'od[;��ov����to��p9�~��Ҍt�o7�,q;�`�ukam!aŲ)�L]C#9�i�C􌣐����I��s�
,k����ᢢ*�T�f�k�i[�'��/q�����{����B	�n9��F�0�H��[�uwg�jl�&KVO�r�خ7��|
�4A5*;�9n�U� ��J�&���z�?FHwf�7�R����Ae�&��~�`���{.*)���N>,R���8����Q��8�qk_��cy����Zo޸����aNme�-�M��&�� )������	Δ�b�
�����L���]�.�y`���T%�����H��:��#�(��o�v���-[���kV�X^l��Ѥ_Q��	�ߏ$��ED�t�G5ҁ�*l{����%r�AD8%�J���w-{X���<1y�W�G��+�����Q =kC��s��2� B���x��z�is|�6Z͈������Š�����\Gex�v��!J�3^����s�ES����x���a9a~�Y�o�K�R��!�H���F����K�Ғ+��4/��A<�D�CxQ�f���C��2�t�!Y{�s���_}��8�8��f���R�J���'' lف�o�]I�S�0z_�f@0 Ӿ?隘�ފּ��h����m�q���R���@>dC�����x�=.AIQ���S{Q6o�?~���LHU��-n�]a\���{pVv��3������㊑����k���W5h�c�p2u�\DT��U����D�k������=�,.��)���� ��r�P@̸���Og�_�yΓ&�L.BWa�ImnHF�_���Ԇ�0�gU�(,?$}ᅝ�B�q�a�MK�`86^1�����w���gʸ�n8��.I��d�8P�B���^6_T�Ǒfl7������ތ�~���ޠ�9��el���qW!P�Ř��,؟evX��}h�@���NuX��݅/Q>J��,��~��5ς���ʵZ�Z�_.B���#���R��w���cAxbT�����!�A�S���iZ�<q��x1������i)��q|����'�P߅��I���(���Ɓ��3)��&���MS�JЧ#�f��Z
���qR#�����k���_q��+�j1��ZF�+�acz[yV�����yqd���=�s���'=�,������礩�&�m��b�E5"*�L���¦I%&8Y�`Ņ*f��ǜ�R�r��e�#"�g�D�X� �B�.SZ2�(�z���H�n3^a�^L��Y�-]L�[��r���x�d
�t�Da(��$�<��@�%h�}�s����F3���Lz��t�V��\��v��/��4K�r;3�M��s�<H�)vv\qt�����g��͘���8���sR}M������vєE�Ld^[��i_�u�Ζ�fޚ L2�ͼ�ڰ �e���qA��h�鈰B'8��ݎZkS�{�o@���;�o$Ǖ�:a��^�N�y>m`^&dN|@S�J�a��)�x�G�Nǒ:�c`����l@ا���X��5_g�x�轫��f�B�u��cZ���.�C���}(�\F!J󥙎b`�z�mN����ZN�*�&r=}�oS�;��q��X�g�Z�r:���N�X>�T�w��3
� ���%�^�='�|�����e���҅�[.�8�D:-V�$�{������!��t��>ge�&T�����{�!�@HT�O���w�����{!�A��NN����ݧ����qA5�Z����7[ꮢ�B����Gc}��
V�-B-z�����Q~6:ދj�A�`Z����Y�p׽��/f��׷��F황`fxՌB�-�M�`�_�P��E�4���ps�z2����1���A�R
z�U!ES������~�e6�\(�_��f����jN|`ZI1�,Ww��Y1�	���L����	����{��n-@:^.T�f���#���Ns���FG��dO$��fզ>�$�Nq`��d��+kGΠcX|����R����Ke���$<��V����3N�";⡷W8_3X� u�.������;C�3E5�>Nl������,X=)�o��]�؀�L��x�����:4����;FU
�_7|�_c��?��!�^�82z��W5iɫ�:�����3�/��,���ZB8��΋9�fc"�<��n��f���އL�Zf
1�~�U�]�εtj�H9�V�:������;�x�R�|�P�H �����g�Iv����(���ڰ���R`�P�A҈�+oi�#����1���'|��gA��t8Z%8����K��06�����DNl?ʹK�ٚf���֠��Wm��� �����vjF��b29���z3 �E;�>_�9��#�ct�>)+�h-�&��\Ͱ���ݞwɞ���84��i9��~� �<��-S����ꖶ3C�d��UD�	"
�4�U��u��i4a��MQ ���d����<������|�`v��L$n���f�P��71ʊJG�v4�c���\�xb3yB>���F��� W���ɁC�IFz��B��Y�6��ˏ¾�:~�A��J�}(�
��c����A��Su%�;�*��{�?��5Q��-�)�$�֏������uݣ�����2��>���g�0�[?��a-�:>Kn9�Q��I�^�6Z_Zx�6��Kb������V�tα��>�K-�T��OM��}�A���؏��X��D
Wx&c��l�B�����l��D<��ش!��gzQ�R/f���e�{H�(�W�%N%�-.� G��12�	�#����/
�ü�y*��>}���X�H/�J�lD}�]��g`T/x$|�O�k$���ɻהq{�k��7p��*
j�@�%!���]��}����Vh�i����{|c�c�.o�k�jn�{�ɐUXi|�{e��f�̍I�V1�v2���i)
=49αZQ��D)2:x�TĦ���j��X.��C���"9[�x�ʰe�$3����R�ƶt�/5��<����m�ŀ�#�v+V����']$�r �$u�2[T/&�y&��$I��١:��, \�ג�|s���~s�i����-S��Ć\����Z��?d1�r��F{��>N��L�"*��i�qF[zzߍ7�hsڏ����\�����˜�%/�-��Rg�8sTؙ̳pkN��������H��d����m
���VU5@x�1��A�G�B�=A����QO�N�3_";���<`�zj���n}�[8�Ū�P���\XǓq5��R�H���g�W`Lgq�ζt׹RِX��.�xa����)���^c�|�65v\��Z��6�uY�Ҹ���q��G�߽6:�(��{?�3�б��K8�n�l̄��yO��EA�Z%F���'d����K� �g�ͼz�g��FiI�i8m���C`�[���%-O�3e��r�=0QZ8�7Ίtx�XlDkq �����z���N��Nk,��ٛ�=_�=f��5��#Q���o�XZ/���E�Ջ��W�toʦb��yCG�]S������:�z���xKx���֥&��N"#Zo���0Jd.�)θ��b�\&���U������A�(YP����)g�����6�q��xP�:~�O2��C��8ن_q���H�o<�l�g/Q�%`y����>�qݯ~�&��̺����
��4IF��b�9*���U�kL�1���7(��C;��������H�S��0Y��g" òd��L�I��mk��!A�dgF��i��Z�(���*�7�M񖟃�����2:���5��KL��Ȃ}�N;P��ԓ�t�ؽ�,��bH���F��'=l��oj{�& HL4�V����������r�+����Qp���!��Ɠ�]�~l[��遨r��/��$��\K�c�Fc�{��JW`a.�==������F�p��;�R��������>:m�ua�n0}:*m�e�Ǥm,
��@x�a��B5Z�w��2h7%P
�DL����j%���(� ��+�Y���>ڹ�j
N=�R�������JN2�^��YN>&|�T���t>t}9~���	~��6�	b�H�L�y��e�Q�!��]ko�ⷵ�Y�N�H�j΢J�f6��y�&����D�qM��y��ӘУ�r�D�cH�;��&�}��Ӈy��)���3eϝ���*���,�!��[���?C�ɶ?���T匷�m�@`
9Щy���;��ÓfqՈ���yz*�92�П�v��$.�����<������z�_}���c�)��B:�Ҩo\��/5���-q��%������i<̅5��bq�qC
����ޭ/���A,�����mfJ����gt	F�GGèW��~�%��L�?A����ך��)g%葇��v9`F� �!L0j||%�S����9k�	U�cF\��$�w�玐0U�	�8v��t�k��F���DF�NWŮ�~Z"�v�rA<�Q�kȔq[�AJ�b��-�Հ�\�{S�[� G��=�@�2'�h��,���.6�L��1j:�;�Z�Y�d�F�l�L{mњ�]�T'3P�}�U�`�
�)� /&�B�J�K=�Nm�3��ƪ����c�GQb����JMh0y?�T�37�J�7������Q�]��tJs�Ɛ�Qp/�e��ƒE3��Lx���?��4�/�������/�Ú�St�����j�j���v��� ���"ҿZ7���^=�d�*B�%�}Rk6�?E�$����e�a���/ٱ����z��q�3�w��j�V�hl`�>�C,VH#�Ab9�>-CN����A	9���\��K-�L�� �S�vT3͉��p�؀�-K"�?�7����g@cOJ�~ E���1��<�=�,�v����r��[l���3�z�����2���ϰ�<����:+'�?�eFro?���ٰ��?���`�ҰW��i_\�șC�C���D��c���z�ɜ��~*j�gc��jn�<-����Smd�k��f�W�d���m�����U{I��G%���=p�t�lk��x++ ��&�m�e�� |m�q���r=c�B��h�t���E�"��ze�����׊�����m������xGS���H=�(%� �
��(�º��r���'��#L��6��Sٮ�b�$���<I��>N��П���d�M���o�jHT�6�k��f>�jVL{��W�A�납���H�0��D$#C
xѡ�����Ñ�x��'C�.�^?�bp�ȀȄW����5:�
2��HT+�bq`YZ^�d�7�M�����M���>��|�y��6#&�%.�ǉ���=شlF�yb?T]�s'��Bt��%w�	+�`yJ����APt2�;ǖ���n�M�){�R*�R��ņ$���N���Hψ0�m�4/s's*ҙ��]t�J�FE(�E��x�خ-f�U��m�!=��-f��(^uX�6��K�e��P%����Bo�8w:�5b�H��]��څwg��2���q\(�ܮ�kףH�S�	��CeQ���ި!ࡣݝ���	(��@v�(a�Z���؈6���Ƀ��n���S�����w'}.� ��S��ɿw�lb	GP�����b?�e��o=�j!0{���5�'�b2Q��fg��Ԕ��LL�>FDJ(<��cA���Q�F�m���P�Z46ӳ���x��t�{Z.ɧX���o�����۷����mh%ӟ}W��Ug�2����*�.�nAF���L"��~=.R׸��c�ڮ��.Iаr���� 7��Lh��H6���[ɖ$<��y�/q�	ã�$�?�~��4��Q�Ӵ��bM��t?XŃuנ&��
,Y��R�a�2���a~�"�h�F�8�"�î{:�|G��m�Z�D�boQZ�G��D/Zz��8RY+w�m���Jwΰ���;�"�p�[7��)�s�z�
|�t6'R:/�qx=m�N�S��0
*�4 u�s��]3�ogې�>x�����x���$I(K��n�h$	R�?Q(����ma�6�,I�D��̒�S��:��Z7�ܞ=� d5��% S۽�}�4�W0�PR����7�U�����h޾�YL�Lj`�����I��1�q��&q�΃6�ț�P2�2+�R�кr`;��Ri23K8��H�C�T���O�3#�
�����{�%��.�ho!D��t-VŞR.��뉮�� �s�O��DnpW�����s���, 8aҨ͢�0W�8^k���*KSX��l���ʇL��Φ۳V FR3���M/��tB���>|%B��_�'NP���]�D#�Ǟb\fťZ�<.P=r�W�ꗨQK�y�!����P֤s������c:vȏ�'�& �Cq��GF���G�(/G=���أ���O7`N{U@�c���
ΧO��tc�R[�x��>��0t�a�mcX|9�D�2�S�+vBd �Oi��C���uu��-���T�r�3�'�����l1��˼Dg��[T��"�ZK����I6� �_��+mqӽۢWoY����*�x{�Y����煐�'�}7�G�T8�@�Eq����h ���1��yŦ���H�%B��z�>���ʲ��_���t9�s3'�B��Em�j�*�$]��T��オ�����o��S��^�R>���<�I� �f<k���LK��qN��9��*����?oA��$6���l�dx���^� ��a�K]���\樜�6�re���DF]'d���YX*�id�5Wǯ�`�p��x�E�XG�Ԩ7��o� Zŝ�A�6N
Q��k�*ߧ�Bzʤ)!H��{�����|��0(�}���%���n.��  N�a�x����}�i� �_�p^��D7���#�6�jDLd��� ^�``��dsq�g�CY����h)1�����g���B"�s ���"�؄f�Š���Ѱ��G�(+�U<��<]-�]J�Va�3����ߝ�2��=�!�F��=���8!8�*W����\V��ym%�V��~Xh ܑ;��H��۱=��՝Ɗ�GBb����zb�{��gP����)�e;��&�Q��������lM�i�x�.Ǖzɐ�{�,Fr�d`��v������4>ec}+He����^�],;�ϰ�#�o�2�xQ��|�#����ù�v0ǂ���_|6��`�d
Ά7`܋�
�@ғ.G�4���S�����q,� jh�`�Ŝxu���t,
t��n��J]zЗ���dؙ�����,u��Ce��Q����Ü'+D����X�#o�0�?��jϱ6� �=�Ѻ5�l�6K�=>�฀Lt���U�F���I�DЊ�����~�b�x�ظ��q�Vw1|�R%wȳ��!��Ǆ��L�*!c�W譈��\cR�'ykn�v$��<��E�.0�%��$C�����c�.��
hYA�Y���Jo(���~��
̠���e7��[�5�'3S48p�l�a�UvUD���;gdI�������?��V������6F��/�b��{/�<��'(S��W'K�D��s�-��tF�}*�W�:_XO$]�X�H��	�.1��Z�m2�dWG#a����ܝ�c���a��n���0!�VY�M}ab��&�	�úutى�e�K7�0���(��D�,�_��t� Q��� QN��U~=ׯO-x����X����L�i�Z��6�����	b�]�oߞ�ɣ�3Խ-XV�
r���\�LI�0�E�٤��i�ʾ��g7D��e"'u E����f�[ ��
���R#�H=�=�ٳM�Չ��R�EUQT�F�&C����7�{�;�j��[ĵ^Rc�������)�,
�_��+����L��?N�a
/5�x!w�ښQU�����^��>a��\',R5"�����䮚X��rQ�@�و�S�SR�ewe�S��4\c��1f`�g�(q�c�]����k�;����w�!�����	�DYQ��.һ�^��5�.Wܦ�ab+3��
�NxިC�����8�Xt���k�S�[_��vĉ�O��#��t�l�!CU����R��f�l�i��¦E���>�"Zײ�?g��.2�+W�#�8q���_ؠ#-���z>�����>�F��m�o=o�}]�j�� ��>�t���	`������	��Е�g�#��*��4@��͠(�Ç	g ����0�^0���v7���\bu&�D�*Y)�飨o��mm`��ѩa�AARJ9&��6��[��[���.�JB����쇗�B���a*����~؟ͷ�g|�<����4��C퇘Q���x��?���UR����v�r|�"��+�t�5�9Z�|�5�k�^G����֛�D��-�2��4�m�G���5�("���bzL�M���4������#�������<88���ʦ���d�����`��ȁ<ʙm$�b���l�	[~⎌d��7z!���S�cg�w��V�ou���"����}��p�y+y��g�g�Aq�k�ŕ*� �k��=�Qa�:n�R-���� A4EU�/�t���cC�T1UksaI��na��_�	vu�ڨV��Kst���|\Y�o��8��S�������<���xX�m./E��&�af'eIR�-���y�+7���4�ã�_�����f+OY�V�]s��%A��Sff0�8)�*/3a.�����zg)��^�
j�c�է;��v���Պ�X7;�fY�s����
,��/�����%~�8`p/�S�s��*m���J%b��_`�М�l�$D�
�?Ġx	�*,HVy�;�������}�WNA����v_#~��͒%� L;H/5�f֘�I�]Gs Q:%�k�d�������������'�{k�s�cz���p�6&a�u-�"M%BU�1�Յyܣe���AW���ׅ7��J#�ܘu��s�:w���p���i�5���zE9E@����]ѽ���V"�ᬇ)�8��	��k���������5A��כ�h#I	��xp`����8z��p�S��k���X��`��fO��s�X����\�F�+�f�䑘���i��@�l���#��\0}��GNFf��ZQ)Fs8��h��j�zD�ck�\J��I�<+cP����s�f�3r��,L
˭}N]�vp��Wt��ik/��'�
^	��<��0�k��|x���|^�'��ݓ(O۱*��r��V�+���P@�8�v��v��W��m|!fV� ��r�����=�UU��{������hݗu�/��<k�<�q_"�趑8�S( �Q�\ݤĈ�	�a�E�﬏� N�M^�/E��Uv��|�o�B�q=��<�wq��IA>���K�[���z�.�e�p�<�c���V�:wf9����x�0�ā���c�7_���?��E.*���3N���t*A'���#���61f�� �֥j��6H&i��^_��r�[���+��u�#GLmyNDwδ��,˘���o��6v�&�{��4�w:V��a��J�d.��F�fR��VJ�݄���wg�-3[�h�m��`0�c=~Վ1;y���!���}�0��0F�(�(�Z+�Qd�m!�$���#�'��#}�}{�a[h�e��GYf~B�In�4!N[6y[��QT�#����g�O�	u$|:Eu����5�� f�+��!��� ����2@y�߽L�v�P!b��_"�,q_/0�)���M�>���H>�$��b��3��n��7�<��Q]��R�gq
s��͑%R�%����R��C����k`��,��
��V�8�����9Z�"鲬�y��;셬[ 	���$
���;>�؄9���'+{%�
�3��֡�Q�U����,_��i��u9�KN� @��[�;	ɒ��yLDc��6d��������52r���et}HQ��ܣ^1-�r7�~����r�{�0��&ɝ� ���Y�Z�-X�1��[9#������HR�y����.��l��/���.{���j�ܴ#o<=p0� �q;��r��z2����<@������3>����\��D�lS�tSF�z�D �oD��$�O�����p��y@ߗ���;_�Nhs��]977A�n�㗜��WA(��JlO{9��.ȩg��Be���H�q���^��<$�¨�u�}~�y"7p����sH<$�3e�u�]�k2��V�<������:�+D���_�3�H��(��������hѕ�U0�g2�g�w�$A�0��[�s�y�Jʏo��u(���,(2yO��X�yȟ�������H�z��'1;'i@�$�N�+[�H�*��oK�E�ѹ��h�?�S�3X��{ȦQ���:��q+��/eJɬ.�V �+;؇k{���R\����9�(�r>�l1�+ZTI@�$ֳ���؞�Q����nR(��	���� �o^z%�����	�if�S�@��~;��E��%a����0B�X
g��o�C�Xv�a��՗kpo��T��	�����X�]�����9���u��Kj�\S�`�8L������(
�:?);�;�6�q��O�U��vlI�%��F�tT�6�J.�	6I��>o2��d��%	�����q�demH���I߶�Ÿ�3#�xB�����8Iv*� ���;�a|�喜)g�b爇g]�@Dt�{r�x���,�IC�\�C�Ytn�S��l���9�Z�0if�2���O�5�J9�A��I)�N��0sd���{I/���u��C�󼺤ۺ)Xe$��&e6�!Cm��	��]o7�~	�N�b����~���B�D
T��Z��������)N��8��A�Aե��H2�O�8�kDn��)���̵�#(%�m[�;:XD�ٵk��X���&{2k��B�@�!�$���M/�ʸ0�F�#�衁H��ț-���?�6.+๮�XoaM`Ջ�<f�Y2��f�pȲ+�7�0Y ��x�L�.�[sa�n'vsر\�\��n�V��]1]I�x�[���Ma$�Ԙ/}�?�1z�5�n�mː~5pbs5�8O�L���Lۏ�ǪUa{I&%Vn�9�C��唙����5�a�*���,�E��Y;P�jB�qq���x"P���4����MWK�B�a��&zR�L�^��yD?�g i�u���N�d��)�:~m\�����̈�
�~���(���v�D�'���58ۊX)ȷҡ�Ov�sx�	BOϛ���C�眡ݚt�JmzjzS��׻�^��g����^m	殞�:M��j�� 9fC�.8��w��K����]S���_v�ȝ��r6�~�U�n��A�j���Z��"r%��'�(A�q�;�x� Tӄ�k�j1��4/�E�A5��������x�\��5"�>B���ڠGK�Gͬ�l��!��n�C�}��X���p��7�I|�O�^t��9���j�w��x�C0��/�����f����x�"�m�-�]���\V�������{/2����� 7tI(�jYN<�#���r�~y{�-6SP���3���a���A+ A?�D�M+\tw�Ģ������;_�8�f�Ib�]�*�c�vS9�G�y	�X�L�f�U�>�������+c�g5�o~ާ�ۚ����j��Y��ߠ�\{+H�"�6��M }qQt=�kH�.�Y3���E4{)�+�)�Y�,��7e��ǗoV_�@3����~d)L�/�'!���C[�?�ӭ�3M�
�}�g�z��ָf�yC�/�O��pM�K�saS>B$q��e%��FUَ����pl{�ُj�*孭�~����T�6��$�z
?;�4��"�wB2�=��2�n�d+��u�~J|���H[�et5�9����M֭~��ɑ�P����2�R~�Y�,/��[� 4*X�7��&N��40}̒�.��t9��/�m����gkl�+�GG���8ˇ?U�\�v
���N`��ۏ��"��a���S}�[�7iP;�	�rc�T�t3D�����:5}bJ/T�9IR=��c��	��P<���J9�pJ:�v��TCG��/*�|�UJ��ʸ>
6�bM$�)a|������'��a�cX�L��0�txTC�21���8����k��@wg�tV^�'8Ӹ_�jʬ��#����O)��p̚��p��6�&8����\N���j'Q�P�/��
����0qe��~� �ڔ�_��O��-q9ӮϠ���,�l�ݵG�X�c~Z����o]�2~�7��Q彌�	y�a����pݐQ�;����1S��6*o��� "�n�ɆO�\X�����-������߆!:�b�W�z��߅I�蘙���aב�΁�����VJ�����~� fYk,ŃZ�O�!����	���mv`ߥ�(Y�eg��u��L
�Kt�vﵪ�չ�A�Ab=<]���M�,�e���p�H��S��n����x��0�-�i�.,��kܖ���n'�l�|M�h�l3(7 �<���
E"�'�L���/��-�*��XW�C�g������~j�\T
ѥ�k�'�(�@�	&VDKQ�<��;*�U6vè��+�_�P�݃�b�@#�@kL�O���/�1�:�!�Y°��@�'x����4���*�������e��Bb�Ҥ�/��W�n9u�'%�������k�O�d�����eZ������Y�o',�� �%�٢�J.s(����X�}���h�k#���`���M���B��)%����K�tC�l$��n��
]��JLfb�=¾�՗��t�On��ҫj��v;����xߐ� D�318��v�l��9�x-d�ʴ��N|���D��R���D�|n�4B��?�I�?	q���1?<SG>���*�3��S�f�gΧ�*ρ�{r٭rh�"����>Ζ,�}Q_W	�,x����]�1��r�Տ7(Ͼ�0�6aP����aS*�D�v��j([�%Q>���Ɍ}����V�G����p1�o̾��ϞP?�$Gm�X����v�vݴ�]�j�� �L����ڽ!�s�8pQ��1����5��/�[|g����'N�`�*���8X�+����gFS�2AVk�b�p�ظQ|[�Ǆ5HşL#�rԎl7���?o3���.�,�zHo��d��k�� �N
de�QB�c�=��l�܌�D ȓҐ�
��a9��
)�x6����h�+!
F�8O�VS��!*Q0�4vfP8�������:aWهRCK��nPو�Z�8�{H�I�w�7�%�BJ�..����g>� ���~ޫ�!�n�ϡ�\mjK�u\s���(����)�����R��77c�|�6h�f�$��"�%��0�|�x�è�K��,`�L'o�q���נ�m��yQ1i���lH*��D:���f�7�k�Cd������T����$bP�a�%�0+�%�AJ}pј��i�㯪�U�k~\i��e�$����,}J����.P���7����x�C�@(�NEC��� Ƅ�Q�
����ߜN�fw�1�Z^����lZ�e�W9�eh���#`u�o�7ҽ��)��n����V�ʧ1�p0}��6B��2�9��EAc9E�N�������}	H���|>�6�����n����&����&v�h~�s�%[ ��0xb(?��˻�K�N	����|���r��+2C�
;�p1BR�H*�$:��)�� �I�lb��a��Oqr��c��{���ɯow3Rm����|��z0���%(왻Gq'����J//���J7.W@f���d&��o/VC��t��i��"]X(<�:�A��	d��gK��izaqR_�Խ�	1<��qv���9@�lwk��b[n}�갊�޿6��p߳���~���e��o��yG�S��V����o��k����Ɠ|N�T�h�{���� ~��E�rao�����:]��l)������nm��x��N{'��r�h�N6���7�X| o{x�]Mnʌcw�K�)��SQ�W��.n?r;)v������޺�Nf>?"�_��@*4#7B,#lOTJ:ɡ^��Qi�>m Z6�ԥ#�z_��k��<b~������3�(k����	R�j�3���(5�6O�Ԛ��̒4�0��i��}�Ȳ�g���4������i��O��Iȣ=��M�T0��F]���;���n�	)s�a���{ֱp'���������l�t���bY��KT�Uq�Nځ�c<yӤ�G^��$$�J�a��p�۩R���4l�
o�!c�kȐ�T�� �K��pD�P�Q���JWmt��F��3VA�=I/ �(�vl@�Cx<����hT�J�f^�H:���/���R�a_Hq��K}E.�,f�� ��.�������M<�z�2X�vh���p���Ww���8БL�a]����ޗ��T����dߘ��Cm�#��6Y�I�Lo���{�I�/�̰����9�.Q�nU��-��D��.��&�M%���)dm��0�E�7o�Ge�SШj&�-�J�s�^�9��vy}�e�&��<�_�{%�-c��I0Y�r�����}��V󂅘�@����o����ep|�(�.bb��R��߹Q������΁]ˮ���mC�*��cu;חIu�8��J���z�l�+�6�����$��;+���[��ȶ_���:�I3MD�Ny %��W����G�0?s�3`8ޕ�h;Tg��|}e���o�4=��E�wp��^TVg�I���b�� l�1�a17� f��	��q@S�O��<��-N_cT�[��'�3�=|�=���("4��N���iB&	:�ė/|Glf�g ��h�)C���@���R��g`���r��=	�к���Q�%����_ɋn�nWX9�هa>��C"��GC��6��Pa4?��q,9�u�#X
/?�/҅��A�_[e`��CG�J,DC�ۉ�1�Ǥg�d#k��b����z�.�/�b9S��'��"�9���gQ8]���}=SX����͜��Z����v��{��GU"��"�6�Ɲ=��tʋ!D#p� �#m�,@����{�y��~A�e��ሠ� ���}�b�y���#��c�Zl}��]���&���6�',6��������t�S�d�4����w�1߆�A򏐮/_Z+����� t v�V��<�nK�/�S�_�%зu)��t�B8���H5@蕹�W�F�V�)�i���p�>��f ��){6��ݹ�b)��+�i кW�>5?9�'�� �+,�3�$سU`܇��\��O�@p�C9kr1�Zl/
���`�hՎ���x*ĩ�`O��H�����Rp<	1��[�F�k���Jq�a8�X�!��K�P��
w~���jkHҀ�Pm���΀P��ðP�78	0���F�X[��-68� �	w��.JD~�/��%�#3���	J�zm�[��@���R,��YΞO�素m����8�{��ОI����In4#n�ߴ��5���9�)5���%5��MS�!Bb��I�
+��Z=10ʦ�=���WTe��ߺns�F��Z\q}n耪�A:<�!S��/!�-��]Բ����$�t�G}�̾�U;ϩqg;��N�K�5�4V0���_�P�׳�U'a�C�0��e�� �W'"�#������[ްu"�uG�)l���/����_y&4�T�����dk���C9�/i����R*���찝b]�ze���˖�����^�v��#6>�� ��|Yn`����	Vy�U�{�O���"��/5�7_�Y+ ��P�D۸j#55��v䈑|��8�\�b��+�)@��И�#�����k����&2!�
�񛉦�6،��z'$��񓈐�hևTM���`)t�.f�;tH�G�5���VD�b�3%xi�f��D�%�2�����}r{C�ɿ�Eo�hW��g=�A �}M2n;�۹>2	��L�߅�
+�"��*I�fȜ��c�UCޗ��J6#�(a��y<a.��g+��z&_����>(���;xM�� �$lpJ�%]�d�\>�`��h�$��'X�9֎"&�Ԩ#�:=��K+.��3!�WȖ�L�����tC?��LX3�с�� c�ӞW��8X��-��,(��	��_��ԩ�[�N؛ލ���l��"��:9�^�N�b�D:�Alh�l�(wq����� ��;�!��Pp�24>z��Z���|�eŀZ�\��~��3%ǽS:��\jS\�e1V��(�h�q�8[C�ׂG�^@�$^�����\[����W�vl}©Xd���G�s*��dj��R.!��4�ƹl��l���Ε)��;��~�
��p��I3�0R[�> ��&T�$��
�K慶N��ΖW�a1ULB���g1�N�>�o�b�*�A8t�5,�$��@HT�L)�v�"݄�\�"<���
��٩�N�w�`�-�͹����-� ר3v�VM� �@tK_O��#��w�3W����r���WpX���9	��t�aό��ğ�l��;�sq�������l����f�`_�ϧ��q�-� �,��b(�� ���p�k�+�Nm�F��h⠡U�;2�r����f)���3x���OdP��2	%vύҢ���0uJ*����|c:�j(��jr�����!	���t- �#���:�z�c&ƅK�3��K�7�#g5��s����#/e͈JBW`�
� �x�b���X����Җx���R�r_�"bҨ �t�k+F�t�)��_ɧ`
ސzy��f�!���:�ϔ�CX� �`��d%ÀB�Q�ZՏ�-{-��:��鐾���+S𜩌���7�hod.u`;I6)����O�('����24�c��>J�)�w����6��RLs��z�	�����^%~Gu�@e�y]	����b�#�>����j� j�Q�aI&���m��e����Ϟ�Z��:���j���|z�� ����8D�h������Zᨣ&������Ff�O� w��Ͷ����R#k�F��7��9	� ��d��y�~�t)�6�r/\�vBZ���F�v��3�
r����_\0�1͈"����A\�la'Z��{b���>5�j�K>��'�ŁJ��H���Pt��*X��j�]�)se�q^�w�]si������X̖�r 7���M�D�̍���6)��r_���-d'��ªA�3�R[�9k8~���»]�A�l~}p�)�N�+(s~Ɏ��4��U�����@�!�1����Lc�	�{r�Oup�[̖"o��)~�^���Z�!+���CzK�!�V�q#;�mEA�b���.��(�vrL�$�t�g��Tr&��6n�{n5���J�|�L"��yS�ƄzW���riQ�s�u�Ԡ/=�J�����Mt��X7J��^z	�	�(\J�� �u��g��	�7�aynB1W��I�l��O��Ys_��J���n5�ˈڲT�4�+��!~��N�^�0c��tt{��|�L%�����\�P��QBR��6m�oؔ��Y��P0�{�����V{���Dc%��b,H�Sat�a���U
�r��<��^L�<� �d$��u�i.��I��T����+�y�Ѽ������:aGms��sI]��>�$�C% <���~�? ��??�Ӷ;�y��l1G�aO��u^�-��Y�����!��V����򪚜�y'D<iS�W���Wcݨ��6b�T�d�1�c�X�o�m~���G	���� :�)���,��pz�7���H��-��ek�Ս�����;*٠#�i�����D�
>�l��EMVh��#ë��������:N��u`ۣ���Q&�Tv��r�qҮ�����5�0��i8m8�����g�W��nj�0�2�+v�f����؊�(��;k�B�r2���nc���V'�Oi�g>�ޤ%O)n�4g�B�����Uv��%�i�t�	%�+=xF��:��OKlL� ذG!t�b�������'�pv�������߹ӭ�$��4c�Ę�a� ��4��f��;fO=>��3 �J+�ꇤ��(���">�2�����Nz�|ْS<qw��Ԕ����Y���f)�V��H��(���h�{_IW��*�;<R��f�^�g�z�հf@
��6�8�T���lfK��C9}���)KV���T�wj,�
;��@�iJ�߮�E���y���ê�_�g�#t8��}z�'ͦo)��8���<��XRX�e~�Eǔ�#�t߯��4Hf/$6Q�y���%���U�P�Y.㳄��zm��b��.�=�*���	=��l���)8]��|��M��A9b-PSbcg@ ��$�f�_YB�&�?L�~}3jr��/K����=<N����~w'��.���S`�u�	D�קѤ�����`ܤ�5�0j�:M���w��Lc7��{D�O|�*�d���e��#6~�ӎd���	�7k����OpW��{X���QM a`@����
>�_~ͩ|��C���v9�/1�a�F�x����<��MsX�UH!���޺x%��s�ة���~:�h8�%<E���ܢ�����hE�=ɴ3&T	B���Ȩ8�P-v�M�^l.f��v�$E�W�ab(x���g�e��G�f��*�YKӁ����Ss��{ve���Br_X�#n8���t@�^��ھlP.�u��悔.(���XՕ}�}M�\/�� �>��ˉ��쀌��quj�
�ĥ-�ࢂq~�5���n���/�~>�xY�f ����d�$� �.xr��e��G���4-��'�h
W��0�v&x���L���2�pgjp�Э�<Y�L�02!�PB4�R�E�=�78ǂF�}��_���L�*Y����
\Y8H�wP7�*E��04��,MmL#�+e�y	d�z�A��BI
"#n�)��/P�Kk}S���9@�BZ$x���\�hD�tQ��<zރ�SX�If��Y������P
��Ng�S]� �c����5R��H7="���1��Eg�ʧ�'�%�/!r)p�����?+��!���,� ,N�>���{��[�50Ϲ ����{$�x�e�f ��9qR(\�~��� �d;�	�~��QT��O�X|�	�rM�z��Ģ/�T��RR�!N :��}�c�M,Kq����M�
�3�!�QB6�	WC���v�8���L?q��,k�pπ���Yx9n�}�P��P��8=�N��I��c�&N���mӼ��ZT3&��i�&|�&����{�#�u�O�o� ?�"i���"�f]��m�1���4�K6�}��3(���v<�7�d<F��G�ٙ�w[!bcbǁ��!�X����s$�C�ϔިi�۬3ϜC�P�/o%�lR8�֩}6TA�C2��K�Z�ߪ��97�38�ò�L����+���Q¤�2w!�l�-)�s���V�HO%���~XLT[�3B$��t�UK���	3%��*Fɺ�#1��l5{S��RG�c��G�`C{���vic��r��4��))·Zykf�B�Wa���>��t�Q�B�Q2�Q�cWʻ4Hy`bTy��g�D'N��Xr>�*ډ��i�F���c��|�B������p�~�OR?���e=�������TM���#Z��B�	?��ڹ���>V���y�mlߏ�L-4�J�w)����A�B5��Ůŕm��֛�n�����M[`�%N/���	���A_F���ϖ�M0d��-L�:8�|bq���!��x��Q��+2cQ��d�N��rs�Ӛ�wX��r�8���_��j�!��U~O��U���f�ɉoo�u�Ва��@��Q���!xW��e2��ѹ������
�{X�,����)���4g��`�=~��r(�-L
�h;7���n�%�D|i9�Mo�2u�	R��Ry}CLRc�q�\�<2�/��2Ø	����O�:��M,�s�=�w5�SCP��1.�XƳs8�DQX�77?�޼%�d{����	�~~�,G��m*b}$�����K��G���i�Z��gZ]!�nվL�w_:��_U(]J'����%Lxɡe��q��9_�Ǝƣ�!�Pbs�i�RH�JMG����Y��-C���@����m�sd`����9t5rAR}r�Eg�I:�C�h�TA�'�����V�t~'�5� W�O&�v^ZgY�27O�^~���K��=*�'�̓�������f�p��v��Z�J�퍊�0���«�n�B�iT;��x3��s"�1�H0g ��P�;�9[��a܆1k	��#�GPѨcU�9����kݶq�v}̛�A����G�$�WQ|@��JYw�t�_�B���.�:��Yc�O�4%��F=��&�����}��?kϖ-�?M�;1؉汁N�"�x�W l%Zut|���[q>&*�B�q���_-�e�u����ȷ
���/��m�n�I�ʃK��Ѩ�,sS�_��Jg�JK������x�>� ��U�o���%*�iv1�%`J�]�������9;>�.�]�~�2�ٽl|����G���P����m�E������G����\�ɰ�c"1�Gq�z4|ʖƣ\��eYM�M�[�՞."��䆧�9v�g�0@��;o�[�I5�ԏo̪�����=��.����p��Q��!We�x��U����g��il.�!�?�5[d�{�;�%{@�̓��.78;
�ϛk�č�~r�,�v�y_���sG÷
��6k7Ń��Z&Vwވ%�$����[�z�|�dʚ�ۗ���:q��dE�]��v�u��!�^��ٷ㞒���WB�<$@K�������B�ӆQ�_�(K!M��*;�#�;�X��F�(���L���א���D���4�UToল�Ok��HL�q0��%�y�1Âi�M�0mQ1ɸ�!�yq��k7D��'�>�?���J���O{��aݙ�i�-cI�� (~:˙'�Qr\�yB���f��Q�<vWL�/GXI�,�l����S��+U�f�ߣ]H2o�fM�3�M���Q�c���{���p��!�LK.���h懟�B��O����	��Ks���?x��'�*��q�������h=�ݏWU&�Ǟ���:�y�	A{eY��o��ޡ�= �`ֿ�ӝ1g_�#�C�ܞ8V[���Źd_Ѯ��i�����GKZv�]]'�OD})p�t����{�A!(�Q��3���A�v�ߎ�.x�ۭ����͈D]�v���R�%��"�MR�se�j�$�2M�v(K�p
!US߱we��Ư4~ٛ ,Y����	���?~�g�n�%�M��*2�Q�jJT�>��pf�s܄J�#���n�����zm.�]>�K�Z��Ҫ�4b<r%������d`]ڣ����"��OG�9I��Fױ ��|P��D��59�{��L�Ɍ�+�W����(�v4��� U$;O��7��ƙ>*��eQt;�Ё~�&��	��{�S��2q���RJ]
E��K�8e}��i�f���I��^�Θ<���b����W�0�02΀p��M/nEyQ�˃<"���9�էG&�9�Ԅ0L�,��?�Vb����EAAבW��h�����E�d7�	4?��	�S����Kr��+��D8.���w+�f�����=}eL���(�",{I�@DG�6濐�I
�Q�X�J�8}���R�XWB�g��rsK���t��Qp6����wt9��H�������^����"6��ae�e��No��KL�0���-~�`�<Y( ��f[���7C4�sr���@(Ϊ�{f��/�2�i���S��*�m�\H��+�rA����_9PK�i��]��G�|?}�~8�a�B��{:��� �'�ScM��J�K<^�7����=9���aY�>��q9)\��Be�ĻR��9[�EZ���Jݎnʷb�9�2��$�Mˢ��AtlÛ�  ��=(%� R �M����Z(X0�\�OG�nŬs��h��~��Y�Q",',��*�YQ���8��AQ��Y0 �=͋��*ð�K�]�קИ�`��E�)�`�>�W��� �o��	F#��y��=��V��~�����F�-iGLi9�C
e��7ӊ1�@��ֵ�0�������4�Zm�.�z����bS)	�'/z5d�n"�MS?+��6�*�)(�=c�;���n�����uX��H��=��c�J��`q����d���{�~���WyQԋ���-���.�6�4G� d[���ʱ�;3��,�+�J9�$�*m4QZ�������~�G���T�"����K�B�7 �62��K��	]*)Y���
HHC�c
���K[��X�uxB�t|F��7�����L�7� �^�8�`����R}��,��@�_�����6��]�RC���m�B�rl����S�_�qr�2�\QĦ��S󪥗��x�1&W��p�Cb�0�t�����-���)���M�=Ï>]����H�#�+�8�X=p$�-�[@����ȥ
+M���=pqߤ�:�?�o�����f��,~X:�Ɵ�H���idצ	�;w�hn�"�(��lE�݁[������xa�l5G������X ��������'�M,��MXt��4Oژ����Y��s��_ �?P#�`K� z�'�I��R��{��Ӵд�sr3(J#!3�}M��^�q2��Oe�:���WD�^^�pD�.�L�"��W;��|�xM%/�N3� {��]�v��.�	?�Em�okJª[^����������:+��5F�êq)��6��,$/�x���n��C��%4���υm�nD_�`=�.R��O����-�H��,�Ȃ��G~�c��Z��d��� ���ڿc�K���l�p�撽7e�¨�N�s��&���VOlc05�v�**��G;�4�u\��y栗����1�tB�a��V�O������Y��/q3�8 � ߆�k1d_�"E�5r�8Ta��N�����G���qAt����N�q�P#Ќۜ�(Bv�k�{ֳX�����\��.�Y_�Y9\4`�E���me:���T0a�������][̇�}�� 	$!��S$�Y�>�����j���_MXi��hj��d��G<OԨqG^GC=��)��]� Ԋ�:�<�Bz��$-VeUg�Hr:���]v�����~��I�h��`g��rTE/Rœlm])�D2��x{7nPar�}��x�Y\��V�1�D7������]�?,�Jcp"��5��S(���}�r�}Q�/�AF{1\��Z��\V�W�Ū�ǫ1�H7��"�������>�yM��zRe���$�)�H��J����80��1օ����?2��0')���?|��\���	!?�\^�N�-N�'�t	�f*��>��&,�,TG��YP�j�b&��+N
��G
���@J��ʃ�uE��oh-���zq<{��2W�׻�l����L���>�~e�n�G�K�ʙ���9O��g�#��Π�4��;d�E�/в,������0��\N�$�dKG�KZu��b����]/�i���יo�m��_7w*����}�{�@$�RHk����4oU�t~�q�wޮJĻ!U|���ڶ�H9����v��z�LK��b�lsEk�T�UC�����{�@\������f�����g+2$e�+Ym�w��.�Cd�@���g/	4�5r��P���{�:U2qY�G���BFt�MD���?0V�j����EYf!љ�����p�K[�5�-aj�
s̺Ӊ��e+��䔻�E�9�:@&�;X�%�D\�:�&�i�q���.�#�j�_��nׂb�mSO�	��_0=��Ay9�w'�����'��1+��K��4{��"%c̘�5�s��r=�e���9L�Wx�!�$�5U_�HZ�ā�e.��e9�]ee]>hD_q�~T? �2�H�+DO��a�~��������:p�) &�E#,ѣt�u��(�Lj�O�z3�u�[@����4��m�R�*[�*��A&���,��P fx{���?g�P��Į����n)�j+6ɓ�2�V�Qo�X���$�Z��-��N���[��cX�gj[��=�0!'(a�`�	�2�L|�!j5�4��Y������������\���3�!vA>L-'S~�8N5�о�|�n�� -��Nh��46����˛�|w.$���P����sL �a=���� �~�u�yu6��:�h�0e��Oz�$s^�U��)��Fufv\y͑�����N{B����޵�BG�Hd�@��H�A�N�w�q�93�M�-5���?��k���cutŌ�vn�а֓�#��$ ڝ��\�	+e��±�"o��
[��5j��]�ȶ@���O�!mG�PٛǵЃ���=��*i��\:y��W�W)Ʌ�G��f�'n���6	6�9(D�`0Ŵ��=�#1K:&�:w=
	T��'1��\�FۼԪ�=�B�a���Ǡ/�5C����Z�l�;����T+J��dP�,��4H%Mc>^���o�� x���ް�6�n2~�Q�����C��D%�Q{��W�=3�tV�qH���4"-;�3�M֋���vz�����9i�-OXD3�_ٗի����=�����E�"/�����&�_˕vӻ�ژ׶JKm���_��D��R�Z@~%�����H#8�\��`�^�n"�t��j>8.�Bҩ�Q������:��E�0c�$���oA)D!{Gz��E�˔��� �H�U��Zf����ZWn�.6�/���=9�Ay<�d��Ƒ#ۃ���v9�T�fK�+���:gj��l/��Z#��h����^�26Zx��(t�؁���� �Du��L���\ ����n�]�.�1����]��ap0����q3�1y�(��U�9���@�j�(C9��g�虏�xME�n��/��o��:�N��(:�K:s7�p��L_LTiͤ��ͮi�vȨ��C��ҢW��]5��o�,�>�����P���"h�)c�*�ᗵ��e}h<~�~H��{i�xg�����A5������v4O�S�DN��l���:?>7� ո�f���u/��lQ�`k�"����#K��N�sq뿘4�6D��A�NI���$�H�~���Z�a;��n��xx�3����?�g�s��?%͟"۬��S���7X?�9�g
���BA1F�>C9^qA�IΫh~�`���`F|�����s;���W�(o3����	��$�0�^�v2�	��؜��i�V��6rsG��|A������g�O�@�U�2V\C�*|=;��m�������y�pa�*C���l�MW1��\I�G5�_����&A�p��W���\��Ю��ɼQl�Fy����\���N��ȱD�B-(k��$p���*pZ*c\�����v��6Y�5*���Fs�%fw�Ir��)t��J ]�T��Jȅ"��	����ƴ��,�.p0I�B)qsL`lJ@�^5����W���>ِ����4�n�������_�%esj��7����ؗ��ف'�Yc/��5#(L��5ŏ�	>�&��(�x�mOZ�o��"(�Ƒ��o"89E;�$A�5�8�r
��}+����:��P-a\C��G���vh�� |zp��X"�]�@?�� #1�9n����F�Fa?�;yJ����Vw��M�;i�*{J���76�b��L��ُXg��s$_�6b�vMo�>��a�t�������r
���{����"~Hשü��f�����\d)X�2�*Z3@ܵ�T	˅��̇R;�����'���2Pn���v/n�,49/o|<.!���/j��-V= ���j���H�Cq^���? �C���`#�-�[P���
K%����"[Fm0�֋#A71�Ԃg�oy��q{ aSJ��-�Wu]���*���0ګ��ۃ��֛�'�O���9���!�1�xy������}Q�Du�~�B{��YG�Y�P�]	�[���zا�x1{��L��]E�oXс 6u��u'�M���6��O)^o�Q$��Ci���2J��0��iD5�QN�]3E��j��a�	7�L� S�C�q\�8:�r&Φ��&qXM��,gͲ���	v�<��Y��s0�w�-kc Y��Ê,͟ᢙ~qҡ���_��:�UB���o�d�y�v=}���<p:�ڸ�A��eܓc��16�R��0�e]woV���L���~�^�ec�ˏ3��r���`���ڍt^-&/���p��b & 9�.~�+j�<e�x �PR�3�|�LY�b��h�B}�z�b���'l�G����m�Z����:�ƹ�ٚ�@A��G�P���L�w�@:`&!���:���n��\�`ʎ,�,gU��m�Q1�GLגjU"l7k`��K�o�bd�GY�40RwZ <$�)���C�h��$���aH��1i3Kޒɯ#^Gk���i����y�K��G�3s>�p�*���;��hY���w(�����߶��zx	��{�HX�YEQi���\��8N|�z.�i����ށo��o�����xp��s�4)�V��U�_��k��!���:��1�ˡ�ep�I�
q����ÖO���[�T~axRN��;[��X�F<;ݑ�6���1�,Jk��|6#Wo)�h�������Ϩ�`��͙�4���?�faV�d��&,pBҏ�#跗��t/x�t�����>�	���)<C�!:��9h���b��Wzi� (w"��#;&���C���_�N��2�N����Aj�\��O��#hRv���k�PSuY�W,�{���?�gb�I��Y2����{�E�L?rV��M��O�kT�R��*Urg�M
K�c�&��_��'�9�%0���t�e�ݪ<	�!k�D���B�� ����}�;p�k�F������1�k��;x���)�����(��4=�"J��ϼ���hH���i�ر�� �u֨QY��Q�A��|݁ţ�mvq������6+ ��������c�G4.�d��|���W�*X�4͘������ݻ@����>�&k�����9�o�[�x�a�|�8t�\-jf��:oЕ��w���AT	7�k�&�R�pg�Z���=o���er�^Kk?%k��8'&�e2�\������t�ܯ�-y��p)�����f��\ȋj4V"����@fm!3��$i��?��%���Մ�(�M��Pu��Wn�^Y��H����<�0����q��F^��\z�W	ӌ;���3�^=AV� �_�.]��g���X��eٓ���:�38�]��أ��{�_s���#4M1^%�����υ8��"��ɷz�s�p?Hx�"��l���yx3H:���;4u���/Ft.�ȚZ]#�騴�I�Π��r��"��v���>�/[������UJ�&V�V1�[I��k���ʆ�M���ۛ���d9_�u��-w8c�T�g~gW
�Q���U.r�9g��z��/X��b�vL��H�u�r���p<~^-�ׁ
���%t�&[H�|$�@�oX��?�&}�C@*���6�)qi���85��GWP|��U�R!(�@�Ы�� �~��KA+q^դ,2�5C�y#��]8�f��u��'4���FY�_~^:/�p�������FR�`��5yч��P�5J{u�����(�+�{g*�y���ؖ.�N먦ki��S���y�����{.������%'HYՈY���x��\-��G���~��<�&�H���%=a�v����G�����b�ĺo�9i5��ZD+U$T���69�i;�I��p�x�O&-m�19���[f#YK<�W�K�
s^d�t��N�������A\���̷��`��z,��Mu� `��9�X�w�4�ZfҔ�x.��2�X�`��#$/p�'��<o��:avc����&o�zė�K�+&�ǡ]�s۴�Z�V��&�@�y�S�Uh��BE�rBm��_�x�9�q�8��w�g~ó����w4����ju��9/	.�����,"r�5���P6d�p\$Tc6�#�.�F��s��g�݀�:Rc5w2���K�� 
��k4��PA|g�Q�h�8��u]�f�6�Q�h�T��1,[\�F�J�9���cU� Q�U�O���Zv���y��y���A�L��k��/�U��g-��ʵ5�N�$	,壮�ϱ��}W�	�p����׏��[R~�E��v����dn��1�I�ƝB��֘�#�`��PJ�b����9ֳh}�̌Q����5�'*���u"喠:U�����i�K�����J�B͹͸��j��~�nTӀM2:���Fw��5�_��Q&~�ީ���E��=2?���g>Ո�!�21CQ�v���/��g��=����C��,J߀V��ۀw�3s?#"�jq=m#���^��-I��;�R첉��!�5"nO��S��!"�M�as��A��x��q�� Ŗ���<m�[��)1����a1�	����"���'W�)[��F	�BF��"�t9� N*�w(�H:����d��(A{�fC���9�Lu��,�u�]��O�Fj{lq',-�׮3��yΊV�XBG[r�m�#%��#�<�X�O��f�)�u�pQ�zz��8jk�� �;/hQ�79��]�TB/�K��f��Qژ�%�ly$ꕾ�w�n���1�ݭ���D�3��	8��6	e"& 0Z��m~z���,!��y�z�(t�>�W�d��z6��ا�B/���9��	I\%0�	�P��1.kw��2Co�q���jZM��Cb��zՂ�� �o1��p�'����r�?v�g����G�@�Y�i���
=�ߟ�x��d�����U�
x����p��z.{��e1������S��⇲<�x^�����\�7����#Kcs�3$P#2<��y�0�X؈s%?d���)�SP��<�7n�ɡ[��2|����Zuz��9E��
�)I�gz���Z�R�<�� �f��9��id�=�d��Ժ��sQ=oa�R���g�rdb}F^�r�F���dW���SS�V�q	��x� �C�M��fe����(��@��a��bk�>\��]��Ϫ%���;B��]�G�h��6Sp	YFi�=���>U���w��yܩZRK��g�<ELyd��6����*�Nd8�l� b;��9�|`�e���|�
v��1�j��-��-D"���*S����Gw�cVV��j{>?����>҃d#��X#������������tfD?��U,�nϔa8U���+U�y�8��$�s�����1��@�L��!���A���|���[�4����T�n�=dqA�n$$C<N�@�<��s=��p~�X��/�l���uo�к~���J��Ѷ	〡4�gͧ��u��
�HZ�]���`&��~��-٥�Q�M^�x�<�#/�DK-��>A\*I�=ޜa���B
�b8���
f�p0�aVg㰼� NS����X4�7�}�8�S_g��k�,K������@�)G]�)�S.6���YxT�;�+�Y3��I�*]��0��G�*�W��Sn7�"�y:��1d��|��-�`?��|�A9Ԡf8]���pZ�D���{=�Ld4o����uX#6O��E��N��S�G^1X�^��J���X0_��u�WfT|��!<�6X�G���v�*y�B2��wk<1,^SM�ϑEA��?G��P��WR�����E+vGTx?����#�؀��_��c�����6~�h�ڀD;�B�.jV�e.��k��������S$�i�j����R�~~#�w{��d�/f2�&�~끊>	-���AK�e��$~�����6��6��}L�Dc����P�Ȟ#0<�yD�j�G5S·��5��������\e��ҦAÙ��aJ�
J��M�_�u%<�
'7���{��2L��0 �y�̌Fx���wY��2�~PxHz��rk� Z��J�F��I�O?�nL�Q��m7j:x��l���o	c��?*��*{��z���m3�n3��K�T�R�Րz;\���p1�G��A�8���q����:.������,4��j���"�q;i�m��:_��h����[
���W4ouC�� Ұ�9�^�h�� ��%ċ���H�����|CwV�590-Voښ��������xn���T�һ�,cXm�{���X�]���Ck�|R�qq����>}@��W�5��\}� ��q���"	�3o���������G���ݥ���mH�b%q�A�}"s��l���rׄqg�� ���|��l�����
�5W�b�%����ԍ�;�Whi(4���}]Y�}J0��)�%��%���m/�-��[�{]%�ܘm�JF����8�O���R"��� �(♾*�%hl��e�<�$����H	�f��ڤ�dP�d���r��a܃�*i퀪���m����w�����|�~�ƈ�&Z�5�ֱ��Co����\n��Q��Փv[��h᫚=�Xi��.Iҡ4�]�����6�W㸖��QA>Ư��˟�f�4WtfI�X-���"�����9Vxy,c�r��ʜ�!��w���2�=9�<}������V�SΫ���hj�K9o��ԕ�d-a��^<����7�"��#3ĤVK	{eH���\p���,|��ʕ��U��f
�Wr��8F�P�4I�C�:1^�f/m���̂�}q<�n��	uY$��Ҫ�
�*���U*D��.m5�$��k��Î_]�'D�x/h�{�n�P�����h�暼D�CK��E��G�LHKm�$��}�quh음�J��`XAU�әfK0|���Be�Y��:CZM�Ū|E)&]�9����Fk��[�4kp��~��̪�?��$�����j�i@�nr��X��:S���*��9�lTe���u�
���P�ze�3��tJfz�P��_wL "��4���Q�@��S&%���g%3����L����4��PU�;���lǄ6�O�o ��{?�x��4ғ|d��Qn���2!*��0δQF�{�uVX۹y����`j~�����{el�g1�dvב�RC�TR���n�%���/5wܻЖ��9|,hҡa�d�Zn�$ɼ��x����:������T� �$�t�n�퉴�����+� ���AG�V�����?������@�H�c��ZDł}q��sW�r����Q[����N%��9����mix�-�����>r�Yʸ�%�:��^j�ת�Y5�{��#EuH�'  ��X<%��Eyb#�D�������7��X�[���K��ʾ���8�uR�N
p�:
��*r�~O/QHZi)De<�ˎ������'�t�Lm�����-M�y��6�K�J�Id��P�e7�U� �~@�e�DK����*t��J�U.���*��P1��[�~m�OD�N�cXi_����`ם0�tl!���Ik��A>=�.WՖ0����9�{g�����PN[Vq��S�#ig�&��/���@)��`�����(��|/�֐bػ�� �S�%f)��b� ��r�W?OC����q�!�9��m��c�'+X~�y,@����L��y�B-YW@�q�1���Dl>j��vR��=I'��0�����%e���1E?U���(�
 f��&�#��[���@8$�k�)m��>8�ъl��He�`j������ɠ-μW��ئ?@J����纉�Z�s@o����g-ӦaNv��B�򈵢����p	f��ɐ��z(�d!u�GK�cH�DQ-t���n�hC�BZ��;�^,W�sQ5��]��H���|H�`�,�g�p����&^��X[\)(�*s9���)�V�64�ΐ����Cr��f��/�����3�v���o�����%�s?z<�s�s>�m�!yQ���	��f�FD�ny�| ��y���n����	�5n;/z2Kv �6���o�J�n��+u�(�BG ��;�O�����Ck��7*a4x�� �D�}c���S�3�3�lwWL4v˥ ����|O�L������Yy�oΊT���z���ڶ_(�8�I����z�((��:�$�:;1�4UG��ӱ�[��al-��
�=��c44���`Be���v&h��\�c����7����	#	�u�F��j���c' �s��1۪<��El^c�Q)ut6���6����)�8 ���<����#���$�&쒓]6��tj�r���r�yOCD�)gn�X�pL�C^����q+�>D"U��^�w���0�pb�!�R��uKmܢ�w����.}�_ȏ�KB��K���g\��~T�1�g�9������瀼
�ӑS�Q����f��7�׫9�����\%�!㳽�g	�Ƌ�b�Z�I:�Y-�^���z��Kr�5�<׆vs'm��j&ɆY<���C`�	#��Khz��\�kj�k�ċ�����T77]�s`�<���F2�%�مa%X�,s�y٪�q8��ڹEN��ӊqFP\&�/�_��i&#�J�,[1��zk~�yq7��O�0�@���X'�H^W
�>��	�y��zhQS��&a��b/����	�om���|���G3"k��_iR�^��ě�ݫ��h�D]��j�>��c_���d]���V�V��{��H��ݍwDr��&i>FW���_�LQ���t,̅綁+��9NF0؃9��� H��p�uW��Q�� �p��$8r���A���H1u@�&�<��U���V���{#I��~J����_Ɨ�E�pⴥ*RZ�Ĥ*�����V��d���ǔSj�2kY��"��p]hN�f����rH&%u�w��� �s��K�V�I�<��}��@F�l�3B�>? �h���I'fmf�^��^
V���b�(շH�mb�a��E����Ā�qV�U��'i��%�/�c��vxX����Sfu.�{�~˄I��tO�fz8�ɡ�����j@T���kWzB^q�����؁�n�k��?�?�,蔇d�[�/0j�>Uh�?;��DU����� R9�m���%`بlx�"�O6�����0I>��5��fUu�"_z�Sf>���YH�*�:T��'��t�X3mxpUL�����v����"_;��3a��#"&C�V�)g�g0�8�f(�z��p�7Y� '�ʕn�(w�<������h8M�J�j�&uO͞s7|�i9Kh��FmD��(�w˳������q|a\����Ku�D ݬk��=a�f�+,��Mzer�Ly��Gv��T�>j��'���-]���>���THMxXt`��dt k�R����"������Z���{����ڡ����
�41?���|<@d�ֆI����f���6����E��D�e��ln<���V�X���v�}�B�~��� �}�'L�x֫�8oI�WS,��3%��s����DV�)�f�����RĚ\�sT��w`j�t�+H�.���*jb���g��M(�iPe�]�ރa�W���֍��˟3oa=�K<��\�?�������	U���>��
�Ǘ���=n|�8#9w�*��N��B�����5g���+c�<dd�g$2�� ���(Y�#}%��xb�����j�
˧3�=�p
��_��&s�ddk��P��(�Q��7k4z7����R�GǏt������6����e���9��d^�`��r� �׉�0������(�	����}�xgҚ�	<8��x��!?�*/BR�o��t_��p�o���͍��*����������Y��w�f'e�[.\=
q��;НA�W9���B�'X��&p)rO� ~�grJ `r�sI�iLٞ@��G�6_��e���X����]c�&�.� ���+��i듑*��ִ}��~eq�8���Ã�:%����}q/�����K�������0p�r�=�ll�_�R6*?)�ɾ��8��r{��z��O�O���4JwZ�#���u:�&��;�B��R�1����<�t��Tz���nemn3����F)b�d��o0�i�l�'�Đk������R�������/�;�`%8=�^ �Yvk��OF�/V(���g�'a��b ږ#�޼A�b\|���Zp
�:��@�Ƌ�b<'�T
��=�K/q���qzx#7x��T�K;(s����	=i9NT�\���T�t��PX�"1�΁x����X��҈���\���c�g�t��D�%|%��U�O���mY=�R���H���Cc��/E�JԷ�8��1���y����k`+�z/�	@�UX�sFM�����Ix�D���s�u׽���8]<�ss�H��z�&U3L������P߲�8<k�h�Ʋ��i��v !8�$��M׽ݻ�L4<a�j�ѵ���w[��$J��cU>�PZ�[~W��[�/N4dvGJI��we���U 	�#<DE1��Z�S���=�e`a`^���pk���*s�q���3���H���')?�J��3R��  �����.��@4��m��ҍZk��,"_�r��"��X*���
i��&�W�JP:�`�zj!�r&E1<H��q���#!�.�s�H2f�B�[��Q�OQ1;�߃���%�gԡ�.��GZtX��I����؝&xf��:%���q��⫁�����/NB���/�8� ��E�OI0܁Ț~�\��`����7a�9I�~�>�{�:Q澭�ܱ�\����s��6����e?�N��	$!�?�5i�d;N2A6�Hpkf��Ia�pݦI7.<2W�<��o�qNC�����G�0����ve�M��,"�I&y8�G~i��+�w��Tb@��@�<�7H���Rsn��U�V35R�{@[�R��}��S�4��;N�"ᰦ���<f����q�,����m�Z��}��͞�Z �Cc�=B�gw�*χ7�1�"��Z�h"��eP�q�����~!��s�5���B��ù�=ՃPݕ:����B�[Rˆ�M��"R�O ��jPmRm4P�mY;��7״�H-�{)�����s|��l�,&4��%�T��Z�T'����F�|]]���m��5��(�-�V�4h)U�kԻ1U�U��d���1�� �@��H��m�ϙl�u"$_~��Y���9�U|�'ne%��;)�<P�tT'L��Y������6��ڙ��W��5�KYX��	�{�;�Y���zp�G�cF�A�t���IS]ӡ�TP��ξ4	y��-5]☸Ήx�漎�G[a��uNX�����/���(�6ō�v�i�2��v�:���x��I��AA��dW�azǥ4$���� A�ւu�5�Y2f-��ͧN��&��5g��{�G�Kco���EI���<�w��=v����ϛ��:�b͍��B���Y�t�a-�{�.œ���.�O��&��������l����&j��l�&r����5���a�u﯒���j���ؘgE
w���lj)����h���v�r��kt� q��Մm�ָ�'���/�Ki��K���]���F��	q@疍�gP��hMO�S=%�C�-e�y��g���P���6`.u�ԥ������P��SG����b�Դ6Gj)������=�TۖCy��Ak�ӫ�a�5�ZQ�o�J6V�==I�@A ��
�?�k��OF%k9�
H,6tK[I��h���ҤI3޴���}+��'�_�-J�'� 3>�כ���ݝ��&�0���q.s��Q�7>���]��cA�	 ��o�,uO�z�"yY*�	���y7:f�~����;ǯ�g۩����Ɨ"5%*�v2�;���W�*�ݹG,�6]�_H[?�9�Ǫ���8a�*��c��x�Ih�}��r�Q�Ґ� 'jZ����#����4�~qw�kPE�d���ҵ�����&��JZ��0֢���DH��:gE(�I��-�����-��Mr����I�$r�'9�l#J�5�����R�"Rep.�c"f��:����� g���AH�f���Ay5��1�`��j5��j�Ƽ�P�z�$ |)�u6:���w�צ�o�U����,�����}���y��+D����w������u��MX�6���33^�d����8=b�F[��.��m���G���rdf�i�EC��v��,�^1�T.}iJ�}�� |<ɵUe��ۊJ�`_�̉#7	'�(y�9{+-�n��X������&�nFc��\�|���&�I�e���j�0pY-�������߽`�U&����� g��l�%*òUn�
� O���ka���+��+BmP�#���R���/���2Pz7U��߸2�~)� n��B�q�d�;Hn1?�>��f��W0��L����r�z��ú�,*eiBy���{�J��� �l��I66�r�����y�<�]���ʽqK���p!�p����s6|�Rc�����2�r�W�3@��,h��W��m�Z J̙
#�_���^����=o�Yf�V�@$$�3ص��5>�(V���@�����0��q*e�"w�k��a���y��5��ob�������{m&.X�Rg2D�`���!�`�o�Ɣ�i�)4�4���Ą�տQ5�쬟Pm����Fo��Yfъ���T6��Mׂ�]<�w�iG�ña	_|�n>^��|�+I�>;�K������Dk�D@��R��0��݁;�y���:�����C��)�{�L��iWy;wV}F�BP���V}Ա��E�A�v��i�sf��4��17��wzʙ�=��!H�H�*1!ğqb���r:c��r{���������d#��j�������{�Vgh筭��M�x��R�t�J ����:��J_�JO<ې%�:��x�%��_�W9#�j2,���+�?,�
�#ۥu�A0v�������Ν�)� ��5�zl⬝�5Mо�>���1����3C�-=!%\�<P�&\AQM�0>_h.)gJ�x�J�>��h��]v$��	�$#�o��.�3�1@��v@�kE-���a��j���`l�}�&���v.%�7+'�H����?���T4\0rm�e�m>�f��ӼOz3I�]��N%�(�R����.6�lx�˺9�nk��y[1;��~r�Ky����&�&:��I�(.���d�~�a�}��X�v����9%�|���<�A	Z�Bm�c?[�&��=�DR���q_�s�3_��x9p?�}:�d@�X���|AѴ��l
T�w1 �2���4 ˺ΌuL7��i����s���@�xZy���l�a�X,G��.�:�8'�x�	EC�0{2X]&$IO���[ض@��K+W�A>���A3Y7?׸)7��i�B v;����E����ї����Qf�,����h���Gl�j��`��H����˔�YǑ�)�ؒ"�\8�C(���y�#��L�2AMn����K�&gN4�3�W@��짛�xJ�%���-L��ۻ�zsm�u_K�y��A�˼z4���o�"�7.�vo��.h`�"ޝ��r+o� �s���Q�GV���VO&��1={( �)?���b����=�K���0��L�_�Ԫ��l�YO��qw��B��
�(b�{۩/ŉ���j�Tăa}�C;��",��	��]&���qOY��H�Y�z�߮��v�(D����t}):��=~Sr,`��9��D��('���.&�j��|��@J_%��Ш�j��h�X��Bb�c���h���R}�c�o =�2����;����(ƙ)�@��8ބ2�e-��
�J�lC5��'�0�_��R!%����İ������t�#�w�]�ۭE\��nKI�I����gq;���R=f����@36J�fv8�z�!�6���m�I���2nqQ�����M��yM���\w*{�k��9']ټf����ż��Z����hA�Q�N�껄|�~�B��R&NP���Տ"W�.���k��=��f�?�jS�Pf�K��������̿��3Y_:�%�������w�f��e�~7�C#������T�5=3����ͼ�Daq�{��/(�l�����UY�չ��[/��c��h����j�ʧ�Uಣ��4;����Z����)� ��[��N��@s�;��Ӡ����]�Wݵ���/�>�~�ϒ-�W@�7��#Gi0|��V���q/�jI��j��5�*	�[y���	L�h��WJ��: �v|�u7W���Rǳ�f�X,�ҭ=�I� y��P]���=_n�ZGT�y�Q��b'��J�?����@��|�J�m�� ����Jy~��A�% 
�s�;�׀�o2�:�`��?H�tS��F���j��*e]C����ܐ �⊓�g7wMD� ����?�o3���^v���n�an�2v�/.���Y�d|���9���sne_�w(��Cd�ͨlC��U�ցy{.���M�,.C�XqD}���b\l��w\���)��G�3$4�X��:��`+�w����T�p�/-�bH'M�$3Uy�:+,IV5�ZR���+���#�'w����~�{� ��|@�NS��3��%��������?�R *_`~�|�4���*��WR��@�/S\����+�b/_��q��l�!a���v$5����2�.1���1<�q��� ~��ք��S��5.@�I�V��m��_i�V���ۮ3�C%Hkp�'YO����d�ۢ2�e������C����\��Hg�z���B�w����*�d'��-�/�B������l}p��0L(��בی��zW�ӸE�-D�I���讪��DZ�7B{nh��j<�|�� ����t1�ٶX�jn^NO�Տ��n�$\;l��(����3���xѓz�w�c�@4e7�)�V�r(	201��kxb鄊��-��mw�y'��A�I{��*��J"�V��G��������FX�����/�̗^(����XR��wQ'��xW�����8J1�[H�
.�u`M�Ej#��f�H(IWb����z$Ei���d]w�J#�d��g#�L�5��Re���Rd6�6s���<o��[O����S)���՞k��$bC&M}j��Ik�#�m��Z��?������B�P��m�)��6U��466rW;�VǬB&=���w���=�#�q}��ʿ�)f����gR\�\j�
c���8����\�e��"`��q�N�F~S	Y����=Rp�޳�nв= ���k}�nJԅ��ÌS������ߌM�����LL�T�N�5�m�M.�>�xll�m��)�{�����
�*h��7XSq�r%��5o<`�}��`Uld����uqC+���B�� �(H��dB*���M,3;+��|'��%V� �$�ş��2���k��!������#�NA�����N!�J3��B7��򹈛����P�w{��J�l�Op��s�G�1n��`�h��S;o�NIFq�����S �dސ�F��8�.�����ݐ�D`��/����M�E0#DJ~a3����S7�F끂��o����g=��B�ȼr>���CWoD��wd�g�W)q��iD\�	\��}k��A"4�©�9�����t�C��*%s���l���OC*n�o��PkJ*%�`^y�l3�t-n��e�(N�\Z��|U���x��E�}^H��?[��#bI����ZY:utm'ʪACSZ����O�èa�d�o��&��F����7��J��ܓ�>Gw�F��2]*L|�w��k���:��Gyg��U�#ә��V����8hq��}���)V]�9��Ury��;[�ޅ��#��)���оF#r�����|oV�Ki��82��	��?ׂL��*�d3��z��%
����k��5�����a�k����`���T���CG��t��y�����oj;�{�+�`r�nڪ(�l�`��X�ٌN��Vd|r^�y��rjV�ҟ��V	�F ǠGh��l;+�}_[����ᑈq���Y�M��2_�*/��t��[3��VU�P�F�";��L�������.ƺ/��n��\�6V]�l�"�ђ|Xl7���
H���}"�{Q�h �1�g��P*�!	A�Hإ��$��H�Fz�P�xW�f��2���?���/���}e��lq����kmE�=�5�WN�h��i��`|�6-�i�Jf�O2�a���-�n3m�����I(�j��W#�%�cF9��U�ӣD{<�0/��{�� Q5@y^��f�8�y7f����8�6����ڭ��9������#����Us�2n�&p���3��KbL��)f@�&�qw�d\E�UǍ�?w,硘m�P���7�$�(�ų̣�.�}
��I;n�`,l!�@?�#�ځ=���3�z}����c��[���3R���k|ʚ�
@���1n����te7��mo=i�h]	��cΎ,bȳ�@���aֿ3$���%�ɔ|iP-Oo�!��Vl)!BA����Q�&4<*�t�5G!B��_--u��z��݉ �O�r\��h�����ؒ�CZ�U�+�q�� pע�J��^�K�r[us�e���K]�m�����@����'�R�KS}�DY � �䄿S:��6>��e�5m��0<�i�؉�	�L��_�5]�g�+H��\
e?���z�`�~�b��#;��h}�IArƘ̎4�ܳ��A�]��^�&/U�R+31=T�Ɋ�Г��Y@��Ҡf�q~D�+s�~� �?��u�KaY���x\�ܐ�?�Ɋť�4�J�z��dv�X��r�^E���c�������ܾ��2x�����W���7��k5�ӝ��I��\���j��X1
Ⱦ�3�hv@zD������/Bm�5%�l��J@=ч��A�m�����R��"t i ˦s��l� X*�zcd`��\��<2Чʥ���Ɨ��oO�S��D��������v2�����d��Q�2.���E~6)R\i�n�Q�����z[:�������T�l��Kh`W +���}�;�r,����S"3��-��G��!��gK���,�Xb���I��7�S��Q�Y�G�;>�t��x�f,��~k��0����oS�+�
�VRR��o@����ՒQF��IWbC�9�)9׽��kb���R�_����.�E�E��̃��w5��~i�Q(;9�?>)-ASf|�fל��g�N���r����y�_��AP	���bIm�Y�^�9�]jN)n��ޞ-ma�eZ[���]�+.��,����Yhl��rљ������b���抷n[��8�Am	Y�c�?��㸷�q8J�t����Ĩ��6��=%���P�܃U�ݙ��3��`d��8J4�Csٯ���]Y�h�(pz(i�_�r7T���6�%t�.'�̓�Yb۝
g�XM��Z��[2^�H�G�S������k���Op;z�#�Ŷ~?�}&�W�A����f]�h��mi���M��y�Z�gi��:*�%ԙ:/��Xz0L��l��o�؏��(�_���/}��*����j�I��Ҽ�su%1G�Ha�T�~�چ
~@�9�-���t���������n��9L�󷠰�(��E��'׼J�	�Q�4��t4�LN�MW�3�V�_ȧ���d4���,EN���emiBı>�5�H"���VV	��T:Ń����
��m������2{��KK;��eB�7%�^-�ƃ[9�F;�a�W�z$^(�Μwf�_0�C��jD5�{�|���W�%����Z��k����C�lK��>���JWBO��Vl����~����G�M��
�dJN�q^=-�S��1A�b�A�lG(F�9���y~{��	'Q���VzK	�'5���C�6�f9����WA�;g��!p-�S^�F6�[�#jk��#)���ea\��X��0�s��m������k�G/c��^�y�4����cͲ��\h����M��mG���nyC�b��J#�l�n��o�T�@�r��#R�T��H��k=@�D���xl3�5�lp�Y��d��5	�Ă��j�A���!����"IM&(�B���\�T��QIo�����Rh�N�X�������V֘����m��C5H���q�:��9X�&eKh+3?����yF�8T}$�9�"�0���WM���/J�J�K�z��ʉ��u|���6��N0 Jj�ɾX��s�q��Su�_������j!^�E���e�o�1��XjI��PE	M�n��A\����E�2N��L
�����(U�V��q����
�w� ��Q2Z��8�����ӥC��i��xw��JC�Cq�+�d�A�p�t4��W)�hiS��|j�F�!�Һ�k�*��ێ���d��2������o�D�b��Jŉ��̲�Nz������+)& /�=��Zi��!י�%�3�'	$�����6��E(���ݳ�+�z�&(}D�I�y$]䞦��z+�gt'^�݀�i��6o9��ҏ^S�,D�)U�c��rR����G�� c%t�m�:��2�5wp�T�{�����(;7M���M�kR� 'fH,Z+[{��c_6�cŰ�Pk4!�Gi�l��S숤��\�%�D�6�83�Y���D6 H��~dm�̓?����~�͎@��ݝ����!�H���NK]A���p 5#�&�L`����q��	��K�����k|�n�z�}	��Sk��.��˻���Ħ#ʮ�C�\	�uI�%SY=�Q���#�� *m�����}�*
7�Y�;�c��\+$A�O�(�F�����Wv���a�_*N�	���UՇn���2\��s+]=���Y=�E�H���kAKr�$����j��l�H![�%���	��k�|��)7��A�j�Z)B`���@c/���~(���.اZ��e���<�H�����0�OZ%D��3UQm��^ֲ�y�s���CRJN�U�,����r{�{��oV�~���3]������p}$�+oX�
G��H�G[�t�Y"��K�k{t��3o�y�E��H������W�Uʢ������tmyN��E5��t�Tַ3�Bu�j��>紬%?&B.����s�G�~�Q?+��(���?��,�T?O���M��	���k�c`���C�x�gu&����U���?��M`�h�C��ӯY��_4d �G�*!���&W�m�2�McH�w���\�9M�7��F�q�em�������]3�ϻn:!_��6e5���]�;�ȓ6��A{��x�����t<]��ꗓx�euTK�Z�s�GU*!���� Q�=����ϻH�����7��kP��`����s,�U ����%1�	����l}�Q�xt�~���6��\�2��Q�u.'�
��E0x_����D�o�)�n�fT�(�׭�J�,ps�D}�1��
C�pǣ�R{w1z��5�Y9헪����s?y�]{��D#�?J}X�?�63z6\���S{�C�Z�bM^F�}���W>�I2������25�C�S��Oo�z���jt�	�����{��\سu�a3�<���G�tA�"��r&�>O|HO�i�����g䏥���K�T�����ʗ�x��iL�6Հ_��P��Y��y;*������E��1��B;պY��G4��'��#�n`\ki�"�*��S���{!��+�F��u���7� ��Y���4��d��W��*6K��q�a��8�NJ���٤2����UE��5�Q�q�,j��+R�ػ���59^6��<a����%�-m�&��`�����)�Bo�{7i����k<�&"�����,�&�cC��ޯK}��"˲|������߆���~눾�j�#����A�s]C.eM���]�1���Oe/������IQ�Ϙ��s���;��9�;M��p�*jM����%����4Bᤕ/����� @Lѫ������/����7�.K�h�,�v�1���y�
�����ߧak��1�YQ�~����S�?b��gjM?ƽ:�u�C]�t�\.�\m�K���M@X�AI��{^F��^�~�����
)?p�	+49�߯�L˛�[8��&��Q� �=M��7JFt9 �������J�YHA��Ҽ{��>����Ÿ�^%<��e:7�|'��_�[�d�5u �3"$�K��-��bG�7q�Z���6��E7]���f�q��qS��;�*c�x��7� ��=�B��|�����Eݧ�
����m٠��lR@��!����#����]ɚ��߷�]�.�]���^�z�b��C��-���8h���@2�v^]�����}��iJ����"�鉜�.�⟩Y�
���Q�j��i�]e�g�י ���7���w`MEK��%��OG��B�@���tl�X�E���Ē�ė�0� ѐ��q��|9/��<o[���ag�d���Ϳf��1��@`�KnW7�7���ی��5bjz�����Z:�� > x����t\/%����1�&v5�^=7��]�@��\�l]�G��it�y�+��LӠR8��pB1��&]���lt�DR����h��ȥK �R� �6�^c|����C�]�����'\�I��<J<�n�0n�pR��;i�QI�eե�|/�@"�z>������)�=c=�	�g5���c ��H{Ҥ�!�:6�|�_EuD�X�uv83�����VQ]x�~6@]
��f�LcQE�i�r�S�K�$?�- *���@E(�����x'��H�a8��k;n4���dQ "}��Ғо!���V1��pb��!��!#�E��ߘ#M�p�eN1�L5E���AI:'��5x"R��I6��-,T��Y�� �1��s"�rr-
mΜ1}BtM][@[�ؖ�9 �FRr�4��bp��ӵ!�?��F��&�˖mY�qm���n<�?\�η�	�|KN%(�&=?h��"�ph���^��(8gCz�7ǲ�[[!�[i���6�(�1�J5��߀j=���*�Y! �H�L�3�|����7����0g�TP�W_v~��+!��ߪ�&���XB���4KU���_��_�hRb|�0ɀ�ԭ�Wx���>���早A�K��lW��z�-,
X��x�n�ᓲ�M��3"�,�Jٿ�.Q
=���9]�e�O=%���ޛ��]\�3���W�/9�' 8�v��7&�4n�n��W< 2���s�Eb��֓%u�D��hNnx�,7C����|�=����$<�E��1Y�59���+��tp��P�ōHlA��&s^.x��Z�X��ap�I�Nn�e�:�V�:Ү(�D,x��]�ďIM�ư�t��E,���Y�nƱ�Гꈦ�(�;D#����h�iu�1�V��U����,���;�_��0NRA��5�����P���@���d�����<��֎�"2�m�6�ue_Ujr@wY8��4�f=�i����M���aTQW�.��1'�^��8�����W�������H�h4����\�lG���>��Va��!�]^|Z�mUe>���8�q�#�&�bլ+��sBY���?m��U�}@�I[��z��˹�3�iI�G���A,�Z7:�ZԩnX�^;g'�1��ޛQL#8@�n���PN��y�N�>"ؠ�� c�٨E)ǒ��&�I�B��c�̛yO{,�-LQ !ey"��z�_�h���٧`6�P�mx'�Ed��V���-�Z2���x��p-��PжJ�c��0�������Z ��F�۲����-Ş�ù��0z�éɭt;
\�&tE�/�]/WLVn�#���<l��Ѡ��g��D8k�3��8D(ɞ��撶�+�?/h���z$�=e�P#������:�44��q-���?�e��9 & A�KU�;������g5�!�{��^y�Ϗ��v��(�L��P�][��t�>��
d� �q\{����w�	g����i��,9njO(#i����|�����A̓�Ng�mC��P�7�1	Pj��'i��U��:R�R}���)|�FF�/���7�Zܛ���  ���X��)�LѾH�4=YWEg�g��D������rZ���c�y��Oa��v�2�ی
�W�ffR�	"���Wm���s�7���D+��\�ӗ �)� 7^��]\�W������.��5j�E������p���n����V��H�`(�D3-���$ ~�Z� �*l:���j����a�z��Dϴݚ��� *tf���`)9l��'������k{��}�L+�ӕ����Y�.I��q�Θ���$�^�Q����[���9!c%U)�>Bm�]p���p�`��k%�\�$#˗p����K&��b�Ǵ�	��_-��lqrqʰ�S8-�\�ǻ�x�*~��Z��^:��/��
�.
M�>�R�
�tA�|�h��ǋ�����+��g�H9���C�5��
i�+��N�ʷ�,zG�\��z�:��x0�V���Շq�RtLr0�v��G�q�-�G������~٧qQ�Wc~�E |!�ĥ
H���x�U\���U�I�� �x�z��R��}$����qj9C�L���I���j[8*�\�9�V�K�p*vY�;S2��K��Qv-sZ��a�XY>tD�u��]�&[,[i��~�^�����I"��ׯ�����vN�^D1lR�҂�X��t�{�;�5s���C����a���6Z�����|vT�,h��pN���g6�R��65c�5=��ۛ#t��1���8{��69��[Jke�B�S�ڌ
��	���9�YO=�e-�p��N�u4�kRŚ"+�H�ߵ����]�շ}���[��͘S!�@�F��gh�:�V��Q8�|0聱N��J�Rލuf f�~��Q�?2gOxV�g�$�]&Lz���~R�`H~91P�$4�14;��ݸ�����	��#�)���m�94�F6����5��hW��M1Tby!fz�-H:�XJ�VD��EE.��v�#� �x[N��t_5a�Ҍ�c4�m�$�Go#��*̏���shHC�iP�vy��9 pF?��4M@�3�<����A_'~g��g:��@��R�у`������X�A6�	!p2�!_�t]�����<z�/�$�����\i�)�*$X��/��օ�d�2O��n"-��R[ȡB��qR��&�����Nx=�G��hc؈���l5R�Y \� �)��p�K=���"iR4�;��zҦr��ՙ�L4��-��:璘���j��P�����FXRӓ�,n�\��lŔhu�L���:Q�~�	'p���uhDW�ܷQr��1�Uy�]��>�G5H�_n�޽�7��!,�Q��(@R�f��Y�!�1�cK��[��5fY*I�ǎ�{�lUK�i��M�����n�&'@?�g� X��L���W��.�D��^[�&�8�C��w���M"�q��;����y�<(����^:qX�AM�K�3�:T+�?����M#1H2���wݬ�{ Z&:B/���4T�<#��y<���W�׸����B�L-UCP��9=A��m�o!8�}FG'�j��+;/�*�)�0����VI�,t��T��&(��t���%g�k��[�ݹ�YO�u;�I2\)�`V�U�YOq�*�x�:_OĆ�X!��15#u������?�yH$�va�w�tN����ā�0��b��#�tIQo�
sqng�2m��@{P�)�a
=�<�)_�9��&����$^���"7�<�A6���wF}Y0��z�E���G������E����&5@4�Ve�"h�|�*��aM��W���
|z������9y
�H9��E���ʋ6��1b	��
ڳ�2t���HD��m�2�b>�rk�`/��8R~�x�(�:�%�?��&� ��g�m���A���<X�Y�"��.���9���C(W+�	���ŀb@c���J��Ll�)�!6^�o��b����T$4�x����eq8ܵٻ�;Ir飯,�1X1��s15e�KŻv���-5HgL���]�x��"����=��B�8��hR�9������B-�3��������m<��2A!�62��<H^��ن�:_1�- ݓ)Ib�n�@�P���+V���4��X�S�TYL�V���pi ��$R��������B<�e0s;���yj9���fe�i�.��|qX#�,��z<\�Y�}�0��.�<��DڋiٰO��s9�� ��H����5�x^D�=K|�e�+��~�\�O�p�LQxQ�ݥ=$����	8��Ã�G�˳�����4�y��m<K �S)|:��#�f���{��0M|^�,��3�(MA=���\ĀT����,�W'RD�f���s2iˬ3
HRN�]N�n'��X�J��yP�m��P	�]��R�)�ʅKm5�Q�K4���2��c��Ʋf޳��x��>P;�+�s1��5Z_ih`�����had�l�]V�BR&��`����@��Q�8#��$���;t�la_S��� K�����}�vgX�Vg��>��YPT���͐����������Ӟ�6��h`���=��m<:�#��ʱL;9�Tt���ڷ�Ώn�#��'}�j�4j�XYݓ�k),w���5�c��E�!sū�B+�70�,�tj7����3�
�9��A~/��E-�/ �\�����Qx�]�4�כ?ogHx�����`�^\�J���|�7�+�E;��\�A o����T:d��3��t��"�,*:U6
�� jMI���<�D��C�B�u���'��7��p2���͕��{���1z2�#���p%�;a8SX�q�1yT�4���Nmr�����~J9��P]c7n�(�"rL�����f����E����G�ß^]�
#nM=�y��]�#8h��5��U��*���<I�-|e.�� ��+q����"I��i��Ns�Z��$߸�(�!'	�� 3H'߈�F��}QJ#Y+1��5�g��h��d}���?�(���}f����
�/fν�]��/��<���2�;�z�x(/őN��Y~b�/�uD�vR��D�5��=B���yc��t�D��[�ζ��`d�x. �km�LC̐+-��C��@h��[
�h9Q��8�	z�ϓ���q�I�<On	K<�����������7#�5f���,�Kʡ�\� �I�-q��W'�׹!��t����թ�]����w�m�.Bf�[��^�HI����ǧ�UKK��kY����ܢ�`2�ó�E&��MM�Jq�@��6�^��gΰ �R^���ؼ����Er����|����vc~�4Vhܝb�b�|���;�KZV�����xf��=�ԡ�������\o �d[k��Q���S��*�f�<rW7�_���Q3�n�P��A�yٟ��`���M�#V�����>���⮧[�2�6�^�IJ�!��7e�	ţR�XmDd��k�����#��|W���d�ī���,y��3��v�pA�� ���W�Bl�&6M��������}5H��M��-��֞�N~Q|a(��N+��VbTGh�{F;'G���/�N�v݋��fb�G�o|C~�4�`��!�@�RӤ�D	E�8���Y�F���}�d�C�8�'�%V�j!(d5O������q�T�����t��>��hx���?�h��2����1�no�.i�+�rxyb:�]QtĞ D@�k�i���3�~��^~��J�ٕ?9��4$��J��Pq�?���W1
�� ��)/��֔J��LJ �WY����&j�V�ff�Y���� Yh/Q���4_�Km����+��?"Ψ��7Ո	��.5�-�/�t3#xA.j ׃X#{���^��5:�ȲM�-h3����1&�$����s��eJ�q��+������$�=Nz�n&)n�_���j�25l���8�����ͣ?팍��P>�o�H �첸
du�!�
`�[&��m,	-�$�d��|�M�>">k������>;�΃O*r)Z�6KL�+-���&UE����ggR�h�'��;���l��� �]��-���	�ƭ�g�:)��g�Ҝ�K��"�J����"�9}z�)�y ]�C��%<�ЅD֝L�4`,�������hg�C�
�Fk���h@�	G��y���~�* �
�:���bN<���7�ȅM������ޠ��Cț����>� yw�@Q�NͶ�	�w\}���ҵ��ץ~�R��l]�tV׷�fco���{2D1�?�TϓL�=	Pk9jSj���U/3mǁ�~�M��V��7.��~��du�UF��F�������:�٘r����k�?0�X�1#Ů��.��m�҂~���q�&��/B��REm�[u1@��	zGR>��,6jeK���E�n�,瀚 ��7Sd��x�C}xG�"�E�$��q�c�qg�BKx,����Ø�]*<�pYo@�OG�/�_Da�O��`Bc� Δ��f��JL0�M����Y8�Wi3��j��!x!��ˉt�t��E�����St��Ѯ�J��Q���ҕ�Z�i���Z~����E��s��'�d�ڜ���bI|��.�>Ggèe������S����3^o�s)�_��	M�v}�L��6w�� ���ks�mV,N��R$����\F�{�t4�\w �B�f�4��Z� _8 aЄjE����}ۿ��Ҵw޷ܾf$���d7s�+c� ��!�ʧQ��0�j�m��A�&"K�I�-�!'6*������DU�j�W������\.p�on���UkD���'�C:��
$�K��[��^�Z(����1p����%�L���k�'�I�I�n�Udr��`Os�	�Q=�0K��Ҭ۩�G&y�YaPtsd��`b��S|Z+�)������A�4�}yߒ��<�K�NG,N��==���
�Z��OU��H�*O%����R�Ch.�V]�����֧�4?�?���TC~��������>�����m�Ԁr�H*'Y���N�͖gB<����Dyi��cZ	��hA�W4� K���g���K�r$O��5a��w�#���U>$sx����^�q7�[h�4��d�����	S!}�R��g�H_c���&1���M����}~��( �d�S`������Bǻo
o�8t��me�����ah�IZ���*��k����ڲ�!5�9����9`R��/�,�����bOي{q=��#�5�ȣh�Z�$b2���֨���'d¿Z�֣jE5�]�l=���;g-��=��J8��gxAuR�(=�Ic4��#�73��~6J�<���	ѭ���]�1q�ү׊2¨Q��6m�鄗Yr�4�2�բn��:���Zt1�TR�%�ߝ4��7~vd�Jx�PUL'������܆��r'��_K-'0���F׺O�aKW�n�ԩe����u؈z��I�`��&̉&0��2�������E������WY,��~V��؈ڣ���M�Ti��*������hv_���t��$���!��E�z�<0oYUTUSӆ� U�)��=�N!U�s�~�Ұ�D��gf�9�w�:��uk(�?i��6yY�LwW�W�?��n*؜�4���0�@�PtH�$�E#qw���r�BcW�)�B��_�ؿ�!Z��tѫ67�����uo=�u�V�"����NR.�3�ML�U�� -�1�2	;���������9��QO,�u�e�k���N�E���	>�J���
����~G�+�,��#| �����e�R�K�"+R�o0�)&^�U�P����~9+�Z^�}�i��>�S*Pr5F��܉m��s��e�:�.�.eT��O��{���V<�кO*w����#�rA�ce���6��R �Qo�\�2*ԃ�9�}	�p�ָi��Y�b�f����CA0O�9��65l�٣S�nB'A"�a+$سUB$�\����*��n1��H��y�K{��t6!W=�׾H{+�ht�0��0��F�Õ�o�,
��#�Wu�����9�_�����*�Bq��%�B�C����[Ӝ	-��$��j�?�r<Y8i,���iuny��C���X��
�J���[m�@�钩�����1���P[�e�i�[�-�	+O��k��6�/�p�F˽z9Hb4"^��0\��4|�]�}GGH'���VxVU��
�k5�N܆dY>]1�X���*1>�I��0�_HT��G߹�m��km����g�X�>5��H�>�G#��Y�Υј�֘/%^L�@AET�L�o�.��Q�	����`����{.	ە�s�33�5�ŋy�>�*eP|��~ˣ�ϖ@Ei����"���J�ۥk����xZY��QEJ :6kG�j��V���h!\:���P��>���������ZJP?r�
��_#*N4���Z[U���]k�xc .5��5Sٺ�)jY��v��h�"��e�;��י^�ق��Pk�T�^����{�,�7�O� gn�%�n��W����"��h�W����򆕣B�1F�^g�V�����
�q_�B��Q�|�w��#B�u���+2��ȂBaվ�lG��w�'I�>m�.e��	�m����?��)ɓP��9/�b�"��Ԧmr�h�L���NZ���}Y��y:�R�>�͕_�f�6"� �F��*��ub4 u���d2�Q*���A<(G��_�4��s���k�T�#|չ��(N�%I�_K��J��:�$q��u1��ܳS�$��UD��/�a��O(~ $�x0����cBu$BW�#Z��PU=E.G�:-�E����T[Q,�����F� ��!��|���$�6:�ݭ���)�MM�	�󞇉
*���E�����<��w��D�4�gӓU!fW"�� 2� ��'�7�J�EQ�I.�c}(�:�]o��r��|��p���X�Ƞ��ɔv�L1ҋ�̗P��^Q[P�[��a�J<Z'�fx�BM���ߐ!�Y`d��p��Z���=�G�=�����{��[%%1��e��-�X��wf��G�t����`i�5!t[��.��~c\V�k/%�"v�X���MuMzp�qQ��1%��h���_q��C�q��7�qA�rX�@8!(�|�/�^������4+�M�3�I0��ؒy�#G��5�5�^I|���ײ�#�9�s7z3C�xFKQ�� �N�	ݼ�Ղ�6��;�@Ƕ�7��5iv.d	��q�ا�6��S�Nt�6D�Т]ݾֵ�z��%6�g.��(���K����{�n!�=p�5��P)�xi܅�/ު���XQ2xEl:&�	�a(¸N=�����j�Hu9}mc����>tX�r���#�P0gIP?�ط����71Ms�M��!:I�K�>�BE�fP�~y�;����fw�rAN�Vp�o���ec����z�~�F��G��)��8�K���F�������Jc���*-V���8i<6�Hg�+.�#˰���3��L�Ak̯$���EMi���K���7im�]1nWbQSQ���Ds�%�.�}�����������r�F�f�'��U��C1��Fu�(yۆ��X��V�ٖ��C�!��Z�W|�cP�mw��y�<B"���`�d��������o�x*��
�Ff��-�a��[�1K>�9a$0������Vax��&���G��� 9������Z�����ƔȨ��@dQ���$�R8�;�C��V�KZ��BL�`L
�u�"���?����{.\k��kj��}�u&���w����=EH����_Í��.aX?~����k���X���c
�
| �/Ct�1�e ��?�E��wZͬ�n:�#�������D�0�̙��i�p`t��Y�z�uMH0؟�P�$��?��
�Ap��B/��R�,2=��旝����
�&L�q��X��Hpx��n:�.&E'!�k�t-� �qZ��>H?�l�h<�oz�b��Ŵ�:���2-���PQxv7��!��K�mzBZ`qt���ǳ���
X�-<~*VUX����p�:���k��<���e;�'́6���|�U�b�3R'r�&�Ҵlo謵����<E�!t��'sv�Oh�>��|��IN�W\��P�	++V��/�*u�����\Lat��O��ɤ%�s��w~LGWtmm��x)�Ab�.	�sEJz�=u�����+=O���>$�:�hNX��*7,��k�>�sc�|�)bD�P��s�b������� �¢ݕ�u[�1��/��SW�|��-��[ә�#���N�u�kѣ@-&�c��:�R�i$�vE�W����6u��p�It�M�]�C�[������ġ�zi�2��"�� 
F"���&Ol��®����*��h�R�F��G/��S�Ѓ*nk��t��#��F�>t.�d6�j8]g�{A◑��dV1����=��~y���7E����fS>���5s1�__���kr6�)]d����'.�hrNǑy
����,��t�����;�W.1��PZI@�K���#�2{�D��Xu��lkT�BMr�(k�Z����XO������ǧrۄY�ɀ�4�a�D<���PC`���סLk�NX�������5���d��ѵ	kxt뒧EO��$�o��Wd�Iy�{
Ő��//������¸1lp</o.��[02��5�;#B��%+k�����%9)��ʐ/�z,#�XS�̥T�%�{����F+qz<�TX�d�K�����ߪӾ��6�G����@*���l~�嵑��&:E�����	�ۼ�!/}`��ṟ.�\��-jp?�Ui��Z�ǻǽ)��fWv��	Z߇����ɨ>���	&Xg�Ж��RZ����� ��CNF.T6�	��$N@��ڠ�VJ�� ~�Q�)V������%g���+�:�x�$��������m���_v��X�J��\(1�@,U�(j]�:�c
�=�&J�������qp��b0Xa��K��r7�Gk�����{�3m�� �x3[�A����1���`�T��JH�|���P�1���Y����QZ).��Yqn�Fs@�������Z��ʗߓ5L���1��r3���2Dz7�d���J7X�����j�t0e���2p3�4`"�	��ge�����׍���qH���i�P���+��a4_ӀGNu�0>�ir��~,/�O��)�Rl��hK���U�@�y��4Ү��w��ޭN�nX��,@���m��]�㕡��4��<�Y�w�=Zdj�)Zܚ��64J#�EئI��>�pU���w�8�����Z��@��^�mY�Cog��p�ߚ���y}�m���dx�ܐUO�����]�RB�sFI���
|\�ܫ�ʼ�3�#T7��w���4�:A�P�S��b?�TӹBUOW7�wH����SZ�*m�W3HyZ"�>�ߥ.8���t	9n�D�GK�q��?%֫]9�r;O�5�����Q�6H�!��]�����]&R$	�F2p�&Pi=n�[�A�$�Xہ�66;摼�n�2//5ਡ����y(xm���
������� E
AN����������p�M/�X��"�.�=/�x�R��n8���Ѥ���V$$U;IfN�S8Jt�>�k���&�1�C�hS����t�
efѭ�>��;3r$����J���$d;}kLX�T3��&B�z�O���4�Mۗ.%�%�-����l������3�F��~�d�����t�uV�$�$!���)Z����\����/Lp�|<-,;`ʐ�z��|�s+�����_]����_�ς�����N�DLa���9�2����
"�p�@�t�V~d@
�B�y�!%D� ���^�ee"}��� U�bLxLʻHxN�oF�����S8������W�z1�����:ZE���~��d�D���8聙�q΀�s=��ܾXu��}�\Uz���yA�v�r��jUZ�J�m�J�ul��4�G�K@�(d\N����� 
}&���r���t�
�0;ۘ\-��G�"�+2�⻸;�c���<m�o�
��/��XR�a�1�3�ÐA�����0��*S�O8]V�TΑ.�WnN�Z=\Q�ͭR��|Vs���{8�S���G��G�WPw+����h��?��҆ƌ���#i�dl����8����`(a�	"��C�!�Wb��ck7�����ڽG�?�4��*}7SІ�*��<�'y�g
��N���C ��3�o��_/q��i�eBΨ.}���}e6��^�c�{Y5�,�4��!�,��	S\��~�㸧g�0)�Q˛�l�Jh#k���o K��AvM�x��w=D��,����������|�@x��>���oQ��w����V��g��@f�$zڟ~g�1��ZxAVP16OM��БUƏ�<�L3��cS�vY�z���{�0�dSt��n{���_`�E�y��Qt����1�P��`_WA���m/u�	��Jz-a������MVr��<o��TFy��:��8`	ł���:���tI�Lo�
�-m$t桲�\�Hk�U�a�HKwR�ڶ�5�t/
ٮ�� �D;��.��#D�wfa�D�!��u�i��HP���ph�����Y+X2c��q�زK�Q��ﴶ�7@�$�X�&i��囔��������]�m�?�v����@A�Dͨq�O�:���O��Jm2F��m��lt�Z��`��>�A�j��R�r��kP0~�E���tˀ��Ӎ��d��k��Vq��,�Fޜ���a��쭩	m3�8�-K�,��6<����r\9�����bw��6�g���y��4�g��u�z��GϘG��ҿ��8蘺C�͊%Sh�tu� D�y�]��4�;%�\
S)���gAͽ:�C��0m*�}k/�%;���:�\P ��k�LQ��z�q��@�����<C�xPos�&2Y��a��}ĒM2L(m;�1��^8�{��橩�nQ�Z�"��{1�2,�Ք<�>}#�|�$����|� v\��O�@�f�V�_
��x I�H�I$���h��q=;��zJ+�z�����.�<uO�-$T�aSF�W���1fƑ��W���ldt�᪼���~$��{�� �yO5A+���ej����a�Ę��*Ҝ�����Ȑ���H�?s��{ﶀ�e�����mS��ϋLBzq��P>��� ޏ4�ǋ�)	���~������|��w&�y�<�v�����f9'J�vs���.\��B�ڊF-9�\�;�W\}�nB�7���_T'fvh˹<wi����es�E]�b�Y��vS�!�b�2k7}u1.�]l�� ^�!5!9�����U½��n3�[����c���X�i��&	���d�o\��,�Q����F��X��D�/�!P��W��n%#/�!�	��'Q�4�TV�)=5�H{��`ɍ�/��jC]@�S���㾹����W~H����]+L��P��"�~}��UR��aE���P���Ј��U�Z�%ñ�sb]�,v�mc�`��U�NP�~�\�6�����j��F7F��g�h5W?�����ߕ#����]�m�fPW��1�dW��Qbs����*�T%a��z2\Z&��qv��.�[F���=d9����E�H2��<�����^V���WaTZ�Y�!)��`f0�`ٖ��V�F��j#ډp�P!� �2n�	kH7�2]Q��C���]�JG�!����O��Nx�Qu)��d�jj��|.�7v5�-���Ӽ'W:2u$}ߺ�Z��SD��n��:v�d�4���~7��Z�4���.������&u�Rf����p�ܮ��ҳ�J���?=�S���������͍��L���>(����&���1@G��)��$\FF�#���O��&_`S��Yq��� }r���1�\�U�r�8�M���\ �L�=��F�%�'�U�>����s/"łB�O��������?�>�����A�c>�,����F��͋��U�x��^ޕ��k�I���xe�p�����J�����:���!�u~h8t�f��ȳW(R�pO_	��K��P�<�`qU~���?��mD�pL+��֬�u�t�?�� 8	O�Y����$yᕉwz�-027��0Ϻ��� ��Aw_y(�T2�����E!�H)�V��7-F�$�s�>�oh`^�=-�M�3Y��Y'��[雯b�5�k��v;�&���]K �����K�B�X�X�i�����W[U�(Z~1����؊��Jhqcn�_N@tn�W����)�4Z�Q��dJF�K]��ԛZ�i��J �@t����_�|�ώ	��6k�6t������p��q'��1rD����QK�9s�]M_�F���W�����ΙCmR�6�ΐ���b�#��O������Py�,+D����l�N�0�� (	`�TJ#����R�s����7C�ŉB���J���Ә.�W�p��n�4� ���WZ�O�~�%&�R��X�zu���K�D�ܱV����̽��}ϼ����\گ�A���x5t\%���iE`LF�U�.�� �Q�l��+| %�pF�'.X�u�$vޚ��NN�rӃp�ʔ�`�E��!dȾ�A%�,�^f!�)ٴ*�<�)�۲@.[�b�׺�l�=B� 52cHY���O��5z�lj�X�P�?X�6�nM�{�蓹�vH��ƺɍ=N� xy�Nc��d��#Z���wT#E8��3s��d��Γ��3��Š��acp�rԆ�e>�V=U��&&�s�7��*\11��áo8��LOHɮ}o��.�~җ	�53�t270wE��j�,��Z�!1ë3���l��|�stO�7�ӡ�=S*��R%>��2e��֏��/*J�-@=���B-��F��*��3����/���y������3xp�<��V
���^@CV.8������Q+����tE��n�ژ_`�
��!���Չ���3�s꙼�o,�V	}�:<��@���P����A�L��>���֑��+--�"�����we���;�oa��e�I����{��	*�D|��O����B�k���[`�$\ǔ�v.=J�f�Jy߆��L�Ȣ�փZ�6M��|a����N0���+K�b��T��)��6�K*h}��#��ZA��b���*�apS�.�>0��2�5�'�,�XD�]G��Ց@�XsLc.=yK��:U00Iն��{�+���<�6�ȕ@`=�nMW��Ҋ8.f��J?+��� �%nF>�Ό�u��*�2��`��\�����z�l%H ^�W�Gs2�#�ޔ�9�A�����,�ͧ��MZ㊈w=�8ñqdOO��h9c+�&����J|��r3�a#ͦ�����5�����'f�f��/��fKU�[*�1��p����k�^�juԙ���/[�ZR�v!�s<O�Oc7rA�H��N/��ٰO,�
\	�O���k�{ܐ�Qu��PdІ��A5p�Ԥ=`HR��p�3�;�<l"���$�DZP
���AA�`��]D�b��L@���h�1'��.��б��lCB6e�P�ʺ	(W��_�ma�b�����g�M ��WG�;�,�Ua�-���Bᐠ���%"&�Z�aj�N/����J�����wY��	�NW�hH[��(��j�Y�qqE8�Uü0��dQ������n#�^Z*���|4��x��
�j�X6�7�U����7�A�����נ�9,��s���o)D��P`�6�5�ܱh)gb��C\R�L���@�N�;ǯ���S�i ��J����G}6�NX��PYM ={և���˫���@�u��S���s�C�px��`�U�����#y��^��'�d9f�z��Vs.$2b���U#Fś���9}t�O
H�p�ǒ�Ѽ����ߵ���O��Ņ��HU�ګ�p��$y)�z<��BH��-2Lf��^٩���Fc�d�1����6�#y*/�C�>u��K��v��k|@������20(��fhQ�j+x�������O�'B���Eg���l��ou��J�A���^�9��uf�>��a�úݜ�2�b�5,h��@�T�'���V.���͕Y���CI�/7�I����L��	~��+����DX^_�#�L9�*M����T�C�PX���F�	�<��R���=/�2�V��`��a�uAV�{N��'���ݍ�9L1�@9U�Dn7�6�����	}�@��,*�;I��?D���qt{�:E6�����a00k�E}Z
��K��r��ܴ2����j���D�˓/�y�g�%[�(k�TwO�F6�d6���3`��jzk�q�h�
>VOw�g�v	����E<u�S=�q +�Ȝ]�N����V^�pNϒ�nb�$Y[DAy��}�j���5��K�q�.���K���/�JW \_sh$��p��e�yگ�<Z���5H8��a2UF�]��;���s��a~�7���T�{�-S���dG3�]��x�
+��0���BpkM��O�� ��謑�;tp����q��6`G<xL�Nb��my�t	��oCsWY�� �'D���ʃ�>��aِ�5_U'��-�Q�%��(�������&S�hHnv�J�m(r+~��f�U����C�Zr�n*�`�׭=��x����n�ꉡV���@��DAD럖2�ʀ�\���^z��X�� RMnx�U
��b�~⺝N}n�(�	��J3e/a��"�].�<�@� ��hd8�T���j�۱lش��E�^�֟L��L� ���UI�,��,����B���T���Gz�O�4��w�Il(�D������}]�l_e;���< vȞ��Jy*t�k�o�~,����@��J`E�:\Ҋ?�HU!���S� �a�t�5I�G��kd:!�#�ZT�6�������-iץ��&�^uN@>�m)���+�7o��X�ۣ0�1�&���L=��{oST�D�(._y�8�q�L���/�'�R8P�C��(}�'hb��52��hpA핝�b���٭�G�i$�y�@κ 3�������*~��b�8���NG]�6T���[<
&����FP5���"n�l�*�����,�������8�Ѹ G�� �PT��*��vV:%8aH٦STs�`n�G�Yls��Η&���4�-����{_s��k��}9�[gzFé�	ҝ2O@��(��D�B�}�h�l9���)���^5�]]��ޔb%��m�Kk��pᖝJ�����zA�_��sΈV�O�D2�,��W	�2��+��n����G�q���� �;�D��cz��paI��qLL�� #,=�E��l����!���(�[uulJ1I��]��8|Ǌ���O#ζ��΀9�7����h��A��H����u�/b���2��tل��ت�pi2��^�>[knh72Р���c7����_/M�a޶#�z[Q]�5C�����4N+���?��E�yJ� ���J8��2��;�|3�n��ڸ��Ӆ��W�Nd*��;��O ��%.Ȑ�'~�����4)��6�Mf8�����yl������%���<X�N�C_��J��>��KQyE�� �ű�IHbܖ�޻뱥�y'J���i��j�^�a3`;oi����h�!q���C)X���i9i��^L�#������ib"���E�Eq�V��I��e�9�� ��l�E�n�����HQaq7�f�¹pXA�_�cl懥^�j���F�B�uW�}8NLҲtm؆�?���4A�+U�#e����.��d�dY�
%�Yw�:��v'O���t��(��
Kg�>O��V
��,Ù�H,�lʾӢ^$���1�J�6��{o1D�dP�A��fUJhVlL�t31p�ĢA�tQ�����'�_Ѻޔ4�8=KA�P������9��Zֱ"I��_Q�u�L,�!3��I2�Z]���;�՟v����B�7G���3L���ZI������.��>%yڣj�W��_�{
�����T�S5FDE.�y� 9��Y��oq�/�6j��T�nWrk͟!��d٪1�W-�r5÷�,z�:�n�`���q-��vO��?>��5�8kT� �Crm~U�j���j�Y�-��ȝI{;|zQՓ;�-�B/+$�O��bo������&��|:���ݑ��[�[���cTob����/��;Ply�cr~.@'D�s��x�Y.F���l].���b'hN
��a�5�9�XTӳR����J����Q�t�6�官��su���z����`�>���;�+#�X���Ɖh�eFj���Ѕ���qi��٠w�y$6��J��~�N
s6�O3�F�m2��K;��b�ƺ��&�:C�*�X�N��7n�	`���x���/�V�v%&� Y�U<�Q�ܚ���"�*��u���W��3�c������o%��b'Q1�Y����u�5Z����*���=�"�~H[������3��(����7�)����cԕ��$�
�~�s��|J��FҸ��:�w��X�V��" M!U;1�6�q��j�Q��p�����,�e�xR���������w<3?*���=��JdN��`WR|��J����xB�HҤ���I�#��g���V�V����FkHqUkC���P-�UŶ^�d��c}��%���_�]��d�m�^���Q��L� �e���%3��w����zz���~��������O���W#e�,�gmP]FKu43xu��Ȫ�?Ը�2Hp����d���<�0�ͯ�c��L������qj��BB0��P�aH\3B����Z�)���3�3��4���| ,�B�L�ߒt�oeY:�]0�~��(2���6p� �p�.�:TN�X�3��>�\��~������d&�9���QZ�d]Q������%۷�;|P��-���a��ORU��
���-A�śϵz���X�^m�n���&�>m�Ŗ���`xg��:��Jy/[dB0ӅL ��f'�w��#��V-��T�w;s~��Ju^���E���_Ң���ҿw�M�Q7or�o�z�����-�
TR�J4ذw��Sh��U$GG���A{	V�zǐ=p�}�����F�Kϟ
�u�Uoե�����rJ����ޒ�>�f-g5@�|{2�5����?��E�����t,�l��`�"�l-u:s��e6Ob⎼7]n+�S:�H���7f���'$���,GڙR�Fi���Gg���Kѫ��D�Rb���Z��[��v�?ykИ��
E��Ba�(HX�7���z��i��͑���	B�k-�}߂�(rs���!��1��?
 1e����+�X`��N@�\�݉<�V�n�WbЉa&��MU��<��e��[;J�u�v"���}��͇�ڳ��T�Nl�5]�(����G@ѪP��^����a�~d�y^�d,Np��|Ghk[��ԥ�մ�Gf�������6�,��
�n�|���FE�{�Z��	��C�x-�����#�[i�J#��Z*�����b���\�Y1 Z���J��2�Z� Ǒ��E��k��F��[ %2WZF*`f
RQX�[O0�4���ܫ~%��x�\LY˜��x�6)-��vT����޷U�fLM��1(��ur�RaR,G�c7a�B�!�6�Eo�WH"y�6�W��&�`�1�m�����0�x����k�`ƄL��^Na��]�&)�,�[�h��ғ�Wx?MM%�7R2��/�'Ё�>@�X�C�>�a@�ÃQ�V�����oyDz��3�"�U��}p���$D��Xox�B��LwO���6f��'��Ej�'t���vB�|d?4����"����G���.��n�G��Ͽ1ſ_vw���lU������i�sI�1�N��/q`�z���Ɲ"��v*?=l�D���� |01J"enb�%�w��S��&P*7��� ����$8�sy�kd�ܿ��ue��x��:
�@�����A4`5{S�W� ��mI�jN�`)(}k��nRoK=P�^D�z*\���A��VD�s����L��E�q��%�
Y	%��/��j=Hy)�L���c���Oo�N�;L�����ü/!�8�\�n�k~^�),�Y��ϣ�9r ��X���,��N?c�&,v<���HHf��ߖ����Z:���&��g��Bw��@җ�_�OS �aq򧘣�w.jC�������
m0�ܒx`ONJ�R�u����U�}#T����>�FU�# ����n�w�?��� y��?�H��Ὅ�6���>G�$	�v]B3�#�ga]��t%� H2#��Mm�߄Jma�Y�x���\��H=���܀�Y����)�p��Λm�Z�S����'��K;sBՔAP���*���-���0y�8ٺ���%��Ő`��O�8O���G�<�.��)o��O�u���"���xW�n�z{9L�t�f��>���.|�����*/��?�z����1W���$ԡp�Ӹ��"ꃸ��Q��f,��w8l�Ԧ(�V�C"�0O�̭)WK,P�Q���8Gn�ϡ��rh,?w o\��w�����1�k�:e/�0YD�����م�ރK�>5�[��9�^��/�oU�3[M��c��A�+@�JY�m���ۀ��a �vY;0Z�daԠZ�첁���M���gb��$�����ڒ�t��D��)ۮ`�N�¥d�7]S�����M��A��t!3�Й����g��U�;�pG��B�%=�%>�1����W����9m]�$p�xd�Q����C}��em�)G��쥕�~kX.��Ò8���0�`lݍ7���D��p%�ʔ�|�YX�A������?C�kD'>3N�i��>�L.!"����&�~��l���9�\�YXF��N����Ô����9�']۰����ʜ�>-d� %ds�]�q'j�%��r�?̭�����H�I��;$+L�^E��n���,��C2�����.l���I��+Ԅ�Y���4��3�p�%�\�O��X��^��!�d9�,$�����&��\B�)b�id�S�J���[�0�6C�ND�ll�W��s�,0�i3�oO�R1���E}S͜R���5�N�g��a\�,�R3O$ޮ}���'NF��M���-��0��48�p�4��f����(��=6O{�w�öa��ZP�lt�Mo��<F&�RA_#�}���m~�q,\�e��q��M�iUD���f�j�w�@�&�˪��D���w_���M�಄�ΒbDް�[f��ط�ۏA�;J��`����a@��@0k?M�!��(y�B��˶��eiMO�tr����!�:��L�U%���/o&���3�z��"�?��p�dK��� �z���2�Z�$�С��HF�4���8�R���Iwc�|=EjP�0���p^���q5��V\f�[r����4�`���h�-�=2���$u��y�X�z��Z)��()%�z�A��E8SF<�5��IEo��n7�N��4��W���;D��L�h�It����Jmr�j�z�ߘ¥�D��y*�K8����h�Գ�U�Z,�cI�&��Ͼ��s����CA�z֐Ф�uoK�_��bU����Ɛ�H��i�
j;�C�ܡ��l��Ǡx�n��:yk0psmCL�ɾr�2����1�e���t5XԽ<�k"d��Stނ��[*��Nz��)P5��Ă8�}-���'�7��e��C���S�K�A�8�Rg�jӶ`���I�*��͐����PPn0�z7k�ډ�"S�0l�X��r�-� ��PҊ:	HV�(�Х-�W�S�[�J�:��<�u5(S�$VHr��ꋈ�����TM�9	M�~i�a�&�������Wb�l8�?�m�%�<Q��K�y]��ㅭ�h��L�,J�>�Sp��++�cG��<dåQ�5����}������\�ܖ����Y��)�`���}7�0izźק���g2�mO��X&�1�P��{�Z*ߟ8�0ڂ� ��^I�C0�H	�����l-v���|��8��/�^�K�p������r�0����(_��I��8� ��)����Vۉ]��!��^4�L�쏱��⏳�K���Q��=�v��{�������v��M��$H��<������j��@��q�i��n�����yg����3��T��0��3$$u<��_����>�I畇�����e��I�[1����Y��5��r<̠5�4Gt�����OR�{<��9׷^Q�Q�R� J��V�ޜ�c(G�Ά��ב�E>�yk,f�m��A�;\���~_���.��+��I�2gmn��񎑈�<���:NĚ��$ �x/$0[&�s�O�N�)^VWV8��3%.�|5��f`�4)��.� ���
�~໷H2{e�>~��eg�:��q��!$��l�b�猷�֏�K�i�G�6A��Dڝ�R�n�V��_�rG�Y
�Ų��"�����Xon!��	ŖW�u�?ba��0�@�n�9
�w� �ǂ��X(�`'\�|� 
	��H� ������}��l}��D�F��R�+^:zv��kq�$ܐN�7�K	���~�<�:H���P���d$���i�G���9� ��A��}i���v<7�oCS
L\vK�P��.��^uZ�w	1d�,kC�M�+�t����!�2�?f�q�LA��3g0Bpq�2�!��C�
i��r�ƇQE��F0�Չ� ����`4�M����|x����u��UV��n��ԁ)�����
i���>0�I��%��T���c�"���$�_�2ѫu�~�Z�-�ʥ3�.^$Bag�tC�k�$�y�Ku_j�*Y;Ц���S��{!��Sp���	Eͬ%��;� J��Y�u�	���f5��?��@�z�Si%� 5�S�L�9�X���|9lz)��d}��a�ǆ>��8{[6$�Hƣ-���tM��Zlr5/��=������so[�;��n��m ͱ�9�՘�3|][X���s"J=>1�8Z|�[0u��ׄd�����؞������ƻ�C�'��R���S�1ڕV�������H��Y1�h���
��?W�A"�Vθ�;QJI�d����*
U?4��-�x6�go��uqp���d3���j�� �֝�͜�zU�@������w���\Cjh!r��,A�f�U#ċ/yjϟ�<��$�D���M������Y
��+��uy$T����f��d�F�l҈�;���⟱�i���]A|�yI���n2�b�_a�p�]�p?�MRm�>�A���.�Fm��i5y�䎼�oky��!dLZǷ�Ђ���	+��
Eغ�-�va8|GL}e&�c�S�裠U��EgQ� *��xu��S���A=�o��"4���Ԫ��+e�I�]z��U��c-���6D[�[����Q�D3��q�uȽ9����=6�;�='+����M�ٹX���!L#����n��T���ƻje5R� {N�tr��G{4��Cp82,��4e�AL�-D!,SH���e�o>Ga&�	��3�b�'���̓��]B4��5��MXl�ߡxh�H;���§��!����vN�E6%��%����╟�g��	f�B�#�3JHܬ��o@�?�!qj����w�{l�e�1/E�2��fv������N����ຶ�gd6>������z���ݕ�.rX4w�;��_	'FgtD��s�H�륃�j4oe]�ßOSl]�ɺ��M��x�Pv�#ʓr����gL�-��/0�'�_V��z�����=1d(k: 5�>�B$�L��.U�(>ь���ΑxዸdW.��g���/�)��;R�H�Tg��I�!���m�B!j"�y���a�v���nˀ���Tx��T��ߥg���yR_k��oy�Xyl*�VI�Aܚ��S�p'El�Qa{ԋZN��0C����RI-,r�JHG�A�|�8?LW-����E�N��>��4+�HWf����+�8|��csx�%��e)e�-ºoF�����m�J$�J}C�9�5G
-x�������yV���Y�J�<�p߭h��F���`-�F��:<E#�d]A$B� ��d�b��k")��׮N�e��G��D��	�����s�0���7Փ6,�2<����I�0K�����(�����.LS���(Ǚ���b0#).`R�U.ܛ7��<��i�0��<U�PR�b��m�b��$�bH����`�iog���Ҡ�M��H0��{B�؊uDv�,7�ә[�5P���jT�"�E>#�0��!2�&o ����&?L���Zy�_t���F����a6��>���eJ0O��H�{MK��@r�j�ȩ�`�s�"�v������Q����r��!�h�ϙ��j��:Y�wyg��T@�ҍ +n��6!,Qjf����$c�:]bnGi'�<�R��۽u�$��"+5����m���i�+�9�B��]	�bRL�Js5��08����  �V	"\x�d"�O����s֢�#+��6͑o���h#�*Z{�1�pΣt�i�~B<ŋc"�F��׾��W	��h[[������>︷����F�*�q�����	��,@���d��hDv��|1+��N<2����d��/��X���u�R"ނ����'X�i����Y@H�d�2hu�u����Q���|���z*,�N��P����~��}���d��bBV�	Ō.(��.��� �7�堰��n����{+�K�^�SB��5��jc�^�tR���u��	&8�]��:w���SCP4�̛N������]�J�����)�W�qO�QSv�K\k���F��"4�B9� .�ĕ;��Ol�O4�����#2C��jﰄ��Җ��9�1NUp(7~x5����?j#r���==s�@�T�����HpE"QD���P�:��@kt��V'��_�����e�O��ݩbe
ne��k��d��> ��w��	���CY��יX��,�~}#���Oy�}�K���vc*���D�K'���oǞ�a<(��n���)�-��T��䤺�7d��_���@��>�j��P���<��m"��#�_�Of�|e��&t�6~к�&�(PL��!"?�׏Ά����v �E��l�YBp{R�ʷ�����ȹ�L+�%��5�SV@	]\��2���r����8*��o"�TЀZ�\-<L����m������ˎ��Q�$. ���oA�gقa��j	M�Ö�h��÷:��Yp+
'�.`�܁X���e<�(�6�z��>!y�!=_:��k�0�	��eA��N5�4f��yɌ�'8�R/c��3�{��B+mD�7���~���d��W|xӑ\w����u�w`'�T;B�mõ,%@-�:�O���_�*��.*w����گ�@̇?���C��yg�V���@ms���U�E�Z}$�ڼ���,i懕=�����۷Nn( ׇ��G4-��ϳ��TV�b3������r�'��O��S�RkPe��G������*@Q�HM�r����:��M��;`C����MM&fbm-Kd:\*Qk[�����/=+�3���^/R!,�٘_�a�dp{n��4]�Psf�@�5#���QIM�}�Y��I�do�ݞA�<\X�d�\"^�o�ZJ�`b~��2����y�Rï],0��S&��v�ۊ��=����.����7�l��L;J�w�_$���W�Mޥ�x���yó+��Y��y��T����^o��}ũ0��Knm�[�Fi���+#(�=I0'������Ļh==�P�I䏐Sp���Gӂ��`�*��b�� ���>+��T�ރ�E��Q1��Cٯ�P�Vu���j̍�n��z&�˔���æZ�[o���h�����0�,�_�+w�0�=��.9>�-�o0�u������C�f���*==���W�4���%^W��H����w�����7��zY�?��L�iD�$�o���9�h��u6�C�d�-��+�*h��+U{H�£�,�	����|El
� �T�^j�c�ב�v$|ſ)�.5֗8?�-�*ro�6�S����V
�_�""[�����M��W�\��.� ��d�ߍU
���a����lZ�nXE��8��'c�}	S`�����y֑�.��á�UC�y��2��t7+�G3Dؒ3�����e��2�}`5&�5v���3�����n�}x1#�%_����z\hWD��nBjn����T5��e�{M��#Y��Z�H��iY)�G���_~�ݔ�� �MӹM��q�Yb��#JY-oEz�.3�į4A���bE��!'?yv,QZ+Fc 㲔���#�Em$�'o��#����h�u�i*1֤��� ��oԍ�o�^�6��;���=x�>Yc� >['"���0��a�;�<?�o�V��md-y>�t�Y������I˅�����(i���l�xx���-5Jf�1Ѳv��%j�%-sƕ��J��e;���_ ��2=�3�{��W;�Ɩ��֣����-�F�Ak�i���]#ߖ1���<UH/�� �������+�3[��~���h��q�6�D|N���؄�9J0h�tYy�i��u۲ L�'R���vɡ���3�1�nF����S�7�q��҇��J����A̿6��HF>��w��z�
�w���{����&DR��@-$��y���$%|�RR؛�s�w��0Z�&��{�� p(�D
������
g�
jxȼ~�C�(�p��x�X���R�W�"sk���v�W�ƌ]g�Ө� �5G���)���o]r�]ꕐ��Mq��¢��3��L�x�M��S2*���YyJ�Y�}'�
9������l�7g��g�^ץ���_1eF�"��Aۻ���X�w���-��{�Y��ĳ�Ry֮���s<<���pz*��Ao7��|0Uް�3`�?�=��;��OLmF�̷����x	͙��9(dDGF��0\{q�>����c�&�ZΤ���-*ec�*:�ٰ�DO�X�@s*2y��6
�����͵���Ѿ5���y#�7�^�NL4��� hv��D'��#4�!�(�F����x�#�o�kE�*��e���?W@�k�^4�֨�Ja��d�t���7��:�W�ng"Rc�?_���.Zfl���V���εմ�F��FL6�h\�>Ǫ*�!"T*�-�����"�x��R������5s�L�5�\G��r*� 9�ň3�BH�2f��É�lX����0f�1���K�30���" G������S[�E���*@u��j��qy"
�����k��Dc���+҆���ޭR���}�KE�(	^�R[��Y�$د�Pg��#�ۥ��׍6�m�$V3 �6R��&�s���2�8e��9�ħ�{vJW�;ܥW��X=�!�Yh>Yg��HY~����[F}����ۈn/�0=��f0M1�'���2�8���P
{;�% ����YP����f�g��GhWƓT���cH�ZPc(���<��Ԓ1��M�N��fV8-�H.�f�*ͩ0�c-dL)�[ B3��s�WK���Yݓ�n��w�i^��<d~_O{�8!�@f��РNmI9���a���
�֡��~�����*%�tr�J�`��S|Uש�fL��~��q� ��A�>���l��Q��<��ˇ$k�bgl]��f]k�]��eTRk�Z�Ȟ1~J%}��#��U�U*�E%��d5r�YlK(#F�$p_�5r]����l�3]e�Eb�U�o�EGI	��F޶��W�^�j�K��!'�өMF?�̙�&o�1��\�8*.���׹n0S�N>ޯ�F��Qd)!��q�c=�ZWN,�>��^���S��.�
�h)1�(�H2V�*i�X_"��5�[e�dĆ��%�<��i	Ap����+;1�l-f�>(�j�� ��|5[�̡��o�������C���R��jp���}5`�}H���E7m��w޳���,M$$���9���h�vmh��w�&?���BfJg����
�(%�a|n��-BÖ�;a�=��H����ԏz��)�d{��xפ�@O���饫z�4�S����Ӂ��1� p�#�ΣÖ�}X��{�� y!�y�)����:��2���U�ӳ��,2>��Ƃ+�t�.��]��xZ�9\	꣨GY���9�͇@#�Ⱥ��\q��+�Q�,�i��(�s"m�$]�q���ZF�Իb��_>�'s]`���h�C�"4V-�~\q,]짲)7�FI�{f�y�t���Q�,�kr������*;���=� ó
���b�k��2O1Ԃiْ���=�_վ��Դ��9$�����8�E�{�q�CjV�t��
*�YN	��|��5�v��٠q��9�4�7fD+s��bF���{�\��d�L|�Ƶ ���͛��0R:�Ҍ��@�,�U�nS�^��׽_��Z:���T��
x��_��C@U:�!,#K��,��;]��&B/��Ǡ[Ъ�2j���ϊ���pu;P=�����D;3����x=}��*>��ծy��W[����D� |C+9R{n۟@o�gZ�#>�n�ɹ����V�$-m!��4l����D�C��yx�]�,����,U��wx��Nf"�?,9C��b���[߄�����8�/�Mllcӈ��z �V�Y��3�5=�֯� zISɛ�%�s�� �����~��XZv���`w�l���5��B�a�m���(b��@��E(O	��ޏ���M�F�P�ǩ)�����Si0m$�=�1#&W>�@��@8��yo��F�L�螓�N.Z���	�	jZ��(#��w�wC�D�&�� M\�p����s%�$�1e�ڛ|��%X�p��Q�/��B�� ^�`C����f�w����Ֆ,��ճ?��j��)EY6�+e(�u|��R�?�Ջ�$`���cV���MK >ŋV?PJ�څSƆ���=��Ȣ����qp�e,V�Ӊ�_~kk^ ���tQ-�y檐�'�h����#8��.b�<��g(�Q[
�%�q�Q����M�2o�I�(�#�ool��h<����:3Iz<�-	7^���3`���e?��cΏ��k�b�B0��X����J�5�jB�~�_���yv�����Y�a�h[1(�n���*�Aɼ�v8�|>L���>�����[@<��l4��h�����%\Ӫ�E[��P��|��{���\��vO�L~��o�7Pg�\���������+\����'�����:��p���D��?#���t!m����H��=*+.���I��51af�������a����y`Ϊ�O��޹:���ljNj���'����M#��fD�3��kN�^�hBj�a<�ʋ{��]3a�蒻9K������ ������?Hʷ��'��s�B��@�p;���OKŉݸ�ҡ�:��P*�o��@>h\�<7v3;3f��� �S�M�����ϡ��յ?I�xBōo��

+�� x�;�@�Wʷ�/�6R{,��')�N$�>O��ƂP�T@fc����'{&?�0+3�0Y�&*�xK�;u��w^��B�/0��J��_!C@�oc��G�Ms A����Ϳ��4Ϭz�t�G٣t�"�Hi�`�~E��wim�|iF���hqJ��1[4�rFP�Lf�
xa����C�yt�t}~R6�I�߾LxX�i�R���틺;,� }����<5�[h�Y��y
b�cQ����ǝLL��`_DH�P�荼O����s����>U�o�1$$P@��V��I��ϴ*W���@�Y�^h�ӄ�����3�܈��Wɶ9��7���dY�B��j	���+�	{#�t� ��ާ�G��b�E
�'�D|0��v��sI��^����䉵���<�������~ȗ�Y�!_U�'�4��l���<B[��6K�{�ނ�uP�Lx�Y��C�!_"*�!�nN��<x��&��S�u8�VnN�k/��9���m(�Y��x�9��ռ�<Y{썋	,�o���-���v4�6X�-ʙ�E��}թ�jE�I(�C3�i�ܨ���N�����V>��LK����sX��b��S�{9Nڂ� +�R�H�W�ߒ��.�j���I��}��+╧h�xAnI�to-۾7V�c�f��m��Y�:P����((zA���m/܍��ͱN*��K-������$r�ٴ  ~l��N�]y��R�O�Ť�K�ôR��fB��v8�1%�B��*T�c�"!�hn�� �����v�D��z�0h���#�킩��`FA���\%;�l�f��A��cO��,l�۹U^�b�&���]RoHX� �����F���γ~I�{*y#���4��[ca���N�4[w��=Q	g��Cz�L&Y����v3fdw@N��r#�=�L��� �Vo��',�$f�;�4d�G�X���_q�<B�L��2��9��n6[��!ϸ�{f?��y�_u���CtLp���:��C$�eIr��~e�)at����U��)��=
k5�g���"��0��8�\�~a����v͒�^�̉����g����zhxv0U|���~����m�;���>�Y��t���K��y6K�}0y>EvnI}��{F >��Mm�U�vLi��E�G͎����������ϴI�5���ᵎ��'go������LG�<�U~P�����NƔ��:)��������/A�g!?o�6o<���p ��UN8�j�����K����L?������)\�O�Yx�-Z����Y��?����g.�?l��t�.��24����V0�Q�J��r��b~,���i��]����͕<��"�ls
���`��[�
�c��G�P�{� ��0yγ����R�5�-���;��9��f�4�z�R��En���^k"���:��7���O���c�+n��"�u��dq�^O�o|���l#E�šunI
B���;�F�=��'K�$�y��i�����u��߷�.�t���3.���e�ѫ�ڌHl���ưa�0�T-�ن^�$Ϗǁ�B����"�\/
ɜ�})�����."{�≵)��Z�#�L7�xˤ��x	�,lE��H�#����=Q��C�tU?ppQF�ٝ�"s7EPn�}����pc�MB��(��vJ�ӗ#s�/��!/B�4*׌��J����J��զ�i�'ǵF0,�Z7"t�t��5������.~|hA�����N�ubG��c[����',L[p;�Yߤ�\۪V~��cZ��$�5�$��]W"����1��J�R����]�*���z�m�q����xM<�[N'=�n�Cɗ1��w�6�+�F修M*��5�H��ۂᴐFQ¹Ih����.�6�ڝ|���U���E?ꢽ(7r^ѹW���,���
�H��h~��x��)C�Þ=�T���X@N�/��Ͷ�l�	�Z�]�::Q,�p:�j���"Ī�3�v��ln��r�A�o�9IP�eN�EכD��dB����!�:�j�b}>��s��11�+�r"ăC�BȺ�!c� [���& �9��a-�~VC�'_$�XR*�h���"2)�z����M��co}��L�,�Mn]���`��m^T:�l�k�is�S�Ƒ^G���ťנ���/��D3�6���0�Tֽ�_�Ƒ���
�u�O#��A�b���=�;�s�9J�=���j�'<fa$�	'	���T���LU�.�-��l�"�fE��LȪǔ)V��KӀ3�<`��R@ j-�;��)��s�\o�ziv}o!���B��f�_5�H�1�*�2�-��0���Ј����ɩZ:w}����X���[�<2�ah��x�0�����^G��2�r�f9�E��N[-وw*����D17�n���P�|	YNَ9I1�I[h�>�"�-�9��{o=���md�`-#>~Z�;b����B#( @����Cw��E��ARv����a�!a��ӿ�T+,m9/.b��1~x�����߿�f ^>��K�}�S��w�Z�Ɲ�V�<��<�ʐ��>5�eb��b�6�1��g�_d�%^?�}i;��у���	}���j���}t��]��A?-@��w~3�ɤ'��&����#���-�T��6X=آ��Jp��#jA(h�:��f���y�Y�5"��>��[d�I����d�)��������p6��"*5M�?��R��~�;��VXU1��4px�d��!Gd�?h]b���ql ������G�.��бr	����;Z�M�5ڪ ��P�!�U��̂aqE(G8Æ�)g.��{� �w�O�.,GMV�^���O�`��טㅓ�����F)±�1'� ���쓡�e�fG����<�=�2PӻH�'������q��K�Q�۬뚼�?�l_�fClw��'ڤ� g8�h�sŤ:�,�!�х`����$�j��H��A�ۣ<�a�����Q�б��5���>�C�vR.7�R�J˲:J��q��iC370���\����x����$%��W�7�.!U�9���J]�u�<�R�L囏�y\X8v�l��{�`��4ĕ!4�^����``��\�����Ka�[�n�4�WZ��I�Gۀ�j��3����AO�޷�:hkZ�e�i�0�����͐8�2��K�D�x]xD�XA��Pچ8	cdJ&�� ��%��JZ~0��t��mp�4
�����6�ݔ�y�ፋ"����վ�pw4����:���si�������-n�&?�B	$�_�)CE<�ܶ�	@��F����J �9~�b&�Jޓ�1c67�q���z�����b&t�&���D�r�m!M�����L��٫���K��������Y�%l��2���H���9��3��=��?�PLS��{ �@����*0�m�����nU��F��oǜ�]�Hꁿ�#[�qA!�9�K��M�~6�S���@��9sl�՞�T06����#	e�J�Q� �5�����\����!�6�L9FҞL�hx���b�������I����$�L�	cZ/�2yԈ���8Aj�^P'U0ҦAR$�| �TA >qY>��,���R�[J�����a��[{*�8�DM۽�Q��;�]׆���L��A*�Ѿ(�"� �/{tP�x�����rXż�m 07�E��R!�j�yM�?gFH��G��hd�%Ng0��ꨐ߰�:�`g/wɢ��C�@W����Ez��A0#yͩz�Dg����xKھ�����g�pL~�Иu���:?�V��){I�b�&�����us]�S7���s�׃K�������\��W� T#		n�5M۟��+\O�7J�o<C�28ȅ�N�����xĘ�6᣺tU�7qAJ�!��P�$Ҭ%]����I��������C��$Ԗ�<��1[�$��v�����4�d�� ׁ	 �x�gy�O�d�p��o�q����+�,��;k��lt��MKB�K=8!) 
Ѡ�;��O���R
��rP>�2�>�G7�
8�)����ۦ���[��rs�o` W�#��7���gC2v鑷��hg�V��9�wY9�H��1ń��% 5}s�pq�+ө��Ɍ�/N�°R�P�*���ʣ,c;���"uh��	�Ö���~\����)����a�i�jڲ��Ä���^�C�v7:����7�o�J±5���<�LJ\8�y����d3��s�k&Sg����w+>��������{� �k' ��Ɉ���R��S�8(����-�y���?�V�?�7Ev�C��:R��Ro,�?�R�'�����>Q��y<�c��\�<���	?8�f�ݠ��o���x*>A��7E�X�����9hd���e��*`s�wAЈPf5h��}U�u��1��U�o^´{�EE��J�:S���7���?)�H���2��B�i�P������ %�I��8��;w�ރ����]Դ�s5��*���\�Co�C���oQ���p��/��ȕ�Rs���t-�mVj'g���M)
�Z��,F矅ȓ%��x^s���E�Hu����<K��T{j�C40��^{6�{i�m��!����8�֘��~@����ZC�*�d!!�����������7܆�����4�Ԧ�l�%/}]��>O��g�s�k}�#h��8�ӻ�� w(d�r؞��Nr�	����;+��AEO$O�4q�ֿ���z�����f��:�)wd�x����r��Z58�G��L��e�X���4;_/p�#��A��t �B��*�`HrWX>�@xh��"�\v}�)�J�z����2n��-�m�{��iWyQ]��6��2Bc��X%F�H[z4<���\�(ס��ب���y����Q1��@����=��KB61Y��V Xy(�kO�	8��czu�질���$/83͔�Sn�>��6"��ڑ�q�p`ڕ�h�����t3
Ss"���G�0%`Y�&�ϝ�� � ���[+j")1���6�T.�Q�bx��(��~ozs
3ˤ����x�����gC��	��uSUz�	/_�;d���������cg��2��5�
�&���+׮�[�T����*��<��Y��G.9���1hVTѨRs�(?��(7�*'�:��p�kF@66+�rN���}��aS��V8��Q	�w_H�
�h�iJ���E�.�}�REKZ����Q�z2j�ucºղ���4/��γڟ�Aխ��q�È��.9�� ?�������<���M��2��.�a��p~���,^!l6�e�r/x��<cc_#�s��H�i(�����]c#2��=����$2�)��|�xxE��H��J�k+��x@p�llY��f�+��R�w}�Rc�m�:J�k��@V@4R�-� &��~�N모��a���g,]h���g�`ۓ/Ԁ�����^�]�O�5��.f�m
�jnǐa�?��/�Z
J�s�|C�(8�}]��KC�U)7�`L�����=u�oa�������83V�ڸ��ل��2���"�,6��6z��n�,�I�Aa�_:%>W��Y�7�����������&�&j�sK�I(H��.Uϙ�L�i���3]��_��^�(�'2qqF�)-<��V-ّ4�×�$��?(�)v�Zk���$�'�9�B���W6ܫz���j[�H,U	��su|ᷱ��4rݚ����}�UO\X�;�N��J�-!$�xԳ���$�M����?a�fIk��Caƞ��p6������G�9�Rg�K��Pã-�ZթTԬ�WR���@~��{�'�C1��k�3K9��1V-����#�%��A�u��k��Ag;��8�<������S�N2�B��?�*���+�7wY>V�+���#/��X#"��
`0�cJ:A=l���f���Y8G���c�� �|��݆lk�l[NQ+X�gS2!W�f~���@7����z_��hsY����"?#���v!Q��x����߲���6�9�u͝��@ٱ`��&pU���������5��i0$�u�R����>�܆��G�/�.�G)᰻���s0�M	nܭ���.���OK��������e�!������x�\h�y-S��579���Oއ}.hϙq�\B��m)~տ���/�u�Ä���` ��s���h>�~0����a6�����KC2mA?�QD)��qE�k�r�"����_��n�X2���ʺ�jW���Hf:ʊ;���$!��jF3���j��p��pn2� ���v�C���%�����iX����,t��墙�N��+����տ�7�s����A�:d�H� a�m%��y�v�g��c~Ys��w�Ow���$�'E�Q�+*�*�ު��/g��3H��@�����JT���|ʞ��>Ӳ�GI6��&C��=�T��C��䵇�m#�Cs�ۖ�{6��$��5����'��HYjB����f�*�[C�ߎG(�3R*دTtE��5S��}X�b�����/�qׁ��� ���<,�_�6�~r�@uڗ$�����w���G�gHr���*���c`��M:�
��m�&�����S��Ƀ��Um�-_!��3}:ڍ�:�EVWV�j 
��L �/�REt7�i�a�9��N���e)�7�U��%�����$��c0�����B�)�.����o�T*�ux�4���΍�ߺ*�m���\�M��$C:k�BHj�'b'����G��O`�rp�ݻ����>��.���F�F�+#�����ί�I�f�ۃ�-0��U��>�
ɀ(o	it��E���M���3Za#�,�J�Y�@6R���$y|^ǅ0i��{&H\�nE��k`�,��HT*h|�q�'�����>cEx�G���y���?6�v� %L��6˻�K�7P�(w
@|��B̇x�� r"e��#W����r����ơt:�@��N-0O�����FZR�WV�G�>k"�H�4�����{_*;c@!�m��ݠ��������KXN|D��XY�4��ö��c�$�1�(���Je��фD`��������%�[\1�Am��.=~x�(!'�Q2�'��g�ᔶ�CHM53�h�HG���X-�@Yn�	�=�ZCnd����� WƉ����[D'XC�N_d�&���`)���v�ꏾ]}�����D�,��"V�6�����ྗ�؀){WK��&b�2����Yr�OH�h�??g��TI�P�0�d�*W������uF�r2�3xi�2���h+)l�Cڂ�H4v��<�O�l��d��c�=�R��ݦO���Ƿ虬#�� U�$
�`��M`�w�Q4���p~6���� �9�5�-�G�w:�UjA�e*�{�T��혧�s������|̰�|!-��� �R�p��.�j��<��nmP��Oe�F$������k���G;D���Q�tkQ?K�5.-u��J�H�б����c\r���̥M�G���	��X�l�	,�vf��F�@�>Ǧ5����7������;	f�`��=7�x�;?j�<�Ey�xQ©r?DV��u�e5y�>055��liGH���Y?�?"XRr�$���ͥ_+y݃�qba*�����Ûg95�̙B�~LsE9���Q�C��L(�r��)����A�GO.�0L#��h��~tN .���]����#+p�@����>3"
��>���ϼ92
>Se�h�ʐ��Nqי�!�j��_ǩ_Tt�d��%�"�S�,�Tو�G"�a�����r�Jk*C;4݄T��1w�G���4j�J�� �q�����dii3p2+s8��m�
�v��T(��>n����籊�������@擙���ŵZ<�dybCR.T�ʦ�N.�^�{[~�4�$E��`����aF�{V��p�/��!��$7!#S�a���O#�Y2�/t���~����#�K[+��Q��b�;:�i�"K�'d����t��4��R?̔�r�� ^������ܑe4��pҊ����^���uo�KV���LBi	Ou���&�a�
0vy�lR:nAԮlO��[K���u�ɔ�2w�KGn��?Y���>�%�e�Χ�EK&N� /J궉��3&�eæ7���#��� 	U�Xʇ�aA4Ő lZ���9�#;�v%osI[U(6�(��Zyv�$# ,�P��m��#p�{)G>�S���^��n�!)�g�O��ĺ�hw��pb)�;�q.�{�{N������:Zv%f��Ÿ}�m�=q;o䈡CD����z�����L�lR%����6|�_}��:%��}~S	<w�E	<�ψ0'�;O�(�_d���ɏ��)`�o5�-��� 5�_����|���e�T����#Bp��,�\�����Fv��ˎD����Ў��A�wi������.�u�}˩/�ǃ�/�Bp��e����s8�R���s��%�T�:A��.�;t@�*�Q�WkW%�� �ZŅ�rg\^�l�G���W�
��wu���j6��8�E�1��&~�E������X �U2P������@4~��}b���Ti��l�ԧEBLf3	��1YY��j+��_��*�\g��(_4Y�1�V�V��k�f�n�;�W��^htp�ؘ�G� ]���)|�X�n��LΜc�	.h�]�����x��{7����ò��iC�O�p���F�`�2�bMA#�#U���j�J<u�vFZqV �$�Q<������v|'�P<&`��dKg�[z=ƴ��[J�s�!����{�+^2$�e3G� ����9�\�����J"i��(�������qNE֊� ��633ac��ၘ�{
���_���(�Q��k¯�C �����#�
rv1�9n�%3��Z�5�����%�A��U���q#঱�L�5�$^-�T<���Q�@G	ַMWg�^q.�5Y)�v>�Ƈ�!���qZ�:�m�H(q,�(���{�>��O8pX	=Yi��72�>��4YMG��'�5�,�[;h	O��jThX�L'5���G�$T��0�k�d��K�W2�#	C�/2�QR���E�?�k�V<�����~�;zpH:y!l$��+[��;T��79�*�R��wӳ�_ܹB��:��,NI��Ư�3���ݱ�.�K�,���ׇ���Py��%2��#�۔(y���8�3i�_��[e=��P>#��v�i�P���wpF���;[�ӯ����T��L&䧶Y�4u߽؞�c��SAܩꤋ�c\x���ɞ̷Jcw1ܣ��J̴،K�y�����r@��&�d� j��7/�. T�3Y^�Ґ+ࡋZ��AcAb�Ϋyp�O4-�"�R�8vM&�+I�.����+&�����(���!�%�o��b�?p>��;Wc}����%QY���q!���&������g�#�@S�=�؀�#�
�&�x��($�&a��(s��o�} d�P
��f[��:þ�8A5�B�d�~��p0fB�7� }_�J��i
'5j��C�a�f2K�&'�X��d�,�����+i��.�HΥ��� ���Q=���"?���)U�C(������8�0P�����z��Ʃ�r�T�ns����E��Cj���m;/;#�j� Dn����~�����"��O]�������̇�+�e�m)O�w��h:m��A�<rA$a�v�� X�͢,>�T^�Vy~W���.8�u���r�$����K����`�%@��e	ur������77�L�kđ���3�����i��$#;��#� n�Ԇ���F��f���M]%]�Yn�9�2=i5+cfM�gB����R���?���QE!�fR̳�p��ʈEuD�������a�i��{�IjF��=��0�u�3N�ZN�;S+�8n� � ���	>�^҂ȦG�h.�[r��`^�ۘ��_��?.���pq�+ |��v(��N�5�r~m�-�s`�H�� ����+!e��6ebǈo��m	8P(��4��D4�!=GO%��� ������)���iG������%��6���!K�t�����#/��%D�G�	�\)�
W�ɺ/�v�
ϕ�U���W�&�\�Kǯ���߂�I�I��ĉ��x��,��q���WX�tڬ
D���z���7!P���2���G '�G����[-|{�(<j��>'~��Y�HjDM�=էL���@��E$-٨���3���~'����v�L(fx��>�]ꂜ0��z~��{H�6J������E�~+1Vh&���)
$a��t6`2�����Ai@�Z^5{�{Gr�s�]�_~+3osYeo�ޅ�N����(~Y�X���g��QO(MT�$�m �t��ʱ�����_�~jE�FT��w8��e}'�}�n2kv|�dª�3�(��1A�Fd��Yӟ��#�����Q��33'{Z�s�\��X���wl�M�3(�F�B`�����i�W�Ee�yO:��ϴ���)��E-�*w�,hHs�Z}���O�22��w��ה��ད�4�.|f�l愨�p�f@�\7����+�ת�����G�J'4�W�!2N7�4����&ՎX<�@�*��/#j&��`�:�0��V7i��I�X �L��!O;��M�u}%�J|k�F��Ҟ0Y���c��w��K\L���lq��� �/��΂J���|Y����4�)V�������|5q�� +,;��6wO�؅��/c�����#���.fC$i�zC޶��MȨ��\���H�܅�C� ��#,���C�t:�<�&D�P�*��'{>���mdo</o)fP�574R�v�Z�C]���/��TM(�d�<�k�2�3b� �X6_����1�U�eY\pM`��B�#eF p�;'W�@�+2s�%�敿��A[A��P!;<�/x�L�-Mg���xZ߆� 쳆�'LA����sJl��v���-��(�21H.��|\�8���b�)[��9h��x>��D�Vr�A�)��ɇ����_n�bEB���.xDA�rp�Г�O�Ҝ�7εz�(�q���!z�eb�������!z�|�h��cU4�&���P�`�@��d�`�w�&��{�N�d��Ѹ�P�:����*����vg{T��_��

3l�|�>΢u�[]���V�&q��� �ڹ�U_Op�oZ1}ĝ��d >�F��Θ�<�F>E���)��2'	��s��	�,�"<wdj}[��z�h�#_��#���wS�*��M}܊������.��r�b���f���-JntT%e�u��ݻM�3����oPd�bL�FX@6�T��"�B�g������V�Ng%�&�bQd��j�>����:X�ALSw���:O@C`(�l,�@3�>�Ժ���3n��N�p��]�Ik��W�W#t|(�>?ܻ�s��]?2p�#����z�K���pb&f]s�Ƨ`�I.0�H�u�������'ߍ�)�,8_���O[�_�*Y��fy-i�� uE0= ��W��}��Ʊз8�۲�9��"�z�w�|��':��R��ߑjww�E:����|?�e�n~�ǉ�51��� Ь4:��n�������T�����^��fr0+� )'����R�P�#`�6�w�z(FH���&��fc�[ب\[��������h
�%��i�����{�er��3�<*'n�s�ꙅ��F%�$��:�Cq��2>�4"����
�����T�وy�U\Ժ6��,*%խP{�:����/Ҍs��6�?r��]p~�n�/Ԩ�$��de). $�8�����a������o�*�뒅3�:�#�̸��v�u!�G}�:��RT4ҫ��[��2�1;w}Z�[��_���m��5*�1�t�:����%��}�3ɹn�Tگd��J�ڪ��	a�o³� ���Z�9
��[i�'�W(o�1�|�!�7o�Z��x�q�2���L�Զ?���������N����L��bzꌸ�W?F�h�j���O�A��h���UDxO��G:��~b���<Y���C�`c�ɷ��,
���gMq z���VT��1������S�^j.v�v�C*\2VP�A�Ez��툧ׂjh~�*U��ؤ��=�-�rS?�Zw�v+3ͷO�I��(IF��D�uT�]��+��9����~$�9�R**�$�H��A�X��HԵ.,4��k�_{���"В��_���v�2������X}T���mPǑ*b�J\���;[;�iMe	�B&�x9���kIi�-�`:�I�c��/|������>y~&�(�eAv�7U�[��2u>�F^a����~�ˬ=��C�xW�,�i�B�����c�38��c�[+^r%��]m��ߠ��٨r��COwi����@ɪssvO_ l��K�&c�N�ߴ�J���ߍF)�����!k�0&��x��/Y0x5���$�į5�>vL�5��N�
�=�[���}��ݒ�(�O��ힴ����>��R�u\��|tB�ʨ&ո�?��S��I0)ɊbO?Р���d���I��R�F~�@���M�G)�~��&��'���cz;�R�C�� h�x�έ��žXL��*z�ԭ���-�b�"�����Kp��E��=3��!)k�[vUO!���=�!��Pyq,A��LA0j�H5��>n0����H �7�ah4.�[��i�KY��q�����:/sy��L�B�����W�p75)vKi{�Yg���*���n���&�Ě�����>8Ĝ"[���KAk���+(����^��@�W��W]�ќ����Ԛ`�
��^k���˗�
n�W7O���o��Z֙��̈́�A�}"AD��ݴ~̼)�$����T�f\zBO��i��P��~K���A���:"[͡�����Ri(���b�-��{,Z��W�x3��D�#���(� ���K<5�O�Om1�M8�)��l!�e���#(����F���l>��-{xO���!Ns���NA�pYh�>*uWO����.��=����&3��`>R�؊��-�H���Wd���n����F�g�@��'W<6�������e�L��f��* ܾ���y�Pg��R���=ӽ�t��B�造�|�����բG�KVn�y݉#|8Z��JO��J�P���Y|#�ܗ�����@�qC�rd�t����ƢI�y"�!��QTP������-��u�� �8��KO�S��^��R^Ks�A�͜ņ�1	A�b��w+ DG�|	WWbP���$B�{#�ي��+���L}�ORÁ�2��J[��J����'�����'VVj�q�����Ls�lG(ss��fzpݻXc�E;��vA@��w�����U��
"�(9\Mi���/DZmk�GT��n��@Q([d��2�����i�����D$�Y��\�aC�:��zݑ�h��WEl�1�kz��[�s��(��r_��	Y� u?$����Q���@�`���b3MH
O{��t�v%6R��r��`�H�<W3�T6�eD�e`p�[pV�Q�&��K��K2�N��7d��E���""	��`��w;���vK�+?�Y�t���Q)�|Ԧ%�>��UrN���
b.A���\���ψ-�<���?��6\�y�ҭ��5i�x�����D��"�b�VAt�E���@����N>(��S���4.�uWafl�Pã��"�غ�h�V���a�l�/A�:�m��i~j��!��t`T�RN�Z���[�A8����*��U�s*_W:mv.+FH����F����n�*�~�Ӗ@G�Q���k���5sP�Z髾(hoD��e��X��Tϩ�Td����)L��j�w�9�e�[�ƣ�9��(nJ���G͆}Z���Ϯ��@�=Y7]��ݡ��1*5���$�Y2'������$\ԡ뱅ͷ�F�Zq=���Rq�g�L:'�!GS@�qF�g`�L�c���a��>��js�	X*���� `�w�3�-q*�hK����?%�#oBU��3��H �b����(�g�ֹg� <�
�mB�"nh=�����2Ϣ�XC0��Hv��w�"�)�B�����nӖt���4��#��Z�=�t������m����5���z�D��������R���C����
��! E�5���h��Yh_��-�j�;�:�Xɫ�����$�0\i&�A%�*�"&߶�����*�����{&^]T=Ћw9����'�W��
��|�6hq�VZ���K�`�T笺z>��۫�;-�]/�c�C�z�uN���U�~}���m�Y���+�6J���.�I�?�\i��s����ɘ̣�Z���eu���Ik��Y�_�J�q�c{g/��,�3��*컥76�*��&U8��aB� �ѱ�R��n�7z�z<�Y���Ȧ���u��e:
=0���h�����SA��4�gFt�@�d��H	��ho�'����=$�'Ry;Ӑ��>AH��2�P-*m�[����_�����վ�@�U��3�f�&vMԖ��9`iW~�j��?椌�Z��1U,B1 ;^Y69FB9���q�}{\���m�^� �y�>�-N"��+F�}L�h0ѯg@�'q]���;��#k�_~���E� ^��C[��|�r"نe�g�'#H�?��s͛��!j���@~����v��C1�S
�+HYу�D��Ν����L��Ǳ�P2$@YąvJ��o��2`�}�K'�[He���2G�Qi�s3��U��7'{$�}߮D���-i)�������k��L�h>���ص�ί�ֵ�c1s�_�ҢN�^��Pf��4]�%8����_.G�$�Q���@rNΗq`�ҟU*˪˞�w��$��ɘ�kH�f�9`�s��8��,מ�����Μ����c�����TxV D�R�<	>�sz��z�)A��p��b~K�����	����o���������Ĺ����lW��hH���$1�g!��{X�Q��1�W,�c?Ψ׎Ȃ����.�-�V� (�!f�X��oI
*��(�y�gZX�6��i�/J�|Q�Gf �>���P�.���ZZA%>�s��y�`;M-)	qi�|x�����0�ߚ�O2�
)��ir0G��t�˓�٤t9:DVČ?���s�ze��3�'�z��:��6�@��,��R��8�8H �8���=a��^>�-B.#dv�����WA��9��sϪ��gzN��E��୭>����M7�@ $��I�>��QQ*�������-R7����i�E��m���}N{��.Jf�m�fh�bJ���W^���H��y��O�>��(7`捈n�aI�B�>X��I��cѺ$�J����� ��{S�Y����9ˢ�h��l���9"��si\�Q>���6�}ha~���}h�0%S�x��L������b9��o/MW=��O���z�ś�S�h��/�+EO��o����F����~եӂ�� ��*<���N��q!=��dp�Pc���-���g����;�6XM+�)̕]RŸcgl�:ǵߥ��F�O�+���� )�~����kE�#�������ї�cl��Ze]��V��rǹ�q'�E�!���p�vR�5�n�o��m��X��������^����u��S/�p�~���T}J��$�dO���$���'�E����>W�>��+,15&�Pz6�N��  qz?������H�(�WR,��Q=Ar�ݠ>����ԅx���nY�l��;���H��k��� ���=3Sp'�{a_e��+�h�k��>m��vĪ}Ҳ?Z�6'~���F���aێ�$(g�8������~����]��6����t���4]
�(`l���)4�V���M�;�CHrD�(�36V8��ݯ�p�W�����GGYe�F)��_�q����j��Y3D�rTo-�$m[D�<�:�(4Mܖ�̃Q8Z
Y�v��������\��vDOW捕�E��~�[��X@"G�H�^Ǭ�"�&0u�_�
k����_��a�/Y���LB>�=��;�&��Ǎ0���~��Oj*KPZ,<ފ�n���LLf�	���n�����\���H�(&�ۧ���#���<{�����r�ɽ� �5S���4~*�����،�߇�sb����f�v@\9�u�K1�X[�Q����������Ć&\��H���m4�rv�)�����H��!�G
oM�z��_�����+Z>���Fwt�J���f��܎n���'��}���W=d�oI���Ev�I��P ���-������(c���d�%�f��l5�=�%��|<�,H���m`�d'1	[��㐀٨6�yu܈�K�ȾI���;�^mx�c���3֛�ehE&�A���J
���K�nq[6�i�(:���� #�j�t	}
f�s�B �>�#�}��4�.,���ucb�_\��O�2U&�g��k�dlއ���	4�a����5�}�:l�Z/�EA���-D4�n��D�/�:e�J�!�A�Z�n����?��A��c�Kcx�D�<��1KxX��6�ބw�ժ�&:t4#}�\�*�"����/�:[@)L�Z1��uG�`�η�B�)��ds��xr��J�@=��/
O6Nˌ|�Uň���:���, L4�K����g|� �s҈y�3�D��l���줂��o�#�ts�Dje���yş�nժys����[-�r��mq8l>-5�����/�kYI��6NKB���[�.��-~�D��o�(þ%<��[M� �o��15��ܭE�%�-[����$�[���H�V��S���8�. ��j.'K�I/�0N����su�3�Ն�K��ax��(}{�����"�nVW�zM
4q��I�Q=4���mfg~F8kn�� �mgH�WWY�!qa}cY,ay�	�w���J�>5ٟ��&!�_�a��6���4�튞L�m�˹ѣ��O�Om$U�5��y?�����Hʓ�u�(�vw��eS�v�va���p�zg&�-��RSI�"�g� ��Ja9�w�!����jA�kDf��i���[�D�ĕ~��֜c����L��񾽊2�J~��0P��A�2Y�Oш ��Zfhi\�'Q�[��F��X�E�jll�	q ��f��_T5d{\�����qR���.�~X�� x]�e����H+���:'�����\�?��y8�����0"�+܃���ڮ��i�3�cnj9�VN3�9���F� �wۻz��B����V��k�&UU��@:� cy@^/#�A�j�N���ޓt��k�1�w١ܩ�.s�?���Wnږ�D��L�U�OU��i�΀�f�b.�ϔ����Z{۝ϫ�����ɂ����/�J��1���ib@��
�7��
f58�$�bX����ʱ��Z��	\r��O���땳!>Uܔ�W�$�E��M�ِ&�A�ra+���mU��|��G��@���zS�������m�H�g��dg����~�b�����ۚ�X6Tɩ�"�]���9z��p��y�6R��[q�u�Ԁ�`W��60y���l'��hQ�	Y��>���ȧIݿu�D�)K~R��^��(�luO�\���
\?��~yV1R}?VT�2����� ��ʁ
X�)a΅\��՜\�B'�S�K���~IWuC�w��$<j:ap�*�Ꙉ1 �x�N"ۻh'nG{�|-��!��&�q8�*���NUل W��:�:-�W��W�(L@H���������_�H�'r�?�7[�������\���Į�Q���}O�BA�+0�C8��*�$��6���i���~�~i�6!�Rx��Nq�h��K���� O\L�D���̐II=?6�5����mmd�沦Lz���B��E�	�)#l�T�y<M�ƁG�R  �@�Ѓ�r�
����~���-�����P̯��r��/�ԙV:HhW��o�n�SVnV�c�'d&#���롰���d��[��<���gwN���mU��]��Tx��<%�
8��*6� I��O�?tě�W>�(�>w�flxh{�����d��$��g�˄t�_H򕽞��E$�+��3^756soan��uI��˚����d����{�VN47KM�U�LW���>�=�q��Ƹ��;F�OO��9�{I?���lm��2�}���C��̼���z/T_�.�珩kKn���n8ĦQJ#N�<�h�y>V1y���=!��J ��[�ټ��)����\�݄ޜ;�C��#���-ӕ+���k�<�ǽ��5�ϦI���H��3�s�_yL?�+���*d�����D��R�*{J����ƶRf����u���Pm'4�!��B{%,�{�p�$��^'!o~R��W�m�X{��c�/���PZ\������7���	���r��8!���݈R�������6�>q5�g�U4�v-̛�e��^_�	H[A��=��G�ʳ��̓�-�z�V�c�Q5���&�v<e�Ѡn������I�f�=���6��F e�D��^�Mἔ��W�7�}8.\g/�a5b� ��z|�IK��3z;�'��i����.�@�A�M+�@@��w�l��i��B�G��§��0\��~��7���lx�5�®�a����J�A�}w�"���^�M��'�������L�HV�U@x��V ��|�2aŎ��p�U�x�\��xS�ᭋQ� ��r%�(Q!rnJ<�)��4�Y�1��M�-��DdqC�3���a�]�������8,���huP2������co�fS�ID$m�[?,�@:F�Y$?�V�n�Q������P�b�濇��xq��/[t����&��C��G� 5W<Sƈ�Y)�Æ R�l?��blc}]�'�ds�����ͣ�/D�/~�&�J���y>�G"���Ϡ��Ʋ�խ����q��3�۔3���Q�0d�r�Q�5x��w��-�7F�]��C46��g�6���4fo���J9���6����#(\����ojmS�b���U���|PC
� Fׄ���C�Φ}Qx ���Fr��`�I�#�i�h/�Uy�_�$�F庖��}ƽ�d��iR2�ў*8�|m���ʕ��#aʢn�}t0��S=�k���/�����5P�G��X�څ�>9X�"��}6&�,�<%�U�"������E�f�B��
ə5�RM�W��v4�h��55wE��m�xz;գ�)'N���`�z$ኊp��~N��F;Ќg��0���n2����A�W喋�G?��9�űl�	��C)�H7^8�]hR:�؊��v��3a���������rG�x�|+��vseCe��#UZ�g��H�q��Q��7���_J'�\-U�,�-����ơ��39�����J\!-F�$�t�`|����tA�n��"r)ZtJ$���G�ZƎ��2PF�I�Nv��b<�R�.��V��Dh��Xn��|��_Ѕ{"9~�`�Ca9��#8���a��-�Cu4)�nI�4�X���X����>?�M�(u���P�	ϮBL��>1��䢺!��F��k�k�����ʣ��3���PȻ=��F�#���9o ����E �Q�0���&�*��q��ǒ L:��ۉ��px���+;�:Ud�UU�ꌈ�=+��^���q��E�1tX��v�:|���<5�V?+Z�R���f�Sb�]m�e���}.�y�1�3��0��f�~4�i�;�3�gF�r�|�/xpV�y���+�
��j&+�����(b�м�����ű��h�qn�.�5�ęj�7�(Ja���ͺV˵ZaYF.�(:�E㮁�G��B�e�����w�@�����yNq��t�ƙZ��}�>�mb��ν�z_b$��l��u��]	�e+����j�UV�s��F6s/�
s�ՁwB�w�}����E o�>Z�^���x�K���%-0��Ow�ui�&p!���t��'P��']:(���x�!3�+'9�Cɗ^��E��pR�Z��8 3f��tk�fSD>q1����h���Ġ��|���jպT3듇K��" #������W�T�˴���cX�����K����`[��)��p߃Am�4O܂�BǼYPT&����ǲ���%T���|��!*�BG�U��F���'���[�jUL��:���	�DI������([�wr�
>�f�aZ<EK���4�KT�_Q�TDҐ�׀	r���^�����@z �GRT�eQ�f��f��M<�Ʋ�@���A�忂��s� �&���B3��;�k��yA�4�CM���p�8�Ŏ����+5�{�0�t������z�(-�6�-~y+96�tK��_H��}��tY�ټ�CvZ>��2��S��ƃ���T�i5�
�ؘ���A�:�>��Ʋ��e��3�Ʀ��|�S�P0��\��Si�j��bJ�&�_z�t�����)���K�_�\�{�0ڟ��n���æ��<ʹprc��h�9<w���By��tj�0���x�Q�r��7�9�S����aO��SOBYA>Τ��ZV.� g����&�����]'N���'��Kbzfe'�*�����<�A�:5��2��c[����׻�Z��$�Gc�cW�<����O>�b���TƧ��`�A_t�;պa{�pj1V��&�nZ��m�:��{`��
=֧�ڟ���w�����fwyip�I��B�䔃ZPv&]�&��\U��R>u�M��!��9�2�|���9W^�$����s}	ez����2��_D���kN\�(t���{y�/�:F[�w���җ��@������`�+kܺ�G�5̤�8�hr��1ݥ�?��0��s�m��PN@�k�@�.&V=�"��j����,�DԔjN�4՛l�c��PS��	�� m*������V�������Q9��37E�t;���2��Bi��X�� +�D�Q�|�g��,���"�`# v����:�e�s��'
����� �d�
ǎ́���1]������D�)�IӒ�{!�&����;�Ѥz��s7�6P|�wh���|��t
>�i	I�tz�u����`���]_�)�����v�=<���>��C�YǶ+�@��uvy�a��@��-�l��g���7q��+���w�G���,19,Zk�5�MR5��i�B���_���(���0%���Q��6����*x�dcada��q�F,��}���9,���H�?�����DE�������O���3ךx7���O%*phe��re��uZZ�Aq>�\c��	��!���3t�Cޖ���kՋ���5@�Hk�D9G!~=\��!�6_+�� �����D ���ʓQt�2�>�F-d�o�:0�?-�55�kj��P�M�09��S|��� �T�*[!D�|
|�-�h�
V�Q}qB�]�����=u��.U�S�/���Y��D�Js���m�b/1���#��1�����<c��Ƌ6)���Px�A�Дmn����B�W�����0ЦK�P�
��w��=y��Q��Aj�U�4���č��ɭk0��8��G�7�V27k �������
�߻d�2�\��|�dd������.�~��2���"�Fn�\��k��w;�/��>}��#���S�+-zG�$�huhOe��<dUhUD5%c/B1��.sJ�0���?J���q~�>�b�w�!|�S=�s��Z�ë��|$3(����Ӿ�r���jt�Y��跷t����ޜ���s�]@,i,1�t(|�F�4\����Z{�%'�;�;;��O��iO��j��CX��{*��o0Vר����,����WHT�E"@�*%/���9�v�!] ǵgj��B���
y�b��W�����`��?��h3R���[�9�I[�[T_�T�m^"�U"��,閯Td{�n��)���g�u�A[D��s�<vg��8�����e�Y� �'�G�.xǰ h�~��R ���o�k3�ǥ�b�^,8̯�H��c�����v�t:Ip&�xa�=�g��*%�f��>�E���Ej2�d3^8c�έgзE��e������~����;�h�{�ɱNx��-�4�^�֤��)+\V�$�
�gA�M
��L��fn@	��+���ڑ)�!���XQ��b��7����w
��F�_���r/�b}�����Dp�/��˔��x���p�|��O��K?�E3�Zş�q `v�u�b����X=Ǖe���Z���xL8��^	 l)+�����*��F������]cl�/ˢʔwo��檟iFV-e��\09��hwhAf�P\f"���(��:�&�~,�֦y�&�>�2<,�w%��������&�u�:|V�AMQr�$5^��"�/$3uĽ_�� M�5��ˁ�D8�5jzB�3�h��n�.IbH!��sC��}�� >�ƪ�\&("۝nRD�sKS�8v!=G�Β)�L������{�A��ψ���6j�q�lx<�P^�#�_���;���\CZ�c?K��\g�B嬇=M������t�?�
��2qѵ%R�K�2axqkp	:�qN�r4�v��@ 7���`���|�W���8CO���v�~�T�|�zݘ���R��%�ܨ�W���0*aE�)��r�t/l�R��sq^�=W�Ҍ�:XSnˤ��ށ|sm��aҔ��nr@hkk;)����vpǊ�d��)�����[𦟛L'v�������X�,�j5o��L�
�g��in��?��m�	�I�s���+��8p�KU��@(�0�,%�a1�=v�>��qD!�hD5-����m�3^��͚�ǎ ��8�</��s;]���[���m����9AX��9���¡����m���1�����C��W� ���)y�?9�d�. �3�@I[�q0�B(����&i�΃3KK���S#�u%�Av-�ņb�q��=9�hʌ�̊�1F�-kCT��}���8f9�s%�9|bU+O��4�����4�Er���X��$d��䤸�����K�'��Oړ�{�v'RY]��["���'���*mVd��t���Ӟ�bb0S v�y�VW�7�.ΎQQEI˺��|X�$]�ʒ�����E��z�R/!Y��glt�+���<�k��.����Q/8j���S�9{~8!Y0)���/\$�]݆$�fD��Q!T�~����G��_�C��<cx�6^0����N�Ik�
�9�ϼ��1k�$Y�Jl�qQc�8�Lm�W�����o�X|`6;{�1*�|ܠ7�����FP<��O��CP�c�}֥Hw��y-rߓ[��xl�'�[����gZ���_� �VJ�81_���j�_�� ��OD�̸E�����]�|�0l皹^Z�,�_ܾ)U$7�,���f�k�Jr3�3�X��d0`�炈� >����)Av)5��p�C�y�ѧ��Hz���� �}�)
y�5���QyOֺ|��+CN�S&��H06�s�Ʈ���ڑ�� _uX�'\��+�v�KЕ��,J<%>k-^ql;*����>2ŹcK"ߚ5]��X��I	%�gJ���ͬ�f��F_�r��+�Gx�z�W���@��:�տ:1w�`��MK �w��v���;D��^�2࿞G)aZP="�+&�x��A��HL#=���A��)�,�-ڬu�(�s�B]��×�WT�P=���Avov��zf[9��?���(�OX�N�>G�lv��m��|�#�U�;5v�@ԡ	�`UJX[	��������eT��Hl�+��+M���>3���R��%]̏�}�~=ɡx�(qzhv�hkw��zQG= �fg��ߋb�n-�˥�����A4̆���j��L�'�$�w�
�g�c_��K#�7�|���*3�lx��������F��J�x�.&�����L��a�ck��̹��Q�?��̔G����1}t
@�*��L�0���Zo�J߁tQ1����C����a�>��nl��ب�\�sJ-�~֊��
��cʧ�"S^9&W�s��Gd4lr����W��>@#�k� Ʊk^��. ^E�rؤ4j#�cU��ʀ��t��z�����^�8�SCM�
֕�2#��\����cLӐ�D���xV�u����� �����,��GH�9��`�`�M�v �t�T^~><��x�ԑ"�if lR�F6�P��Dx��)��PY�_�H5�vBZ�I���Q�:g5v���E��NO�=��yf8�8f�^F�&�1�������;�sm����c��mY�]MXq�]^c{����c}��LcMդ�b��=�W�Nn��D�.F �NJl�3ߖs�}���E��E������nPO�x2e��$͡HT#�5%��J�S}m�=Y�(����Ȓ�1���A�ws����c���p�c<ҵAQ��;�*L���w��I����x�d �j��Yd�VL���u��*�	$����Ҧ#�o�6j"�S*�$j�G���T�!�����l�CW`#��0(�1�r�<�7��,Έѯn�;��[����N�;�ބ�V쾲pH�[H�g�M�F��l`o	?l2�V�����5
u���j*����
��J_�����m�Y�1y�X[��O+�&�
ߍ7����q͖k���"t(���<z�_})jo�l�^���~\� ��KP)�柤T>!���	��I�����K�Q�315�1�51��CQ�'7p^��u_��9�J-)e�HM�D�OgE�5�U�G>�'_���J����{Ӿpv6�KY����#��X�}� �Q��kh�	�g�0�,���X-�P_1R�F�]��{R6F��zy�f��C�W��Եzx${Z���t�CN�E����b�E<��%B�Mm'ﺆ���R�3�kT+Yʼ.���{� ᤄ4���~ai�Yz+�U�j�'ûj[	��~]�|�C�<�4�AW�/�4t"�RZ��8��r^A^��x��i�5����rj\�*ƶ�/�@3Ð��.T����8<�����E�_����PXk<������b���B�B=�zÄi�~ vs}�Q��E�����iW��^㇉
<g�Y[���Ueup�bUU"sʟX�(�N�eS!P�s�0G0*[��3�vwg�~�a��:�U���"��Q
���Ӊ�1JC���0���y����a�Q���t�% ���� d�hu�
u����4V�P?)Z�Z?(1d-�}a|��P
h6`�6�B�wHLe��Q�H��*�E�.���֪ٛF\^�
l�%F����!�t�_{�d�g��r�O��H0�x'�Hts" �X�`�K�35쵽i�&�q�~`����4�?�lr��!e�k�M�cP�+"��k>�j��@����*��M��~ى!�ʔ7`��n�⍮���AM��+�z��%8�=�hKdb1
6:��Igу.߁u��b�W��'-��W��,֘v?Z�+��C�����')����V�lD�߶Ѿ\|�?s'-<l��i=u��FI��qQ�镼j�`݇,b
�XC��ykv�l�+�\�����)Q��97��n�G�%�ؘ�vS`�����.�l����.2�f�\��N
�lA�f�i��蛖a����{��Nlk�O��θ� ��E��������p��ٿ�B�
� ��]!�6T����ŀgw��W���7���Ć%� ��	�ebE�M�36%��$���^���Q���m/b23�Ӛ�W���4o�*�u�ll��}��=J�|i{�.4wƆz�s6��cpc��nB��q�[mkSdr%��>2���g��͑Ap�J�̀!�2,��Pk�"�&Cc�4Z�+a����	�l�'wnn�򞷤Q��K��A��݇�ҋ���d4��}�['[�����R\c>7C?��q$$�_k�~W~5�*��4Ҁ���H'�G�
%��F��������M:x����l'i���|d���9a*�v;�fn$��A�5;Z�A� �I�,�u�xp�yz����$Ic�G�8��><��V�.��ꕄ� ���'�L	0�q��1�ݚ�)����*�5���%wuS�����:nR+�Fi������2R/�ḇ�ȴS�]�tS�}���y�X�gի���j�mԴ��1��9�5����N�cߊ���z�I�l� �����F��tA�ol*F(I�B;����&�R�w��0�U�>¨͋���}�㞮����n~�M�~���T��~G�g!�K�V�c�D{�E�6*�f>�@���rA�%W�����_'����}��K� �uh�y�m���0�,��[��T�s�G̟)2��7��$wSA�T�P�a&hQ��s�>���3�(���'�v>#�4r4S�������p$@y�5���n�_�{	Fy�St�\;q��Z���Jھ��K�.��"B������<ߵ���{EK��Q_`xJ��4�k v�o�h��$�� ��"�l�����)I�8��r	�Z��t���>�Ϯ���$�F2��4��+�ÿ����c�^l�{���lc����cd�^��AO�����̊�xNq�~��[�ܐ��[�����S��Ḷ��H)y�O�8�N[.�w��i�9Q�'9�����)_|$�(�FgRc2�6{Ee�_����;�>��Z��UY�ѽގ�L���O�^O�f���2S�<]SކpD�	,��L�����׾SWH��e;��%���(�W�im��f�����	����Y���ɽ���ap��S��ɢ��?��ɰ!=��n�HP�m�P��;}GʬXU!�9�uS�E�����)��=K�9��f�HEC�5�r�W���^g�Pm�Z�K��4���W�/�t���ғ�62;��h!rkt�E�8�c�bv�M �yƗq��j���Fe�
r]9��-���_��]��t��A����;]8��C��c�Q=@��Ԓ�1h��$(��cm9E0�q�n!��H���#�%�c"���{d�Z��o����kV@�t����&l����B��h�!����ȃ�>ێ-b(DvSe�BF��ؑ����_�b�P�����v{�]��j����L5��z~Θl�I�K�����v��;�QH|qa��i�r��IdFPW|U�Q��X{�z��1�������/nնC]ke*-�;�J��G;1�q�Ŏ���Lm�.�Req������L�<�@�;:��`ƁX��N��Tɫd5�J{>Q�?����S )�/��Bl�@���K�̠e��-�oM��ɵtr�;^`k �<�=OH�$kTg��W��$~l����pV�q&��zmo-�A����f�9r�5c@�<��8=v����tz8��}P-t񚸀!i]���f-�Act�Ƭ�z�L�| MN��]�dg�7�qSGk*Ph��_��\-((�0J<�����  Z�D���h��K�����~F}oZ�Dt�w�g�Ȏ"�WK?�&�@! 7�)?ͅ�����0Q�%u�QCz��N��M|f�b?r?"�F}4J��Fz[P�Nk��<���f�8?�=\,.T_Q�ĺ8z�f�(�gaTi�)����t]?V�`i�daֆ�׉X?�������W}�s��Q%�H;���N�{Mx�.�0q �B�.�ג�1�ʱ؛������iL�e�;�ͬ�v�b�����b� l�Q�X��R��þۚ�dUI���oXf\}Ϸ���k�ʹ��Ѫmd�B49��a%������4��O�HBH$mKP�x/��j�*p�j�7_��$ww\;ϱX[��iPQ�(������/$�,ڍ�cU�k:�H؜E�L�7�[(j�R�8R�1%[A�#�������3��M�����G�{�,u^�D�$c�k�QӪ���y�~Z��.+Hܲ�0Ŵi�)iw�y6iytbݠ�ki?Vs"��~٥�v�8�Z�hӉ����%�����QǑ&{�WϷ����Ś/V�����T����խ�E�.�8�� o��w�c�A�l6��,�g�D����O�V�`ªHN�������]���"'��t�^�L��d�x���Jwt?�
!ɳOLe
�*�H7��랷b��Ə��1�4���Kv�oh_�p��T?����jG���j����=g̫���q��u�Py�!�{-�[M�kG4%1����5]����y��'�w�EԯJ��P���3w/���B(�PM �ebCH����Υ"R��
.�y,g��
*�QW1�M�[�.ۣǬ��`W��V
2Y��O!����\�G��F��+���J����k���D�.i���Z���$Z�|������Nru�y2��n���UYkI�t'|�����4�'h���\8�'֢U0>.v:���?d5k'�h-��o��R݋"�:��{Ջ]�����T9+���H���N�i�w���J&���s������˻�S�pwY��i�&{+�[�I�B��No?2��Mt��3�i��7�Ll�@ɳB�M ?�q�0n���hs�h���!β�����~I���&�=�J%х	�/*���6�%��Q�^���J:A4������lo��k������(�5�0�u�48o�Z�3��]th����O���o��,*���m�qK��Fj}� �+��-Il�:� 韗ɬ!5�ƚ���ֺ���q"�I�i$,R/�ܦ���w��/��Hf􊽆sK�Q,#��qfu�!�S���I��(X﫱���k�A�����g���T ��n=boD`@bˬ]L�!z��ȶ_Pa�����q+�y\�Sqp�3� 4��v��X
Tk� �)�In?�V�kP��ib��_.�oN-T6�^���w�[�F�!�]�z��מߑ�4Ђ"3r(���*>�&@��h��$�ʽ9fF+���ǖ�YHM͗�｣�D���E�0�)��U��u�O�v��Z��6���#D}��RE�ˬU�+r��s�w��D�]5�ǔVH���p��P�!JJۡ���oݭ���C��1}ͨ�&j��aq�n�����H���]����W>g"���vf��
�eT$�v���34���aY�����D�p��ᰭY�a�� ]���N8��:��A���=Y��i�L,��a�S�π�4.� �7
_��X��_�5�����`�݃��g�_o��8�-���'����.�䈴(��_X�P��wL�eʃ���wz3�~=W7���Pp�L@��<��=t����dS�^����#
�k��z{�=����|L�&����kl��E�qLm��1GL�w�6&t����d��r�MU��?�e�{v� 	>}z!��J)L�o���2*mU�i0���Ѽ�@�H���hF�¨������LZeڸ8:5�O�"Ŋ�聯�!�4 ԏI�\*ZX�����\m<�I�s m)h��ů����Fx�D%B���?b��� Ѷ?&/��@�u�-	@H�!h�@�b��?a�
��uڣn�+�E�{�Y�۪�(U^����(5^����	�"'��|ُ���eWa��tT}~���M~t����F{f�T<^P�{��M��$����!)x{E�cAC�ۯMo�D�7��R�e�gl��Q-�9���hC��?�k _>9��[��>�g�Т!�*p�������^��Z_5��A��":q�܄|C��q5zm/�gHv%����R�lnvaH��ع�F��ߐB��,B����cߟ�u�~x=f#e�ܷΨJH\�x�p����N�,����Ve4NY����5���?�:	vT!ų��L����C���D��u^�&9��L���>�[����(��RԱ3�'�F�>��V4�8�9I͂�l��g��v��H\B�Bu�9�!�?�Әi)bF��+-� ��^�Ǹ�a�ڬ����u��/��PQ� (ϊ�=��t6�������c�NU���H�����-�KBY	��0�8��X�D+�G�;C�������%�' �>�6�}g#��Y��NA�Ps1�K���<�����YibK�;�5��m��~��)Y�[R�֎^A)�76(	�ٟ���Ddp�v��S�C�;,��PD�.�or�<%�Z+!$��~}�C�([�
��9�
ֹ͠��焲���|o3*]�zOMO� ��Ⱦ���B/TnV��H>��U�uB/�J����N
�K�"`�1�f�<Ǘp�P����BL�XE�u�t����O�b�*9���		��{�OF�������0�Ju	x��W�nWIO�0��z��������͌4	`��H3
�#�� yu���0P
� �ø��`�h"i{������떯�=�F%$�O�I@��処��kp-kA���?�i��%&�{�ޅb�.�IVm���-y
�-����G���Ur�w:�A��,��u����L%��·�t&���&��C���3��}�� �0/{/�G)��RCg�g�d�l��J��I���I�
Jo�~���;$%�3��A�����U6�XÆ,Tx���>�,ݖ2�^������I�� |e��訥�=fFO�fW<Ś�铉g�����h�~ج�r��8VJF���0% �_��+�ޱ&�C@���K��j���e��е��T�� <�~�o�x�H�W.-]K7������7)B�HƬ^���ޟ%	�5�ķ$e�De0М �K:�ӥ�6�Ⳟ?Z���
��7f7슰��L�M�Jc0�T�� Cu��� ���OWV��j܎���l��c꺠!�L K�n#�����D�^o���g�����v�R��?0"���<H��tX�G�ܲ\�
d�N�T���|
�!zF�� �r�<3,���[\ǷZ�Ǒ���8q)6|� [D��`0S?y%0Sd�b���vM��Q��{�3�u0�Pt��r�x	���&[j���쑑�B�D$�'�썯��촫ܾ��@��̀�B�t�%=miH{r�6�K�R��;���f���� ��h�(�Y��6'�"�Fy�IL��e��n�\�~'3����x��"�~Y�l(�hͨH�&@�2T*����y{�H�Q$��W�,$��d�J��H��}��ⶵW����$Ɏ���,ʁL��a��}���%�&�������j�hHzˢ�9[��tv��q������HS=%b��A�O'�g�1}U��h�	܏���FmK���X[�߁N��p�����^���Ɏ�+��D���3�G����d8|������,�͞M�j�0g��`�*�sNnvWU���P:7ˊs����-�O����{�B�G��-ŝ֓i�V�Y�˭�W�%��<Fk�[��;,��g�?��#w���j)�U� D5�dL��D�V8� ���Լ�~��Wꭃ5t�����i���&hk�^��+��n�<m�_E�:$�a�07�Ss���f�8���/Z�B�������ש����|_��k���T.����.2=�H*'���)�o�l��@���
`��lM~p�R""��
b�����2�Xs0"�3�T�E���S��wX -9Q�nr�8y5��솱Yd]o�oI7L��,w�@c�	�������vnCn|۾��(W�r�	}fgLo*
�ꃾ}�	MF%��U�������s���r�Y�j�塪^��mI��E��
/�j#�A�8����.&T�
���&���,W���1���N,�.5�KI� Y��]�6 we�<����H
*I����� )ɞ��ȡ"�H�8��)����#�A��Yz(iχw���^��9c�1h�����S� ,��{6	��{6Q֗8�ә��wX����{cR�r�װ�;@݄�7?�)Hُ�@C���[�^��7Iڀy�
�q�EG�S� �"�"�\b�(���N7{ 	%�����W�0xW�s;�Y��ؾ��@�'�|j�x��&��E(��A;��%�j��9�@����#�En�
9��K��G�`��U0+��3�;�B&�뉷����N+;��G��T/��L�i^Akғ��!�5y��~�@!Ż9��������L;�8������pg����R�c���)�1�V�)�-��W/�!5����8Q���XV��a�mM��aH��d�d�����<pH��?���ʜh	�ç��ck輎e����f>*�s�9�4S8n�s�@)�y7JLL^�~T�<��+���~	'��]D�w�c3i���)0�zD7�.Q����5���IOp�(�z>�)!R������O������ޚ�n����G��i���I���c�$���tM��Z��]�c"���r�����R�QBZ�9[[B�e�yV���ӷ��C������8%��b�|v��+)ԍ����p�����
��_y�@����J۵L���ş��;�Tx�Aj��be�*$%+��Fn��sC���[=6��� �rc͆m	�M@�(��a���=/�ꈠ�����}����u=M!��_\^���n?��D�1IS�?6�E�J�6�Q����4%fA[���(_zFe�d׸��︊��a��i����q�
H��gb�G�M,<�{�ij٦o���� x@F��S��0�g�]hS��C|�n�ZP�̏���3���	�5�8�n��Y3�A�k-�d��^��	���x�=J��d16�����I{�w��k!��W]�~~����}��XTfĢ/�m��Nݵ�>ax�8���&��ʖ]�<����"�>�G7����2U�U+;��`?L�HWљ���a˱7��Jp�u�&�	�
|�-�M3��K?^�z|C����74�]wο4U�&RL:4\�����,�Q
��,Al��l�\'-��P��qm�n)����W蕃n!]�*I�� �ܷm8^,�OC�,c#3n��v�\-�3�01�R\K��4@�RU|�8;r�˰�cRY�h�Y��^-����2����eCa���ݰmF���P��/S��f��t��e�!�eR�?�Z��F$h�5l�ԡY�� �:<{�Ak�ْɕnC�چ�gU�=,ִ�^tqG��s�Q!��ܐS"��60���X���X��c�N�+���p;GQw�q�
�D�|Sڏ��6�e1雏�U�r����;�(�Nd[�z�Qz�?��p�󦭮�t{�����
>ZG��G�]��m�5콲����� �2���rb��Z�9�~�k`_�e��>[���J����]���iF�ve���A���xN�!����8��*�0W<���N�ӕ�N��#!���=�ud�h���Vq�P�p�j"����՗P��SH2RUV�Y���������c	̭�=EՕrq�%����PJn�����m��ߠC#�~��a8���N=~]��',�G�?f�(�jV
��֜*9���-a��E���f���� ִ�ݾ:YrO��!�I��L�%#oTʽŕ���6~���ߚ��f�D�FeKƽ�/ xIF�<�r�[}�V����O*���ѯ��<s9Kk����,.ٛ�h�:�9�H�g�2j�����$�b�N�uy�y"/��!s�N3咶�G.z�b�������뛭ʫ�n��
���"��f�@K
Q{!X�4�O�ƽ'��@ ;VZ��4�3qK�7���&|�$<��ʈ��o҇��n˜�`��F���"L����5n�)����� t��^%���ٴ64$�L�x]f�\6.��;e}V��@���'��h��U����R�Xxȥ��/z�E���9\�V�x"�c1�R�K@�$�{���U4��@%S�{����W�rJ�G����|��i4�? ���Qc�##a��@��OΛ�O�#�R�k {ڜP��6���_��#$�(������Oì0R Yz�i��X���>�Ԥ���p�b�u����*U.��[u���HÔ�Q���$�p���8��xE�A���
M)B�����OR�76%���������q	S����]�E�hpD�!g�<��r��N�{>�=zukn'��s��2"Έ�#)���$E��q�m`vP=ܟ�y@�匟�Ν�%�kd�w��@��8pf3S�v����,%)�0��]�f���=f.��zt^�<�r��v%'G�|W���H�_�++�tp��F������c�CL�i��Z�jz.��s۩Mi7��0�?M둞�Hǃ�� �z�E%��/G��s�\��}ua�B+,��$���;�M*��Ż1��V1Gi2��t�$���4�;�1�5��E  �����kwtߢ(W�կ��[��� ��ʝqY~����*�� 3ay���y^��I�=�ԝ�wy	4�Ҕ��a ���jڜ���Y��Y�@�E�e�dM��d�ǒ�~z�հ �i�n���噞>���������"���^�B<V�v�DWTF��w�y�Ou�e�lF��.F8(��iǗ>w�3׻k؆�O��3���e�%~���z�~��	�|��g��=�G4��d�۠�с�l��O��͡�^���+�������oW�(Wo��b�ઔ;��~���)u;]����r�&�.�G/����c��"cQm�)k�Ћ��B�S�4�zs��������he�݇[�HS�&u���0R����)�i�ot:_��9*M�\�5x��J5l�ڭ�@�=ʬMv�^ȗ �-B���J�E�B�c�>�U6���OW��Ҕy� :\��:��^J�/����d�S����wZ9����H!7�Y_�mU���!�+������l�[hpQ,\��\�\$�8���/��rY�*�j�Ə����CN������",>�	��e��GlgHn
	��jm���t�YN�@]�ݽ��k��S~�C�Z�;�\:ݼ&���5eDeͫ+���]9gzU�A5��xD�Z���,���o�Ax8���/��5#��qQ���S��J�qݖ�ci�x�(a��|#�:�����>j�v���
�I��V�����%��s��k�,�S�uE�q2���
jf�%ZC�ֱT��z~��_��Md�裠㹍�,�Zgu���H.78\�R�����2Sd翹����bRJ�݂��}�f�w�qw��w�ԗ�c�T���̒�C�L��nY�D���Kyd8D7��enaŪ��^�1����s�2�z�o��:���0�i��7�d��PMi���~Dĭ)2���.B���>B�� +���ý8�Z��s���o�,˱O�)�Q�)���IHJ1���f�=G����Gpd`F?Zsk-:���Vӄ-VE]��7��v�ϓ�,�����$žQ,�G]�i�(.,J��*Թ^�45�RA�� Om�fK���/f+�%.ݷTw��m�8z$����۬���4�xјnj� ����qsާ2:�Æ����y���Q
٫E�ּ�5�~��L��\��%��DF�n���Vn
��Oq����m#���[��7��b�R1
W���C�۱��;m�щqx���G��D����a��1頞��W�-d	��]�G!,;g]��:9���"\���p���g�&��J�� ��cA��s�e��}麹k�i�$5�G����^��؍�s ��b<�ݰJ��f���*�>�Q,�K�C��j����4Q]������%���m�=��_�[����:ڈOgl��k2/�8O2n�jc�b�F0�w����dr���S�ᑱ��ȧ��A�Z�I��Ǖ��e�a�)�+S�}qR~ѵ�*�
� :'���@Mi2���3�hvb�@���Qty-�U5��8��e z�����c������S!�J�=��B��(w��/��vd�������oQM1��"�7��ƌ������;�{�ŵI=��O%|�[?xa*���d�ߗk����E
$"�\Z'��4B�<�8\mQ�B\{�"A�5\�S,���-b�����y�PT��j&x{0��Õyi�T���vy`�﯊7����_	Y���H�Sۖ}3�f��sYk&��.��`�`Zɺ��g��F��m�;�,��JE��݆���=�Ť�P�*��0:5�-�-5��l��c��.�򝑁�]�!��bEW���R<X��-&��Y��x<u)�~�>Q�������2�C��P2Tn`��"ܝܷPM��k���B*oUd~�����H�������2X�u��.�����[���*
4���$*-	#Hs�R����f�OK^ך<*.��m�^����Y�<2}��һ�f(���ͩ㺡j�.����C���W�{��آ`���e�����l<!��kc*1:?`䧆�DtT����{��"���v꫾�h���!u
n�]l	~l�%�Xt�$f"]B(���LQD�_�i�7��r�ז� tx��..�-��#�O�_��p��ņ����R�P4�*�]`��:���2���٢��[�}��H�O���hu6�����@�� �T	M�DZ�4?�g/��r�j�^�IZ7��q�d���N����w�}�����3� ��aTV��$kXQ������xSy�ˣą[��(���.0:$6���Ŝ�xN f���[zE��Rqr|��^B�J7dOL�ҁ���hYi�^��h]/�ƹ���)6Yx�s)'��!.���K�� �כ@R��P'���O*�2s��,0��or�L)�^�E4��6Zx��Z_g!	u�a�I�]*�<�R~����E��"��?�_]���A��*�*�&De��6br1$Fzת*���`^*~��u{#���_(O�\}&ޭit=���T#o�Sl�Ӷ�
h���?�B��
�$��B8ٙ�B �x�R_�Z0�6��:�X
K��i�� ��ΰioa[��q���Rn(ӟt���Q�<#�|>F��2�]��_�x��� ���\k����2]j̫��x��Rj�0U�P�Jj���Z請e��Ӷ�8���Ԛ�+]���X\:?������ZP��]��i2�Fy�Ia%|�\�<w����c���m5�ɶIy;��wՠ֜���n���e����YA�b"�2;�Y&����:���~���E�A��g#�
l�Fe�8����G��=�6
ت"0�.�.LDW ���:���J�YnI�O^�l$�'M�D�b�m4(A���Nu�����\��D#��������p�K�̾��l:���M�.go�������Ʃ���{��E��������K�+�	(ƔoNL0�M�~�x9*���J�G+s^�ڏ��р���M��g�Ƌ�>�5�,��j�~��S�ݴ�]CI�8�lh?��%�ʚ~��żx{D���}f�ٰ�Qf��Fw� �r���%/vdEӝ�D�1�����yT1b1i�����0�3%�!�O �e�kHD�j>�b⻯�~���^��G�C��H8H6����~s��
��gVJ����BF�nCX�0q|;��. I��)�w�0i��X�E42�e^{a�C��0cOR��N�}Zmڎ�6�IɤQJ��;G�F��B��g::��P�$�c�tֳ	ˣ�����C�%�g��7���g�_ћ��#ܖ����[Z����~����&̼K@B����w�ߴ��<�?ka�"2aq�Aq5�k{�������W��oB�c �$�V���W�p2�3�kAY�m�AX��˟Yj��47r�a\)��P�f2�]���U��JTH���� ��\
�4��Pn��	��]S��x�3���,�� cσl*H)�9��'�5�_�k)D��g���)����Jf�<z��F�d돡k�K��3��woS��=b����)���,o��@mU"`�ϓ�^� _�'���[���E��4��0F�`'�s��8c�󘇙]qbh�YL^����V��z�Ρ3_��0�R���`�c͏��6�y�S����[���K�>��7�1��x��l�L�^Aǫ��_�@���m$f|}Ӭ2H�GӼ�G��Id7*Nk,[�ְ#�ޣ_eȺ:Ζ�q}�ð�e #2`�	��}���`���$4wa$��?|�U��P��ٷ���`*��G�ܩ�N�C���|�X��Tk蕣P2�xZ��C���f�����f�R=�tz�L'g�������
��>����vC+���o/�-�G̍�xJ��E �Z�t��� u:��r��V�ri��fN-v�S�)���g�@��c*���T�l�n)~$^�\|���)�e��)@9���su��U�,���>��x�p�.#T�p�&���2�IyA��op�]�uC�@v�m�P��m�#���Ow��T[��Y�i�!�Q�YP�ͩ��{��T�$T$Ki�� :Ȯ�4��O�x��~����=��,�b� NS�*q�����y
I�}�E�����<4IUc��U7 �J����4d-�ϯڀ�0���5��+#��1JЊ�U��N���Z����Kӷ5�?��/�y��]z�ڛ�����(�1%�˩�n��E�7 ��Z�-+e;ZZS���%O���Q~���a���§�f��҇W��{��������b0)��l�q�O��	=��6T�3M�3����'����&����k�7;�/������{u�^�R�&g,�I�93��Y9Ec�����(��.(8�.U���ABfb��y���iȌ(��en��3;���_yVg�(�R�Jt���H:є0�U���V-�Yg�/s�V�y�oj�MY[M�}�ǅ+'0�ax<���YH�����zE�YI��/r�c�i(�df,��J{dZ���ɜ��
r�cB��BM��r��`	*zI��v��N ws�3���W��Y�0�pѻ}���u�_�$Ӱ��_�џ�<�zhv(4�T(���8[9
����r$�t��׹�/yu�#\��)��Z���A�������U3�d�VT��'���,�!#f�}DlH(��8��Q���q�D7A>��"�����F�^�_6F�2���6;�����+J�z�PV�lY)�o^-��
Y<�ݶ<���C����UtT�#W/�s�h���quf���?���1�>F+����T�t�ݚ���-[�	yY4���0&J_�t�@���7$��8�d�P�e�o�ժߤXT�ܼ�-���p�ќ&��s�7���9�u��
����u�vRw��T]|����h7C$�,Q}�{Z����(�gy�<�}��F�ר'!� X"�9| @H�3��.+�鯧l.1ϱ�X;q�ڽB;N�4&����b	R3���J�֞�f������	-�jl!*:D��a���Wr����^3�0n�f�eb<$dcY�:�V�����\�R!5��+S��^�ݷ��%C���]��I���<���X%P���Z���+�k�=��a{�C��sPA�QX?
����e�9¡w[�,�9w��@�9�7����Z&��	��f�����^���(m}"�Æ(�i�������4��.~4Ba?�%~Z�4�������Ϛ�iH��v'�o�$�D��ͽy�ʝ>����a���ˍ^�����0JPc�]ב�5qm�S+Z1ݸ���1�ps2��}���r�ǐ�g߯��c,<�)��?��R$'ҏ�<�>���:K��'p���te'g�x��C���7���4����W3t��x�"<X�+3d����N*~WҾ�rJo-SY���-s��|��fqD��%W����w����;0��>�0��mb7QI�q�ݺ�vNd�����9���S;,Fb�c/���\��;+�4"�n$�7�*|¤��vH;���\�(��K�ٱlC��#0�&�:k�/��]v�ȿ祴)2�o��#���{��f����,���M�9������-A�C3���*�����e���`��q�i�!%�u�~K�!QEnQ�tT��)YSWc@#�kj�s�(��m�[�(
��gڸWmٲ�����O��%�cʃ��Ӣ+�Ƚ>�g��Q"���SB�mK�2!�*Y(l{Őछ�	0�k$�&:��z�sfU)2�Qm.��[=�@�!��nm�~��JbzJ�Ӧd���T�U� 調�*Sx>���Vi�q��^ST�R�9��2��SMF������v��W���!!+5��^N/���Sv��Ϥ��X���U|'�5����;x�`@6pN��$ǳ
��;K�'�^����i��AK��l���Qb~QB�&�c�l�5���G��3�)����T%��B"O�<� X�N@$�i*k@c�y�rˆ��<}�^%Wԅbk�z�r��@��c�=����역��ЂV�S�C�����[���Iu�d��E�$J��Q�5�(W�����Ua'���1L|�w@���������./�\-.����I��簝o��oƉ�!w��]Vxj���F�� s��04�w��̶�v�Xi��ȯ}�%�;'�s�����J�v7������@Q�"/�ujz��l����T��/$�}mt��V�G����l'�(	��G;٦�t�{|�B.�e;&0���Jl��4 �6��>!C;G2,�;�#�Ԓ�%��[ΦX3�_��	�\k�{�U�7�w��E��Z"T���M���!��K&�}��Fy 9���ޜ~�Id�b�|�D�t�\ɠ�e�k�t������	�����aF��ʢ��z�@N��7�݌J�J���=N�� b�^2�~���~�4q)W�(sܓuļ�.(]�p7���'̂�Gm��m+�hX/ݲZ��S�����0��3���3����G`�De���z�|�*���yW]gͪ%f^LA��a��ʻ�81��Q�Z\��Q�"����n�z��6�ԅ���媆tS��NP��J<L̋�W� q�P}�|��ή[�$S�A��=��ؽ:5�A��亗��K#C�
�xK�I0�RE�*W��	�؇ڞ���ÓF Qkk���h��n�����vR���!?z� ��8e}&�p�0���dl�I'�@����xj���̛c�?6"�����jo����
Ѧ���p�N�>���J��%��=�=A>���>�6�9�1��y�!2�~� � �[�J�ב�	���ị�k�� ;���>E\�4�w��	a���a�����ir�m �U�9�`&,�Mi�x68B�(�x��ki�&�ݲә��"��C�|���u�S~�'�N��b�3�V5�m���A���Ԗ��w{�t`�Ȑ����Mh ��j������jA�˥ɮ��aK��=�4ԉ�薫i���ZK�����J(��͵I��]�2ݐ~�<��x\BK�dJ����I�̒�ݕ��F�く2p&�0#��?OC}y������q�ӷ:_�|���O|�	U���;E'II"�D>t~7�s�?���d��x�x*��b����x;�dd��:�{��Ṕ$���Û+���a�Wԝ�r@�@�O���*��hsX�aޥd��O�+ ?~I�Q>�D��v�{Dn`j8,�T�y��P���nr�j�]}�@\H�#���������D<<��U��w[��L�/��[&յ�o��L#�3����
2�x���i�%M�,R�F5\�x��OZӅZ�ٗV!Rr`c�iV�ɢ�x������6���r�;ݞi⡹
4ֹU|w0��L�.�;%G�_�ҡ�5��3�yl���(��,T�H��Vc�
=X�V}`^Q�gS�\�<~A�Hk��D�9�$��YD��_ƛ&D6,��B��}����}C����\�@lr��P6�4�~/
� ���}G���Ӝ�c���@�� 2�fZ�l�b�(��4j~c��˦�Ef=G-�k8@��c���p��c�9X�B�}p�ܵ��Me�f�}��#h(�K�'Ί @��S��E�C��[RG�	6��s#�W��V�ݱD��L�Ϯ�7��~���4��O�O���	>Z�Z�`F�O�꫍�k��Xp8��� jY��-�o��n�LCtF;MT�0���$2��q� �(���Q���U�8߇ 18�s�+�A�����􁦺�.��#֖�68t�KY�i����%�b�p�-�g5�������zn'm'�W������Cw���P�5���]HG&�YW}dR��G���2QvZ_n���m~9lI���,�?`�'(g�޹FQ|����s�!o4bn��T�x��6�l�afy{Z�;�ւ�B� �DSf�XG&�8JG�@'t9�m�� �sԔ�Nx�.v!�,���O�t_���݁o��P.	
T�~K�(��;�́�G:�h@�N�Zؙ��l��r���eɒ��~{���e1)��g!��}�6YV�2��� (�^��&u�����^0�d�@�H���c?&<0��ig����lH��o�?CD�ަ�/S���:yF�ֻ5�#0��y���{�J����!y�[��m%	�䲭=�H��#�JW}Y��QcC�r�����j	Rs�	G��SR�1�^��H���Ǝ��̀q�h�ZXa�0��+?������-N���b�ǎ�=Qc������gI� �����w�m����P���3L3]吢̖֓�[�B���D�m����h��?+R����S?64"D��{o�����zª��(/�cQI��eG�#x߱ �{4���%�w��bL��8�_�����$�E�����nt�b'D[t�+��
tGVVL�ܼ�����b�ef�Mr�A���mw)f9��V>5.wQ�a(���"��M�i�,>���Nbx��>ߝ9�\�Ƅ�Dr+j'�����~hy��v/(c�X@:ջ6,Q-aՙ��X2����?y���ַ��������s���y)Jn,>����긄�b�m��8ʾ5Y��v`/,ߐ�����3 m���kk�S�ّaf�9�,Ѽ �s�l��'NӼ�����Xt�L�b4�Yf�\ک���[�I�t�~�fŏ�m��>��A@����@��v~a=�T+%�7ɬ��~t^�)n)W�'�;��l��@��l�V�./�{@��X����au�~��1C�ٕ�ad͉Y��ǆu�4�}
��EǲK\��QJ���_R�d��� �4��f �S��S/�r�+��O���]7�c�)/��XToM�f� ����e=�~�&Z�x����G�5`/i�Z}0���'�G��]�ǎ�D]2�`����m48Gn����*%�r���4�s`��9��J���u�ZH���.��.��{ �;��ܜ6��S�HYx���D�����*tP�`+�C^k��X�!�d�@��f��f�ۗ�V����Z";i�.2�/��7H�	<�^n���S�PkL�#���a��9)7�a���QbT.�`!8-�?�	�@�R-�ѧx�ېx8<1cJ��5>�T��$�&PļĹSa%��D�[%��&�3��nv���^�:�D>�7�w��3(-�N�V�s�gN���E��(>�E�S`yVL������Wv)g�=�W��C}��
�R2��u���c���"�x����4�~�eB�tÇsŴ"���3w0��3�o%��H�dXw�A�ڡ-h���H��({�����'q��r'ֿ����Yh��<�Ԋ�5i��ΈR�b��43���#wp�')�O�k�QJ0���c��e����Kwc�,�j�����"HO�hwD8�^Rk���J]N��7�k+k5oC���B�9,qP.��l�b��̓�[�iT�` ���y��Oݴ��)zW_,6\��`̠�x��0P���z��2`ݣ���2�6 ��ovsde�\�e��P'��6�����䰙��B��!�%l2�����y�����m�0.w�A�ȍ��q��3�<�%5 ��� ���e�by���w6O2�����v�z=ȶ��|��_��'aD���l T,'�����f�5h{Qoҏ�H��0����j���Yf6�g���^^1r_d糮�}3&L,��?T��[��!䫍&yi�*o��SVJ X[����/��-K��dev���'H2��L���lV�'m9�``�BQ�����ٝ��:XqL�B{�~��0�Wy ��"R������ࢩBBy7߈�з�?T��}ɷ��	*���~�:UT.׺�9K�&G�ᨳ����הVb�CAD����CuC�"����D���+�kuvQ�(�tԬ�:Y��h<LO;�9�A|p��B��S�k7�\��B(xfI��}���g7�����I
@<H^р�����V���MpZ��uh?'\� M��D�-����S˱���.�b+��N�P��R&��?�9}*\�O�������%U��[$�:k�D|d)e@��Z)��,il�W(����Q��&]o��0`��"����Es�d
F�^L�H���w�6N�o���{�^(����������,��>{�6G�`��CSq���UA`�7���OQ2�w�b����tL=��P�ds�C�S-u0��^Ly����p��ʌ���a>���^xՔ�v��f����լ%q�x���sb�9���0�ͦxF=w�)̆��@WJt�s��<STH�-�dI��-�.��n�(��-�e@Qڝ!#ީ����n��b��v��N�󒩫�:J������1K�x>*�Q�Ak7�k�Z579)2O�n�$[C�A�\��_��pKzZ&��縕���b��Bj�K��������R&���lZV��=ܲ3}�>��'s�aD��F��F�6l�6����XA]��i�Z�!JN�����S�u�(A#(e��%��!ӿ��wBS��В�%D�� t�>�A���!�{iEb��N��ޖ�5q)�J3��N1~��0 �k*6O@v�$ľ�O\��@`r�=��,�~�ɯ�2ƽ�?A��Dp�Y�to����،���K)9�5`�큨}dJӶy� ��@z �f����^�SJ�s�Eʴo��BP�� ��`5��	}Hf�D�V�[�8�}��EKz�c��(p���;�:�����M��>m =r�)�YQJ�й6���d�<��z�i�/�Ǹ�x��4��Q��@N�S����$���*E���o$;��Z%��5˹�]�*+~`��R�B"�kՆ���ʔ}�OL����Z��?�)�0 �)b��;�|j����c�b�
��,�"�O�
�;�k��J	��;B��޴1ɀ}>��qz��X�d2�9з�i�)�T���{����bP��"�S\݋���k�Mv�@��$Q�GIm���s�'����sN ��)s��'&$T2?{�@.����k���u����߂������T^��l���zִ��;⽷��${�4��ʓR3�� `�Nb������y�Rl$� �哼#0[��6A6!ĩ-ϕ����������&��d�4T��*����7db�0CS�D��;r�I6_��V��6ѫ���&��.Wa�ť~��v~o�J\%DeL�V��H���3:���,��86���x�EC>��	�?�r<�T�j�����>!�H4ͱWy�}J�h���Z;aڜ��,�J%}��0�x��Y�T�/�1MK�2$��Z������:qԅӒ���&��z��h"���b= ��Cl	��QS��c}q�p���OHЃ�.��?�fCV�1>�,���(`�?�T�i׭Xƒ�?��*������{f8�J�0A~���jڏ��c�?��f��K�G��>�b��Ĺ�`r�.�Q�8}/����?�gG�}+z�.���l�Q|��^&y�MO��@������R�:VOf�����Ȱ lCP��Mԥ��3�$�LPB�=��|C歆=a�cE�^ad������v�z@h�Y�}���d�&Od|�h*�̥#tn�;��q@.{�ϨU{�p���;x8&�i�嚕1:�Ȍ;����]����vK�� ]H��7�I�P*mՎ�]R���'5�X@�kA��,�i���.L�:V*�,����3K�.����J�l͉[�&4b�]ծ�@s[�z���F���
�;,]6%��.�T��]�vvmB�A�a&�J�2TWl���~+������>DD�ۮ^p2@��0$�m�c��1V7�����x�*�w���`�"�Jgrqv��
Գ������:����zs���}2gvV7ll����� �%3�P$�����A���`�7�x���lV�T�i$�mH��A[>ڲsx�k�FdQ��d���K�W���Gq����-B�͒��F��i�6F)�'�p��D�"oqy.��O�Tꄰk��<Y��S��"J�#�qN�;yN)&������I�K���A��=z�n�|f��O���H��<ۡ􆐛l[#��M��wi�)>�xo�5lM���=2M`�3�:2���?A�,v� �~���<�J�i�?��da�@�����BS��H@��K1H��_5���`d-��zl0�TdeT�!x��\�N�,^?νBJZ��[ۛ�����(�sײ��=�fu������5�pR�!�Is�Y�jTH�jYSu+�|w:-1~�y��8���E�FaO˪��U����s�P����Ljd��͸��2���N�K�ye@eI�?��`NCc4S�ǝ���\N@��=3tH����[��2I�C��#cmz��'��xX5��By�\��rL���?~��OwI��7@�(ڐ02�dǧ�N�!c��t"�D��S�Y��d�$��t"t��O�%�?&����v���+B�!�-�-�Ď����-*`:��N��C x�`����W��u�sh��6�	B5�l�+���R�90��;�`���#�l��s}_�㨫��y�6M������0��Lǫ��p&��/��RH$�E�CĂԟ�����?8�3(KF���o�`܋7�	��r��3ك\1T΃�j��;ێHҊ�9�ĮH&�$�(�ro��K˹B�ڋ�6�ۯި��w]u��晶�(�<ҧ �x�" nc�|֞ד#��.P��sXZt��Ph�З�oau�T׹���$d��o�
\4���S۵a��l��D�ϖ�Nj��v�$8��J�oj��g�<`� R,H�L�CH�J)5��L��!d���c\
LG9�|�"ZRgt>m�8k~S�Lo9���C~~p�F=	����n��8��V"g(T������G�>,<�S/?��O�ؗ��8Yr_�)��Ϭ���b�t��m�("Xd�/P���^"s�W��>7��9L�w�PC�1o�i��s뚑~v��f��4��-G�'b
�Z!�x��G��-�O�H�^v˹k2��~�L��p����,��q���#��|@ĿKǖZ�V����F�.��Q:H򅻮�=���u���2���κ���3:\'�8�����e���i�����NU�̜C�&��G�C��G��4r�Z�3�I�V+���EI�[���K!�~�i�!d� ! ���t��[���+�g��jĜ��ཬ?�A����^�&��b�b@���j#��'a˾�q�ؿa�!o�[�$w�T��ؿ��ma����}Eû��_ӎV%U���{�B����[Yiz*���D����n㘶
�)[[���K2��F{�g?|��ѣ�^t�kğ�>��owUr��Ygٛ�᷌Zt����$E�`�|��k��xy��� #�Z�����e�$����]�b�q�-�[��,oK
9�F�5���,��^���c�(�~���ΌY���?���\&�n����4�Y�t�!{7�CP.��м0�Ĩ~}�C��ǔ>.�)��v��Ԥ�؜\��,�#j�?@F�kI��w5���/-� ���&�^f�T��[��.Jy<��Ú���e0glGR��z߷���J�]$�����bA%�[R�k��(�b��_��Ȗ�(T띇�g."?�P�cz�$�1��kڞ+L4|�$��0#m !)��{�3.�T�m'�i`�.��P#�<�&������r�L�2�N-5'�pI�^yĥ���g����9���x�!��Tf��\M&���J`�e��P�Ҭ��B���5��MnXWqя�=�+L�k����N�~0#'��[:�ë��mq���I��6�R���_C���}�BeEM����H���D��6a(V�� �Ɛ\۰��W��N�V>�zu�CxHu+��s�d��'�H(v�D����(�"�0o�wc_��CKP_�)ʣ�ISw1h=V�������� YRT�}M��I����M=]CBBY��R@��&�wo��LQv����-��I���IE��}���N�l�T�\���[|�p����._�O�zF2�C]]��>u�­���4�_��vI��I\�I��_���<c�J�A����i�DTf��w��ػĪ���ĥF��~���Tjn��/�v �����;���`6����3h�՞�z�-�;5��	�e���0�UBpA�{��4_-���2v�&���>�FĔ��̷#e�L�.�VĲ�xm}AW�U��z21�ͣ�~��Z
�]s�^���#�5�PR�v�����=r���H(��?q�o�$�����l�9��V8U{*v��F���N�@�K�E�m�'%�y���ղi��Wh+�1��Y"o�e��ݺ�6H��bP��[	�i挼��C�:]��K�	S�_�i��c;�ހ&x7�!r��tҘ�%��翚�3����UB�;j�Դ�Y`�m����1�������j��uFǤ���q��ل��\�-{�	���������OA���r�l���(>ȃ�e�q[�R�@�0ZP���|*�y�DG��P��Ն6xC������/]�+ݑ7WY!�9��e`���\��+ϋ�Y8<xQЕJ+"�y"����mh;cң_1i� eŃ�р�n�M�3
q���@8!�D��T�r+Q�y)9&���
5��'4�t#�H��"Nk*��|9u�p��y��2���b��F"sj�"����<:'�d��oDؿZN��gm
(�N[�?
�YJ[���GQ1-}L�d�� �n��G* t"��Z�� �M�g�FO#��=$\?��/�����&�T�T��)�����`�M�
�����8F�rkbŪ٧4{G^k����D�*����Wh)_zj����[��/8��A��c\��}sl�W	p����	1���_�j�^�,.�gQ�S�-��V,��!q�h5���0SϮJu�x���փ1�R�b/��L�ٱ����i���G��V$�wX��:�b��G�-��wq�?�\�i,�S�� :G��X��r�m�f}Dl��Ks�+~��L�S���h���Ia��y�'���j����th���a�#��[���8��?��TuU�!��M�zvЩq���W7�0�ͪd�;>$���A���\X������DOhy�nB�3p�M\��B���Ւ��MP�{�#*+�>���Π���̏L^뻳EǪ��V&��D�f�`BW �Lo�7����a�5��O8��3���=��O�eD	���{��I��9���9�FP�@K���D 4L%��ǲ�u5�v7=[��ޛ�иD��m  ��<V2�~��������-q��F#%�ӈ�/"	� �V��;�'�!��^�=A *F,���h��	��3h�G�$\͹�L�;���F�&[N��C=+�ȵ�}�oE���ە4��W�Z:.^��ت��p�\��Qk�p�L��
�!^�?xD�<�v��v�{OQ�z`^�(�4d�l��6{t&7`�|���-e��{x*^nG�Ƞ�7�����&j�s��U�l�s��Ӵ�o�>ja!B_��k+&����zJ{\��KSh�)�=�´��@$�ц��H�	Y�^D�?CZy����|����ؖg�|�=�iH�h�ᤤ]Jv;H��28������
fȩ�f#�|��j��8c� ":�N,5¯1i*���âvm��T���(Mc�
e�� �7����/�|���3+��{�
Y��[�RW(�����#S����ME�DG�4K�����h��f��"����!�Yv&!���*�R)�}���bE�=ty��o�JBn�yx�+�db����Y��m�ǝ�K����<ku4F-bq .n>�a��Q.:8�z�{���R�G�A�S웨$#��GR�k���K�I��?4B,)x��]]z��@�i_���bҫ/��b�+xy�1ifƸ���Q`
���	��-�z�^���O�к��{�VY��1)��x�_ClN@MscK��}q/�z�9�z��q�@(O��E�stZ���a.ח��[��@ �f�Eڰ� ��djk5 9$K�Y�R�8�	VO��1��s��3�;"^�;5�Hw�yI[j�/�Q�3624�����g֭�b�+Ȁx$Lz�8�1U�4�l�O�FI��f�pp8�փ9����}��e��E �}��밮���%sI��82.'�U�o�~g�@����=pun�9ʳ&RW�j-��S�X����y�b�H�^����(�������a0w��o&-ڋ�^a�~ʸ%�]����4?�\N^;Y�֧���O?�E�T)�z�=?���+t~=���An��f������P+��s~�A��6����R��m�.�������Ϙ�Ӗm�m�728�`����W��n�	67"c��T �"sC;����V�b�@4/K;�{O]I��;��� �h,�Y_����c���tx��8�O2��0uFS��T���<�������Xe�įΡ���<������S�s�s����$�>�����Ϫ!M���m܁$%1A�;`�3؁��(�53�H����D&��k	`ߋ�q�i�_�{V�GN��C.r�*��71�wsh�!S�@tE�m�L!�|�iH^����-��~'EI��R����b�(�͆�Z���-	��K�{�G�˯1���-��1��v��tL��꿔����>�)��{c��@��>��UI+G����[��/ע��7���9��ϋ����r��T�!�8`���*��O.�\jf�	5c�ΐ|��1�N"f?$.�5ꞅ�@,� �����η�AT���� ��8�nt=>[�����^"��x�IV�Z��@!��$��>��d��in�հ�A�7	�B)}GS�&5e��d�6t���D(A�������Zё��G ������	 0��A�_�;�C�ש�����a4��N}��ђQםwE�ȕ�߀P��|�ٌ�m��/���^{5�.�ˏɶ�����XșxJ
������>�D��=P/�*~�� r�c<�nGΜhUE�E�	�DS��M���6�!ɹ�Ė��}v[����=훬4ӺN:�lt�+I��^D���#���w��D�c{�#cƄ��G��A;c���my ���-����d��G[�4S�I}����[�����J^��0�ޅ����k�����|�6D[&b����)W%�?\|k���g����)h�-#ˮ��>�����o$�u ��-4�Ed�:�9������R�����9]|A`�]p��m�)��#�)Υ��7h�BKQe�=!T��'u��}�[�H����fJ-ؚ�9:��Dy?�?����B���%�G���"�C�7����Vy�,��{ۭd"�
��Т�ur�:B��bpo�X{�"y�XyA �<,V�Fx���4k���i�ɬ���gkB�
�,^��b����<�n`�O��{���H3�S_�r����'6�\5�f���:R�f҄O���v�<�v�ӑ��T�j�W3�Bv)����2ᗠ,�BX}�l �H�Ǝ7󞄋��8e�yI�N�����YGA:l�h�3��2|.��V;1Qr!g�*��\����cՃ����f(�lv�����W$ݬ�9L)�82~�e;'�!ВH����;<��`s�_kkkl|�%����iX5�hX�I?-�X�!#w϶K 1���\���u_�
k#��cm>K,�Q���������"�C�U�2��6����ՠ,l�+��<���<�Z1���ܩ�mh��U�?�@��)��zp���CD������gW���b�(;��7��5���e8����Y�������qe��9KJ���
�0R�UP��(޹'#Ή�V�Ж�Y����h��-���ٞ���S��~�{�R�$�o{y\����v4�+ g��5��u�g���3��Z�w�J��@�0(�]�*l|�3
�7�������t�y���eJ�Z�.���1a�7@�L�P�C�Yz���U[#�o}�BЍh�K�'�h��gQx��F6�B���1�RvC�m�'`ix�����[V�������⟾�WI�����F\gV|\Znj�T�=���w`l�sKަ)n�ߘ���h�c����ޏc� ˭�}�eW�m��޼.Z���說�vDFl<p�}���]��u��Uk�ҵt�H��WE��l���Ѻ� �-m�����1s@���X+_7�u�u��=�O���UM�v��:��c�,�q��2����:�^�� �+u�x���l74�;I��\%��l Vt:^;���`ƺ�.�����tW)F�=�	'���߻v���5x��dk]k�c���v�a��M��j�ƍ���w�����f�f��N!|$��:8pr�֖�P��K�t�Lo�/PҔ�@��{ݠ��0y��z)L���I��N.{Mu)��+��VY�	_�#m̡;���pP�+v{�:�����g���e�D�S�!�}���̺��k�JL����Gs�V?��c��M>�nc2�U.�D����?���,��Xp���%���)�vc��!_%����G&/8M��v�/�2$��8�^�چ�`�3JL�+;�0��YW��0 k~ҹO��N7?�C��!L��� m��g��j��
UDe���@Q��c,�d�"\+4�)�x����Q4�7Z�5�M���dBwcM͵o���	���*��=1�;�G�դ��)B�'d_숛��n�C
�I�֩I.���e~,U�!jlʙ���N'k& ���므+�%
��h�q |����� ҇"U��b����20r�����|P,0���Ls{�9 ��|w؋D>��w��<+�����3X��|⦧eXڳ�z�2`W(p����
���p@"M�M�6�O��Oi[۰��K���A�X˧�e=��Q�������{8��b���_ӋiR
�q)÷�W�Ơn�M&�EgXv��Q~�s�t�4�Z���vc�s�d�>������v��3jP]  8\%�I����c I�6�|���<AD�J�/�O�yK�3�l�&���VI��!���T+��keC_uGbl��!��Pg�mBs��;�l>�j�z�4 y�I��
�˽#8���'Y�}?�c�mc$�>���\G��I�69LB���0Κ� �8�j���ظ�@(�{���䫛�1U��>@~��5�%\o�=�%IC��A�٣���ݓ}��1c��d��_�G+�JS��2�{R&��9	�l�!lُ�*�kA�P�/��Xk����RR$�$��	�3d�>�9v�� ��lp�p̞�&��oJH�T��@�cEԥ��-U{W|
�g3M�n��X~��G�9Ʌ���M<���'���y����.1��f��܍w V�������JeO�<<UK�~���>�Wg�)B�U&j֣� �)� \|�g�[^��d�=D|�"⧸�,�G�#��-F9`a����hp�,!(���#��k��(:g�d���#"����m�Dt�
�X�61Z��[�*b�:-��4�WD�����6S��s:U��|�l[���
fV���ω7����w�;�(j��`�2ڎh�-��
��]V������"	�D�'!!4w�h�y���6�]|�\��v�SF���0����\���=2�2��3kK'|W�X��2��d��FOܰ��%Kӯ���O�M�'"s�gU�,�觡ι���G�o�m���F�΋|B��:n�
*W��5�-?�b����q�0	*�QD�ݍ �j�e����d6ﰐ]�ќ�Sԩ�q�z�G�𼓿�?g��6�c�i����C�w�,f���d��
<�?��I?������%od>�K���S�Ja��38��͗6�}�܎hmx�U������@IV|�&6ώIJ���:U�*Z[x~�{ͺ�y�ωI�=KP��{??ue#��v"rG�jɨ�G�#,��ך}�J�!�� ~J�sJ3�ҒL�O?�L�W�NNȇ6�H^9��պ ��L U�.?#�CΨ���>�k)�'Y�Y251�uZ$U��."����vǖ%KW1Ƭ�}p��P���+���x^���1_v+k�ăe�2��5%���g�K����K�1��M�DڏQGP1��'��foN~[?n�X�F�:�=jƙ�s�� =מ� �ɼ[HM�d-��#8�P��M�����z��H
ȁ������PQ��(�JaR�n�<�������ì����x?�+|�XÓ	��m��!���g��IaK{�vܦ���*|�i��z~�/�A���l�l��޿cOmn���f\��@�}����+w:������D�i}�$7�a
K����,�L�~�[G�Ua%�Kzy�(�,Q��M��?���>�*���?�{"j~T��ZtE[��1��^ۘ�3���F�k�;�<Ta.{���"�����l��7�絹ƼN��j�B@4�0��Di��Ÿ������#f_�w�����>*�V ��r�!Y{��>O#:�
���z
�UpN�.����YIZ]�y@E��-eOTf�W���'�Zv�Y]��Q�_�9��ϡډW�idy��)�V��pj���z=$�Cg}e!�`c��=�n�$k���j@�Sl�2r��Xߵ����.~Lݵ+8�(F�941�=o�6T\�e��*?=ẌA��Fs�����|f#�A��qJx{޻I;s����I���S{,����T`k�G:��.�]�v -�,$�t��u7�ƹԶ��,-���"�����
���X{]o-|Es��P���0�:�a+��:����Сi^=󕖽jpR�(�3���NMq��*w|�������t��޹DU�3�#2~9h"��Y@���W���CdsJ���%67$:��Jn���Hu�d��+��'$�/�_�ߓp��x�U�>L��Fk�<?��	;58�
�����[�2�T�qK��Ә���������)���`�[rZ�xX�j�R"��4O�d��s#}E��ap�26 ;�
���y��pғ
.�ʱ��w|����$��t�GPB8��Ma�f��	R�z��t8%�b}�~D�BjN
S�}����@�1A������,���Y�Iܝc52T�X�蟬�f�_&�RZVy���vv
b�&`����]�#3��Y��9�A&C萝�(�`f��{�5N��$IXo�e_ɭ~x���^�x���y���y��r�]Δ�/��U~:�\0��IQ�&�Y ��[q���pq$� ����m�P5�x�"�@
z�ē�����p�(�8�LH�
ZFZ}#H�ח&;�|z7�j�S��ßF�'u��Ҁ9�p,��m�Vb���s?��N�쇯��C����e����6fA�L6nԕ{�Y��9~T�����[�����M�5�պ�5�����n^����:�7z�د��w<&��M]z8W����P����ư
�D�_�QP�E����k�U�Ǟ�涙=���~��;F��:�Coٷ
\/��TP$����� &`q$�����c<��w�k�H��}�D'w�b�Ī���W2�K��)�^bg��;����H�;��p�s4��<oiV_��0=}y������Ć���[����
gο�~uF=��v5Zz����'�ˉAl$V������6%�`�~�ޒQh r��n4p��}_�ߊ�����u�s��"��ދE�Zw2.O7NO$Ѫ&�N!��%w�v����Rw!i�u��	� l����ڈ!��U�QxF�XKW2�����j�?빑��Ƃ����榴Gfl��fMa���A����#�s�r���7�B�'jp��ib/ s�xRj�7sU��/�yT�w�����Z��q���Me\�AB`9�#]��1 1�f�Y^�����D��"b`$�V�_���B/��8�Ȕ��ؕ�>�+qf=����.��Hh�tK��g�
A*�&�� ��v�[H9�ͦ1�Nb�+ώ^�"�<53Z)�bPq"��t`�@63� �S��&>���=]��}%�I�b��q�������fd����!��`����'��'EQ��t�18�K=H٨{g�P�9�.��(%����o�����f��kP�HC�)�kZ,qCv7My�B[�t���^�镺+�g�����j^8�Ep�!�`K��"L0�.�;BC^��Q�a8�	�J�m�?S��RE$t	�;#��Q�v��������?`�e�8�O��/��w�2��u0�㊻v�����C�d�[t>opK�f����@l!^T-6����o�o�FI��m͒}�K���E�䃮Z!���^�J�,�[�E}؂ �+(q.��p7�= ��\g���>}㉀�f�e���7�铳x�Lf8��`NQX�f��v|$(����y��T�	`��h��輀����b�e3�WEh����1}"�y��<����V��~��x	!G�u�zo��p�;6����n�!�ྻO�c/��P�S����rÀP7�!��)�qz���4>��k����N��t1�A�Q�F�b��K��)De�/n��̐���9mB.g�!�?��]4�=���\!��is&�o���n�q>�J�>��n1}�M�,�^�cr�sEw+��HW���
f�>v��At1V��ٰG��M��r�[CQF�[ȝ"�j��3j�41�~�i:�K�P)y>d�wk��/
2�(q����-�Z���K�S�pD�m�	�[��¥up�uw����Z�^�Z�pR��М��0xL�7M���q�	��PD����a2T?L��Bi�妁T� ok�y��|��p��	�񄹯���v������jt��N��ا���	qC4mPf�^	5:�M5Oq����3��	����V�![0o��<�s ��;���a(�.�,%J��Y](�<2�D��#[&��9&���:����e�����/����J���Ģ&%��L$EМ�����9�^D��ґ@O�pN�X��8CMlT�������2�H�0��i䲼��_��O�ꬾws�Pa�� -Bg�'���=�i��X t�Tm��0h0B��s������0�ce�>�~�Ѥ��Q��r~�"�Y"t�ɻ��V���P��H�#�ʡ���4w;�K�itVh�Ђʰu8�%��%��	r����-��x�/��@ ��ˬ���r싩�]A4@��=�"	���� '�s��� 0�4�O���B��%پ�%��Meh��3"���p򥎖�)�+���d�#�'G����vmpR3�%�P�)5�I�⑷0�Sb/��G�+�8$vS�t,��U����:N�1�:�	"d��$K��|¶ܹ�kv_I�-�%R�����ͫ����S��]~�T�ٱ׹9߮O�<�꼲̏́3u&R�����z���,_�=�43���>�o���ȭ��u ����8��Yi+R#({7��3=���'B�*l7��n�$a��~��Ͼ%\a�M��_��t?l�) �\�e
����5]������Xd�l��i�lڞ���)�J{y��� �G�q;(O���۲)�q�˶P0�d?���~4��#V�g�L.�P�6���4�=F�ԠA�Y�ŽQ�ШD�ݙ��h�0D����`��ޭ�k����Cj��OBň���7XP�����������A��h��#�MC;u�$$N�{��GXB]���ν�}���o���L�� ѥ3_%{h�P���.fg��Z@rL�e�>F����N�u[�֮b�e�-��H"�0D|m�4̢�u���y��'&�m��/<I� y����j݆���5�V�%P�d�ƿ����� \�2`��&�=)\M�pީs#��WT�����M��z$�'@��9nws�0�������y6�3��� E�3��E�G'be�dݩL���{�< /�X"��Ƥs}?z�� ����T�۴�
5��픋�;�P��+��Rze`f\k��<-$Xù$Y�.�jJ-��}�r���?�t���P0����Y���e��^��GXt�^<�B��y͈wn��U��-I�"�:z_���=#OWO��.�}ԙ��~?�u�`-L�g�ǧp�#�s ˫�|��o�,�"]�<D�()��5��]��Ϙ��j�����L+Њ�]�W�0��.�½5e��)�/��wl�߉6́[W�b\1C���a����_� z1�L�EK�P&z:���b[�a�-����5H5L�U����p=�]Y3e�c��S.+�Q�:ȴ���$<ؙ����5%	Z\~�CH����b��<�	�Xl��[!wj�,e,��x��q�֝�&��B��}�Ud3`�u�Yi�������%��*k�+� (�=�Ч�.�H<�F��:3 G�����@(1��aJ���/L��J<[ɢt���֬�B��]�ħh����V��(&�
9S��\8�T<��"�3|�;:�v�D@�_�ښtQ��{<��`$�y�������:��C��"����8�eJ�q=��
]�~X0MW0S�y�*���UټD����o��%T�#�؉����< �c�9�ι��Y�~�:B�u5����n��Gs�� �NX�Z���2b��F[z��i�cj�oDn��[3� t剉Ƕ������")��iey#հ��ڛ�	��&[�^$VDY�̿���3���9Oe�_�H������U�-��}����8'��{��$$DSB>4cښ&��I?}��<x���E�-��j�9Ρ{FD?���
i&e���Q�GBU)���x��S�p)(P�o�NvF!I�	���1|�=��
-�Q�����y����xx�T�x�1G
�z��n��~N;l�_�h�c�&	to'fZT��U�?���7������O
=�	�n�6_�
�
?�KHF��Q9���풟�&SZ�l]���2V�*Kb�X��\µ�"|M�']!�!нw[2�t��Hz��gЧ����;����{�[�~N�����vC��H��*�j$A���G]�Z'j��DIY�܎7T��&-�..�1�>��Xd
�ܛ o��L�~��9"U�;��%d~��)AG.Z蓉CkY�x�>^� �v����2�k��<��He���8#&���2���$q�~>������q��s~P"�g��><j)k3�$�iC3��ܵ�g��"zYu�z���k_��;{�������}Z7F+d��xeGHu���ä�)@�u������9���Pv�]�I3���zF������D<�;�4��^@
�m�uc�c��Qu�Ή7�\�Ң>��'�9�f��u��蔓�aKc�������1A��;%1��?������g|�^!��B��ɡ�Մ��d�qW@�i�5��E�&�� ؅A*]�B��P/W����R��`���jK�lg���
�ӱk�/�����z�h�|�IyQ�8�p���e�|�
�f�l���� ���I���Lڑ%<������
�3A�t��y�M�3)#��-��DСV�My����^�.
�>i.e���\���ǣ4��t�ޔp��P���Ě��빰�c�s;�9���A^�}�r�XՂ�y(�E�����Z	!����~�|��ұW�W׼J��v%j�%0���FW�b�_%�2T�� P	QV;�!���A�9 ��|���y�٥�.lfu�EBӤ���p��������f7.D� P c�З�V+1�Ж��`G/L��&kY�&����B��Ǝi�O�a��KI��q�@�E�G�:�pL*��;O��v%�~q2}S��T��HPt�K*s��yoE�18 gN�fܻ�pJJU���P1��Ӌ��c��ƷN����R�4A�	Xc�1�tZ�[�.Ad�rw;��^�B�	���lV(�����>Yf3�KTcwT͠�� �*�a��|gTE��(�惯{��h�n֩c+��b9c����6��Qq {~8pD�ʑ����k֭�Ha��0SVRK.�[.O��yו�]8�������M^�����"�]��=��]�.����;m��x!�n�b+�At��jn��[zq��*�)ꦷr�Wi��K�ڒ�e�9��jud<� �áy�����LJ��+��|?�T�����*�(+�[��?�4J&��'ѯ�	9մQ�$���b?��̒fi޵O�ڀS s�ݛ�Yg;`�N�
-ڶ�FV����� !엵7����_�_(]���BYQ���EE)�\�����ݵ�b���3̉�����Lb��O�A?�� �Ĭ�N���<3���\��:+�����a�Ԁ�*lJm�K��@�c�����o1��SF<w�	/���I*�ro1l�!�j��W6u@DE��/�ش)��j��O�
������T���*��,�J�&��(ޕ�ڙ=Q�=���~��9�w��.F��r��Y��U��U�U,]
�R�A=F� b�!8Gx��IQ?o�8O{��u��v�'�ǧ�5��ģ��y쑺7ӎ9��p�3��[Ph
4��i �IaG�"�+f`���~��;s�tȟB��d�t�[)�-�g���}�t�~�~�J�;{X���E`yW����ˀ��,nov�]�ow�,�e�/�L�we�%��,ٌ'X�[�<(�K��.��oZ�|;i��(�����P���^���ҧ�hF��7�临�������J�OHJ���;BE�G��Y�; ���MS���mX�٤�Y�f8MX�UJ��Q� Aq��2�r�����)���s��:�'�̻�,
#I �ćz�2H2��q��ĥ�m�2�ê�֛QRS�!\�G u��-�2`ۗL�G�������_c'K�t1����R�xu|6��[O�[&����6?��IX~��R�_Wr9��im1�%���Ki�8w>�A�~^@\��q[�yd��EPVI�5����9��lR��I� ^���LA����}?�9�ynpCn�Ͻܻ��pz�cl:��BE#��?� �a���8���߄��s�G�H�tX��5*Э�X��Τ/Q��6|^��G��|��ZZ�<|}�҈e!�=�;l��j�>�[��dr�s��6�@u��0�Q�&��t�֏���V�����GJw褲<
�巁Yh�m�ʹ��s3ob��A�ci����<S1�$��R��$�+� ��+������8�`y�do�\	s�v�v����z��L�Vm�]!gK�ʑ�t>���׉����D����p�������L��@��䍍I�D�x��R�X���0Q�[Rw���pJ�X��X����|@j>p�X`XC��Lc'�:�����0�3�׻�% �iAj+��ⅰ�E�����T�;���t������q,W�d.��)ɛ��� Q�^�mxlH߻����ND_\��w��<:s4m�p!h��v�#�o��B(�f�8����t�5�v_��*�d�T! ����s����Fժ��x�3YS��h���%u"ox����V��k_~�
�ސ��d���:}b�+���Ge3��y���R�&S�7�rfҝ��d4���x��w84�Vu�r"m�Oţ�1ڭ�m������y7�TDz��:PP���]�3�a�R�������@���F��h���mMXO��N-��mZˋ��*E[m9���W���4S�Ì��ݥ�BW����q���@;X}Q���HjW�u`�Ր����]�5�e�r�و��0Ӫ������F���q�x�F��"�؛Ć�` v��#Ԑ0��ZV��Q�O~�WBW �Ǘk:^y�a���:t�f�>]l1���Y�u�kb�ó}�V�(ҥ����"�,M�yS� �~Jw�d3����z�ιzY�u��T(T�e�w�\u��k]�&��9'5��N�]�<�a�����9����wZ����j�7rb"P"�\�n2��B�{~|�\h�g�X�C����ّ�ۚդ�&7�����=:��X[������{���K
���	�|�����o�l�C��4�1��aJ"������@^~�΅�4�47!�$ �g��|P��#QF\S�#��Z8��hܷ�p�F�A�O1)oz�aU��U�t,���	���6�)���^3{�W�n/Z#2�������>E6I�1K�ߏ���4��rrz�gI5�y�VA>���rC�7�h�M$'GhXZ��e��%k�P�՟L"GhKO�5y{A�}�l��i�z�'̩W��k�cΔ���$~�� �a�՗A7����9�t�K�	� ���.��m���6�r���ˬ��_&�#D���ڰ�~K�甓�S�|D���.O0��Ak�p���, �j�g�6� ���b�������Y��*����yp���r&��ok�����)1�j�1�~[��Iq�u�cP��E�mr�k�G��oh_��u�*s^�gNp����uR�s���>�k��6�=JA�b�5�1hs���}<ۯ�.#�E4v�U
m��{�o&udˊӢSKT����:��7X������MJͺ��_�I:a܋~�7�;ئs��+3�;���'�.N�l�K��&��2��Vd�KdGA�[{NE���\��ypӕ�b7ʒq^����|�,��I��?�\|jz�{�OVF��>S֧�^�Y�X��w�}Ƞ�O��-��QN�>F堔?�[i��jP3w�p5V�x$T�WK�<�/�Ex�}o�Ǣ��,�7Ӻ�0޾k�b�Q87+�D�Al"�W���v��ZJ��h�Ѧ�Hhl?4V�Yr��2�̼8.����S�s���
�\2��|Y�h���鞓d��Bbd�T�+��9P��H�XB��#�,gh�����x�����]��1��ì��#�[H�U��?�⮕;��[�k ��F鈊��_ٛ���R�h50�/�IU%}�9�&�+V���~�Hs7>rB�kA�^^b{�\a�����"�\e�	�� ��Ӝ����k<�+�p���<��t�?>�sJ�H�܁N�z>��8�K����>�c��i��0���p����EW�����}R6Nуa��{�)��:Q<D��'#�dQ+�m]^Ǻk"���4��ҍ����c����Wb�S8=*ϧ��UTz��@eC V�♧څ�BR9%��cq�K���P4�H
_�%�~�.�?�_?cJ ���]��S��*X�5M/B���*l5�N'	3c���4M߄O �l�D!�����w�kg[�@п��yk�r���ٓ7O�S_���;�$���r�����OƏ}�E)��G���q.�ϖ<}��h.ۿ�c��M���o^�2�T�����U��m"����-%̟1�9�"��3��,��`x�Z��)6c~0��֫��P�jxt�a��ʨ���>��Y���b�bh�B�:��b@Phc�B���k���sy�W�X'��ς�I�H�A��X�I�h���{�@�qv9�r�}��ra �w@�M�r�l\���E�������Z ��3����B��`=Xܪ"��܄�/�1��O��m�ӵo� �Gk�I
��N�����$C���*Z�Mxc�g�L���_��{���q�т�Y_��~q��"s���V~� ����Z(+��SF��]�㋉}c꾏����L����=��z��Og�����Ez2m��,�b�������㌷�=��W��Æ��b⓲�D� 3���,)�������w����]چPk6�5PL�.v��$&� ���9���-�$N�n�'������w��BKy� ���v�@}FAr#�h#�Z���T�:�b�v(�C0K������%=|Yٹ�-�=g!qbγ����G����RZoT�L��v�!��%ђ���V�ŉ5-.�B��8��|� 4��R������g���;M:�֣`��1����!���<y�M�*q�$��Dex��v�F�&�-D���ʯ���!�|��c-{��r��d6:���;PTy}��:����?���h ۏ����B�c�)�5�b�˳UQ��\A�Q�L½r�5[C�͉�ȏ������/T2p �m֖(�;�z��� =���l�u4}�A9�|oZE �o k�Y��Ҟ�>ح�)G���G&�9����*�y�Ra�]!L8�	k�	r��b��JL�vB��d�ղ�>2��ǔ�{1��z�v�8I�	z���܈�B�<���n�<�E\��g�q�и}ҐF����`ǰ07f�_)S��������[��!s�1�8i9���t)�ؚ%�O'0���/'��F�Х�U�����iz3̍-	W�B��[nK<a����(��م�;�Pm���f�TayAgs"?��Ig �ϭ���CR������$Z��Z��+���N@��A۸��ˆ����q��Z��"�B{��ga��'d��_4�9W�&,bs<����f��s0��^��"z��u�?y^P���6
�&`M�/�Kg�����v��cϽ�QQ�ʊ���l��.�{����#S��m:Urx�DD��4����;T0��G�l/?I׺�0B�:��}������DY�i�[��'ZvEP�v�E{N����猘��p�[�<i���¶�Oi^dƏ��b�������Im����C��<�0z�b:δ����\�k
��"��Wya�Q�0� _������uG��ew��o��Wf�~xN�7p8^5�T��@"K�D�r;��D1����7�I�=v�ts,gwn"A �7���j0��C�+}TC�cR�'�=|A?����m����}�)���\{��D�\	�qw�>��Wώ�}	qr�ߕǩ&�R�sw��$!�x#�j����b3�����J;�y�u��~����� �]����F�����9����;�|�%���K�H
kM��_J��p~�l����\:���7�p�k/�V�
���3XE��r�F�YW����֗ Iڷ1�l_�'�gJ��tF1`�6�H��!����r��n����9�j����l������� ["��ԭL?�;D�!ڥ-���V�Qt�ȢM�b0_W�����GAp�-Ҋ
v�������X�.WY�֍�dB��/�K?,K[�+�p��&�?~����f�Ǹ��0� X
(�����ެ�3�S��pT�"���&�,ίS��7�T���l)�
ڋd�E}d�v̳L8�$�߰�}�*�<ےG�ܫ�ym���uJ�+E툠�s;G;;Ca0�j7Ǝ��^v9�����,V��r��,��@��=�S��W�0���0�$��[q�l��忼o�p;;�aqt@�O�+��M%�" 6�b�v̻ ��hžM�Y��#����Y
[��q������W�v?|e�x����9`kYhj���پ1���J��u�L ���?Y��y��[���L���h�uLT$��id� G>$s2���ӿ|�'����Es���{{���՟t{%��s�j��ӱ����*�����l܋8�r����;��e��Û���	F����Cglv.dݯ �)+~V�?����b���u��u��ӟ�6�u�09ь������"�?�M2�_��@w�O�݌�n �u?�Ek�X/��Bq������a�y��?��|&o���ZXh��]Gr���x@P��d��� g~����2��7�����<ol���I�>��܃|��>:x�1PET�c��n� ;���� �}�]+�b�����:`β+�N0��i=>y]�:%p�.���PJ�Iktĳ_�OFM0(���U'ee���o�����у5��|�Ua�j(��^7O�_�R���%GcO��&�U�(+���韷P3h��B�S�9�cg8{��u��}�M��B���5�b+�YR���I\�����(ސ�ql;�e�P�J+��̛���"^A�����S8q>��1#h���:�['s de�� 3����#�A��i�����.�m���N�%����:z�`�^��}�o�<7|#�ӯ�4p�߂�Ú�BM☜Gʍ%�	���&������ѽ��8;�o�.��[�O�Ol���6P2r2�͆��{���_���;:���+��ə��b���V�,�:����Vzd3q�,�P{I���Q��G�g0����S#D^���i	���M���-�������ɜ��Vf*���ӈ�؛"ٝ���]1H�\�Df8�/2t0�[��C0���`I�(���bА/��D�bص��$4|L��	Ҙ��= ���G3�X_!���Q-�*ߟiB�!E��*��o��ϡ ^\�bݿ���p+'�]Ci{R�\%hv�׏���L 6V�4��m��+L�O,�vc?�˥�f��-��(�(�Q��HOWO>,�$6^����	U�@���+y}��b��A_��G `}�LF3m~d������&#���>��8��N<I��~Ǜ�p�M)F���{�j�Y�H�Mt�vɃ��õ=��L#��w�z�Lc���%�8�2t4���m��{q9�SjH� 1�.�E2XQ���߻��|�(�Y���h(r}����%�E�!�҅��6~�,keD�&���m�F�Ƅ�$qC&�%��>�����Qu�)�~/��̽��vJ�'_���Z�
��J�~�������H�*�Xz�a���}�����+�n-tPz9�ܗ��v������	"P���qOکͲ~&��u�����BA�X�R�f��l���4O�4s
F$��a\�9Q�*4��H[���1�67ʆH�v*���	,��������I���'?-���E�}$��n�������V�(�f1$n��7^R%<?�~�t�kYu�����P��r�����Yfr�ju/�]�fG��ED`[�&�F�a��{���Î���v�-)&S�yb	��F���j{�����H|q"e�fWoO�����Q�m%k2�p<1���)�L�Z���;�$f�݄�u��<x����<�@�����Ӄ_�V-�C�9t>���5����b�ӓ��}	��^2��S7Ѷ�}�Î "��+��
.��Z&4d����kbP�\�'�*E�ڍ.`~����?��8�x����i
�����P�=Ȩ���A̎����W����-N�/��T���T| �.���R�c��r��<���0�d��Kt����[,�C��SA�RƏ�	DJ�>����_�F�[�C�y���	�)<�~n��� ��ۙ��x���:�}�]A~nӬ�{�A%��Ty���1 \$�� ��D���<��Qd��5�D��u�t
yTE�E�/�S�I���ɲ��=��{p9������O����YC˶ҦB�5�z��s'��ǁS����+��?eA�=,� ���8Ș? �G�22���qw��d����!]}����F��,�3�;N��N�6{>�|G*S[��&�
��NZ��bR�	;�ϫ��a��I�A�S�� ��ɽ�B�h
;�1ָ����q;A�)*㓚4�L������W�5%�ե-Wl�Ϟ�Q��]$��@r�l%D�$�W4�DY�(T���_�N��q�M�S-:j����벟���My����_�����S+*����S�b�5��(�4C��#�C����,��f�]/���=M8�;�l��e�i�)�x���lv�D؞}|��t�(�F�%������q�K��E�b«-(W�6�K�&a\�="�ZX(�ϓ�Y����;RJ��,}ݣ��ż�a|���	�@��O�����|�DK�v(AxB^߉��I�&YZ��;��H��06M��x��]��r}�A��Mc��!���,��,�˷��ms��!'�L�C[wẵ�]~>�ܟ!�9�P���~p6���GӍ!�jQ�*~i�,����Y��pp����5��$1���vu@��`����B��P��ſ��@�_��U\2�LM�+CC��t�+�:���]Ҋ�џt�Ibv�X�F"6Iˏ�yyB!W����#��\`b��)J渂L�0kTy󪡡���?tk�������O!�DVe��7b� �:�#�9&*/-Mzіk
d�,g�=A��9��6�b�Z��ߎ�B�zT�x��7S�O^�u���zy$�wr4��<�I���@�>I�3S|<v�j27�A�� ޿�D��
讟��ܳ)q���d`���H�"(��R�0�3�� Mj�E-��ײ␸+����3�P�?��{5k��k�^�A��=ћd�
<�ߨ����C_��wA`��Ϡ�Y ���9h�T�}�_��o
�-�m7ę&B��Y�v�G��L)��E����&��[����L�xa�ǁ���Bj�gɄ��ZU��� ����w���Q91��Ց������[RK5�֭����@m!-�F��č�����?�{#��<��T�h�.��=�}ؗ|����O�D�N�z��2]��u�<�m "ݑOs{�3�X7aڐ5'��c�g��y�u��&F��ks���~&:?��N8z"�ܬ�p�_oT���CđM:M��cko����Qx����� ��w/��ӚI+��&��Qx,d&��7{{��|��A���?�9�&�P-�4�ɳ�3p��5P�J6��F�L=�H�.��G^�4JX� 6'v�%/�5+]���h_�9�^n�0ĭ������<Q��˾���uE_A�ђ�#�<�5f���|q4�B�+����9iA�ңT,il���P��un� ,��?��+����f.)9�,I�y�@B�ڢƒ��<{}X+��*�(��f�ZOD�9�DjR�����bY���-�v���NX}�9
J�I �(��Ȗ��H홉��~7���7Q�uEԁ�0	�7 r��͘�+�>Z�g/q���N���	-Y�Xw��7QQ�Om� �@��3���`&I�n)�LBSg9��� ���YUޤ������Z�W�X y���q>�!��ޝ�;�ϊ
��d]�:��R�A���dl�Vjk��t���O
B��f̤��wY4�o<�����&h^���hi�{�|�I4��&���S�4En$��$�<��,��F��u��l�����A��A�M��T�a��[�}�yM���7�L ��C��#��?�t4l�ԕ��Uc�)g
�Y�H���d�� �
�`Q���j)]t)|�2oA�)8IV����QtLv����e��Q6��$��zJ�}J�JJ��: �{ш׭ށJD��҈���$@j}��N�!���� �X�DVBA��,�% ������:� �iu(��ޛR)T*'(�ӳ�g�*Ϛ'�d���w�GKz{&t���oI�u&5�~t�/ڟ��޼����a�k��e_��<��i�諾���>����J�7�в�⯴�\�'�-�L�4��8��t��� ��>�g��^�k�V$��;K�,�&i��V/����`<���?�â�E�C��^�h��k 1�{����ٛ� e�ɸft���Q�T����;�&
��/l�wɒ�|��^������fj�*x;2��;��&��Qˑy���}�A�UV�W��Zq������.A��)��Z�oW�fBF	X�i�x;�|�JK�r<d�S�G��2C����ed��ul8_A.���I��Jf$
��%�\�]�rg��2b�1X�P���]��)O]5H̪�`D����l�dm& $ØU��#���e�C_T�G+3+ ����S1�����v>� jCF "��նlm��i~W��|��ҔL�8^#�d5H?�q����x��}$Íh�oڷ�s�S=����î��
GwmѺ���Ȟ۟ȻNG�����i'�x���|x�����̧����p^S �;���d6�w������u�^.dY�;�-8�i;�k��t�`8E�Ԟ�n�.�������FK1t������	t��?}�%���� ��y���.eb9;�1(�"u��/%�r�0U����%OС���	��']dɷ,����4D�;PA#^	VIR����΍m~?�����s�@T�S�b03�;7��Sn%w�C@�s�-�22\U
~��j����l���A�^0�
�i�`���Ҋ�P�f�
��y�y��^#�{�XyvO�5�s�ñ\��9\���]N�EGl|<�h�@�:��o{sD�G8��/$mg>�����룔�q�K`G��O�"��	���}�¬�<��E#`ӽP����;�Q(�1�0�V+��qWAL�y/�n;�+Rw�j�������gg5�G{	�9%�=�����T��p|������z�bY*G�H�Χ&��_������� @��R�ɠx���;�Gd�=�2r�����s��D�
֏5����Z�3x��ϙ^,D�	ܑ+�ܻ?���k).u�^6��@���r������:Gp�k�Mc��0shD��P�J���<-T�q�:O�����~^K����l�?�R�e�N'�u��r/����_�~�� �h��pc�M��>[�K��EiyҖ�L(����|�ߋ�+njwOQ��H��~¹�Y@*���i�-���6a�a�i�Qf�h�{)�"7ͧ}1���K�$ϼ��tH��4��e��vDm�-}����p����b�p�W#0�2"h?0"Ƭ:q�v�*u��|,j�"�:"�@�Y�L���A%���=�?P���c��������ak^(���
i]یD�)��*��P[L�V�sP�b�U?�̉�[W��?��}KB��0�*�zĽ��d	Z�x ��,*�9��t��]Aj��%�e��i�tF6���SmD�����Ia���K!����r���B�<e~���}x<�A��P��t�e~~0�UJ6����(��#�P�^�J:���Y�b��z�Q=�?f���B�׻�o:�X	���Bu�$�p��̤}R������l��T��@��D��pe�x{�XF��B7�I���P��`;L��@Ub��R��8)p�Pzl�ۦ�a�<����U=<�#�	�I���m`���ͳ�?�j�$H�Bd�S�����F�3�6�zF8�ݑ������K�y%8Jʦݻ� :\����x�d��Sd�����|����u�^��Μ��;�`����&��g=\)�nyo�`�����M{��e@/F�L��:��H:����r[2��]w�s��?B!@�FEb]���>n,��We��`�f�op���:�,vn�R:��ۮ�a���^�O�2 3eO�p�ݩ�2$[&}���`�d���1�cw��5H����ds�i��C�5�F@��������v�1�?[��]W�)�`ӕ`�Bt�4v�BYy���� ;K��e��(��;�TnV`��f��\��K�GO��p�|Hb�0�E�]T�X]���\�T}`��p���6OY��ei��X��o��)+�<R�"�r�I�C����N`������4{��D{w�d�đ�W�����M��~lT�R�
�,�knOW|t��@�kl��v�Ư�ar@WJ����A�4-�݇(tY�X�^$8LOJ�%���������K��z�{u��r��MP\i�.��mP�V�tAa�K�[#oo�B�)�:�H����}�K8����O��͙�5u�=��s��K���q����	�#u�H��'8v\0c=��y�c�%p�P$O}�����C���y-ת^�&R%;�}�h�c�>B�m�M�(�"[[Wp��C��	�n��@��3E$�T��ŏƉ��S@B�"���S���,d��y����[�>������vkz=�{��6��-�.wP�P�"\4��a*��/�p�E��w����&*f���d�Dx�O��jy�K���R��P���D/ i|7D�{l����aIB[�����2��G��L���Cq�^�}Ĺ҆��=x�{�e9��ς.FB#?3�m=�+*�b㢥����]���,%,�\�RK��̞1(du���\p��SD`��.ʼ dZ_�\q�J�3��p���,p�+<o6��z��=�[5���ѷ�K+S�&�ց'���f 1��$%N|��s��\$]���B�%y���p)f\�R�Ai9*���9[\��k�<��.��z��;�B� PU
�����[�� �C�s��.����3�#oԖ��h��U����]�y�0�C�6�漷у#�L�IY�D��NQ��yK��9���U�z�X��Q�dk���,-��P�8A���oQ*|�@���zV��mX�|��C8���fC���y�m6�������Mbt��0ٰ�2O~��*V�qxӁ$JĬ���#��צ�b[ 	c%߿u�_D[�N�m���W�(�#�t:KhMt	r�I>p�����b�O!v�������l/@]��D[~D�íJ�����n5= N������3����_�'�+9�G�M�Z���w��7Z5\3"|���wI��n@YaOa}�'����ś��)U���V;14���Ml����v/���_JNӝc��T�©˷h26�F.t�8O��>��&��$==�{mQ�����/`Al7D�bQ���jr���98w)$X��&� �r_6�P:��'�}��]y���B�	������1C@�YI%�36Ks����{B_|�}q�0au���U"JXf���u�ƇێΧ��*f�+����+:��>��p��>.+,��v��-��t��|�^i�N&�tc`R-y:�^{��h^7�Ò��Ci���C���Z�S��-�r	:�f�&��7�����5�,N��Y����ޏ~�������>�Ƌ��殣��Sc�XSQ�x�̀3L���c,d+�}���>�u(��w��� �Jʞn�xY�?���Ħ��a=:v��m}�ŒG ����E�/�-����ՉpήOiDY���+y��9���I���)h����{֍�������g�p�U�^&˭�B��[[��e��L�P���0�����'�����{?���K�_�=��CϦ/}�}� 
p���=� �� �_��R�v^Y�5u���� ����&�a�G>@��M{�{���@+�}�#օ��8Cѫ�������� ��5���Ha8 �bQ��hћ[�Y�!��+��/�)�	�<b�ڐ��Y]X��v�W ��KB�Z(��`�!��Պ��U=���&�J���j���L��d�!+	ؑ"���;Я��/j^
z;6���d,��W�O)���yw��s��;�4�ӓ��_�J�\�fo�6
��li�?��7̮DE���EQ�3&�������-����k/( �OW,��P�B�W��<yD"[��])�;TX�^��˭ԇ]���{��x]+!��Y
}4����N��uju(,u��ڔ�����.�?7@���t�R*kU)�@�F�����-"�����,Q��V&� ��
��L&�]h���Th�)��rF1�B�&?��0 ��V��!�B>�ځ"����̋N��QC�B��oL�-�=�a�8��
ɻ�$}��8�,�5�4��.�r&6�9Vf8h�l�bD%TFÂJJ?�&Y�G!Q��T�(Ȏ�Ť ԍUfM�
�?>�+R���ƈJ��*X�'���#&�?��?OB�ls���\��o���L����2��Eu�G�)M�:F$���D"�)+����t[O.�4��ĠV�	&A$��7��}6�@�������h[����o���t�f^2H��P61�W����8��x���$:��	���B��pcۏ��ʘum�s�	t��`��֫Z�ݺ5T��ڮ�3��f��<	GU�F��K�$�d�(��#GFdcG��.�ŗ�~��P^���a�6�\Q&�5?ø�v�R
h��ٴ�����J>R���C��y��*<~H�]%�KGx�4^����ە���AɲU'��/�*� �S_���zňA��Ov4���I�,���0�8�]X�r�ڽZ���HTG<D���f��>&EG�CWP$K �3K�M�l��P<�u�k�zl���Ž|R/�[q-"���˴7�=g�5b��H�%����_�+ �ܔ0�YΫ���QT �Q\�dl�);F'� J�v����<���ܮ#�7�c=�����i�ޞv`�%qn��z���i�1%m'��	��Q_�Ub��	�&��t�W��ߧ=����p��wH�j+_̠�׭]\5q���?�p��Q	�q��HH��B�O��&y��P��,�"Do%Ot��������3���a�1!��g�%��")(r��� (K�騡5"Yx%�)�n��t:9�O�xb	�`�/������#���^��zj�g�l�D��,��Ps��[D��8:�|q�c��u�wʽ~���A���nL{�,nku����=D���X��Խ�R`�7Z���&k��gU$1��4ρ��{+�)���J����E���~����@V��46g�0�lD�<��'vq�
�#�B��%�dv�� "��u��k"��>{�{m����E(�o���QL9nob"IJ�t��/�~���nֳ!����"�L=�T2��񴤍��e����]���re{>��XI$�e8
m03�W�p��Ǣ[`��q����e����*��h�s�`ۍ�f�I�t)ϱѯ
�{df�H˭%�M�_˩�Q�x�m�z����nT�I9������f��v?��ox�I�.���{	H)//����F�P�-Rw��ҫ�����Ch�"�"M#�4�D�[��	0�R���#��)�Oj���>E���L}U�&�F���
�!g���,�NE��m��P$uk�X�N�"���-�1��õ�D�<��C��04G����Lq2)����������>�\߇�4Zc��j��Ezҋ��s��O�,lG��ذ� ��q�ό��Z��I��\B&!��$?d������m>��8�!/u��u�������6Wր0�d}�Ҙw�b�z�H���tg��5ʅ1]��8bMj ��6�F�� ��cj�F�S�Z[uW�{4�p�v:�E.հ���l�FpI��ܘ����|��^k=��W՛I��yl�/ʊ`�Q����ް���'K����3K(�l�k�9��b�umה���U��0�-5Na2C��bqDG�7Qs��?���d��ɣ���z4LɭRi�u@�fQѬ�"�>:���0�#I�	�yO8�0�������C�K�y�(V��N�����K�:�#�(����P磱�˳��4���r�g�_OI�ENJ�ư`ρ���B�'����p��qT
����[=�9�ܵ�l��͌!c�n�?�]���<��HwHN�u�k�f l	V�e�5J�'�Ŧ�ا��lJɊ$�F�	XP'X����/�,�=s1��<��}q��:�`��O��C��'�}V�	`����B�w���v2���^Y�r�{�7G7�:���.�!w�X�!&㇖�R+7V,?�l�K�T���J�M��_TfP,�Bm���8iӫ����9rX2S����G�ƜQ]�-:��n���D�
`��Z�O�h�AH0$�β9�tH���� /����V�M��95�$�뵉5кa�Z+VfWL��\`����J�w�uؙ1M�ߖ��Y6�~���+�۞M�%L�/��t+Ei��1�����*�%wC� +�"`m�������|�=�w�y蜺)F_���GJ1��"5�m���U�d�&�Z�4��Ϡm��L �`����q��#	��:g�x3��A���7�5��@?5��ֈ�ͷ�Vm ^_�%��>⚱�,"kmy���2R9a��q�����W>>�{�<��`�+4��o��.���X:�=����Xv� ��D����"�*%�����[��XS��f�f%�zI ͠��˙j�;9o1���7��T���,F$}�$��}�V(�H\��j�Tɨ<����Q���/����A��貘��*�s���8��}t��>�L��0a;�f����hj�uW���V�7�����
�0ϟ��6��:<W���4N]Z����`s6�v�O�=!���7� R+S��U�ҹ�_ʤs)$�E=�M����&?�~�xuZ� u#տc��9�]�P���g�{1#(�W�� ky7A?�K���@?���{��#��:S�.��b�y�2�	�_ex�\n��#^�Ҕ��w ����qf�����Y�d5 ��:��e	��]�=�킽��&j�a�q�S�(�9/Ƚ�Z6b��୲��M� f�t[�ؠ �w�K��qf�d�_��2�R��_�YJ��։F����	t�I<�uX��KЁ�Å�`������[�&�6����E�t��C;�ӣ���
9,3��V<j@|���M�"������C�i~��>X���~����j�&M���bf�~_��mN�5�E�O����o���2�<U�!��f/�6��V
 ��j�B׽��om��t([��O�tP�{>h۸�sFo&G�߽�E�0=�R�㉫uE�|W�ǕZ��q�$����0 ߏ�j�G�:�d����p0z���uD�>q�?��Y�ߪ ���P�	�.g!��4�$�4�<�,R���]��BJ@#j�D�(�1�4���m��#Y�n�J��_��sa�ͥ��ߒ2���ܥ�r[�q��[Nj��6˸���lz���`;�C��f����ǳ�����Qk�>s�{��K�Ι,OP�2��E� N��]�I�x�bo�eD�&L��E�Y��jn���J͈��`뗐#W��"U�h����)�g+�Jt=�*�I�ꕵ�p)�"K���:S,�g]���tؔvi��`���k͚Q��Pǚ�>;��'|W�𮯠(���Q��M�ey&�ݓH�o����eDu�l�����׉7��<WR4�M*��C�����i4s8?</��q�j�b��W:�kdp�*����f/�$�^�O��v`��d�j.h���~&�-{�2S��nS�\ʈ�j��*&��n�֜_74w-%�R���9�<G-�!N|;�)��a��d�|ޓ� ic"%�Ç�3lFZn�@�Q]��6���'R��&��J����'.�b���L��a� J ð�!ϩֆ�]Nht % ����I��{�R�GJ6c!��#��5ӳ~1_4\�U�~�QH��_t]
������J�Z��h&�1�!�e����]J�Ii������+��v�K\i�b����3g�$��ǆZ� �>��/[9��B��9l�?߶��c��[�n9�0bJ;$�_J["�I�0o�q����J���@���<D��u�$z�y��ڳ���sZIxڽI_�Ʊ�rܵ���o]����V�3X�?@��&]�[siQ�����$�5�|��UʇF�X�YY1L���p�d����o�{#���l~<%p'M�t?_�����%�� E�D���c欕[EO������?��'p�~�e830𝍪TkhW�0q[u��5sl'�)�BG�lU����j5�@=m���-ǅ����_�P��I��vWӜC�X�NG��a��f�<:X�F����Y�QijgGf�L�����>�V��������8�2�4їd�NA���ŀ v|��*y�'�cl�&{-�ص���|n���!EU��Y`}'^`��s|��΢�4�c�{6���(��Y�Cֿ�u����s��m�+��zl��v=���TYde��?q�KC'��ԏU�^b��|�T�#5Af����:ޢ���w�3Qn�.���i��c7����(6��x���ROh}�P(̃��g8�'w�n�s�(�p!4�9�l|Ve#�����8|r����<�n�|AE�����������8�Ո�7��t���f@(�n��]gG��4���
�[��Z.U�q����o#KB+�.b9�Ej,o���a��'�@B��K'���z��� '|[�{vC�,v%T�SR
b4�����%�\�ß02!R/������Q�osI��V�G#��)����Br6{�(K
u��[���*�~K�1M�j�*+4�X��ϛ%	̆�Ĩd�v�d�T��	R	��(���LGY�]Xq	����}T�Քv�=��l:g%l��e��9�	�B�e��i�����`����.� J�MGI}�����`��gH���cl������j�X	a#vM�Ә�蘳 -����m&�K
{+�_�6�81��xX���w��Hm�m��rD���1�I�-Y�c�W�`�IyM9~�,\�ل�8vV����i	=�-0�Qr��aE�eUD�����2�������1U]��V֡�]�K>�`M4H#L��8c?���\s)8 V�`���*m�$�Q5!�]����/P��z`a�y��~��mn�A�k�Ǡ6w4>��E��O	�;��H=-���"z���\۵��wGc��G�x�w����d%kY���w���bo�AC�`?�#��Mh����õ-��%*��K8F����͟2Btvm�,��f�B�����ܿߟgg˞֯Z�6.�r+5��y�Q�޷4�����42���x�@m�\�ac�B��6[��bKR��̹����oOV�o����l���<��髢��0������������:S�#����1�(�D��y��JQ��+�.���G�ғwS���>jb��g�}V���}a���$�#sdz$�fh^ܩvgPY[ⅺM�ݼR�� C^�$�S6
dhj-���=�*����1<�Î�c�%���JnI ?�ԁ�������vgᗗ�@�'1�#�fM��a&���9IB��*�q� )�������
���p-�H)lu�O.�ٖ1�X��s-̤]h�9��v�m��Bf����ɹ�=��@&]WG)Th��D�i����:�U�bc�b�>]����W��Q���Q�w��i߲u�����Y[(�O�Ъ����P���դ�����G2���K���:��2�T�v�`��2��_]R1���ᡰZ�	�0���wY�=/xL��AX-��4��ҙ�X.0ڈ} ���}�T����UvW(��)4K&�����0����[w3G��.���2l����Z�r#���-�8��pr��L�(�ޥ]��fZ5yxug�C�2�j3�;Ƅ�x�p\ Gm��;���X\�q���&�+c�z#��Q��L�1�֠�b=$Y�_��IB����P�N*�F��Z������c|������~����w�~�m[F�f����V�vY��	hk_^�h4�h3`?�������g�!1�ْ�R�dt�-j�Ϸ�r�d2T(��dqp��=��8t(�9B����͆�㋞� i{	0�M��|���gP�W�h��Yy
����50'f��/�gњ~�I�z�t�����t��W]�!��<�&����u�x.lY�;�������9�@)�^�!$'�����a><}�~�b5�B�W�������	�=���r=>=9&�T�K�B~���̌t��!����\����w���7 R^s�!�L �;)�Sf��)Tn�Nݲ�!��HG�Ѡ�H����������qUvl5���_�*LZ�Z�黧���ݰcbՑ_�c:�i[u���g�du��O>v6�����5�oZ5]ֻj�Z��0��'U�%�q�g�> 5����>����6�`��d��F�I\�.��3��Ew��0:�p1�\������z�ӡ8~'��A�����箉L�1E�O�7����k:?	�tqJ��W>5o�����Xra<EMGe��Q��KS����S�T�~���ΛԱD��!~�����*�����e��Di���͢�Z�e�Gc��4�{��Z/^T\��K4v����(�i�/MڊE�����	#�hz,^S6ޭ�v����JN�Ǎ�?8T�Ӓ|�݆���A�2�A��40�E^�b�t�}S�s�+ެ9��c�MC��TU�4w���-G�t�-^�:��	��M��L�\a�w�)T��G��\����.{��1f�ծj�N���+��m%XϯсAܿ���/�пGf�Wl;������XiRƥT�Sbd��YS2��V�)(o�����]�������_.���@��^��3逧��Sn��7����	��0�l*-�Q4��VmE��&�ؘ$y8-`x��c��5W�� �
:��Qq�4J:�+�ɱ��p��C:���'PD'�G�{��R�20����@���d����l�F�b��N���J/m���5��x���P]�4vJ��v;�Z駂e���?�s�����'��q�9�|s�d����}iڿ�S���V�0�b���YB�����@=�5
�-�a��|��A�VUN��ڄd.|��d�������֢v��z�Y��rV��m`R�mP��vQ.��b	����e�^^?ʹ#��1�q�.�a����h�<�zE�1O����RVǟ�]��P�}4
�DqА��,L��3�y���$��B�a�+3��8�����Ϊ)w�G�}˴�xvlQ}��Սm����f��|^�+��5+N"=�4}��Ӣ�RE[��|���$�ee>Q|<[��������l�ް��Y�!?�|C�l&,�Ѯk�(�x������.Gj|!=�F���֢h]����)Ŷ� ����z�ڼ
%�h��1�CK��`��c;���l��xh��.��vW;��c�b��l'��P�ΐ��/lm7p ��x0�f��8�%eK؇�6��@X^�
��&��-A��RV0��pee:��e�N_������N�Y?�$>}pNxd���`��j�&�����cٓ��v�]J�>)m�C���{$o�O^3�DŚ�0��?�ATE�a��#�VFk+$��~;��[���OP�y��Z������?��m����������d1��\"�^�(P�G�Tu����)!�([�Hб������R��Bִ��뎫�T�%��B��C�Q;8�HA�9�j�f�]�p�~���|�r� б�̔�X�!\�S{�K��e��|M�eЩ&PA]OMxV�xCɽ����<}��2ek E�Xg�&���an�K%U�Vޜ.��(�Lq�$�b����&6�X��7y]c9��X�Va��Rkw(B� �
W����{v�U�킧�e�e���[��|&N���	��q1��q^Ӷ��Q9Lr`����T:Xgxrƹ�/�|�X��{��}�~����*�rc{'������sf�g͈���(���撩>�!7�����^����Rg�2��I&?�Qi�w^�س#�+G�I������mD���3.o��SL�y5~�Q%�*�&|>Ee��e�CO0��.�M�ݖ�*���$/���hC��X�Ay7�t>+�)9d"�( !^H��f��ATb�Y50�����������(�o���4pr���|�#�e�p'jSt�n\0x �#�ٱ�@��t�lT�f�e>��_�����)�w�Kf�� _ڒX7GT��`���a6J×��X��mC68P��\9E���s3��k3�������Q�����^���E�io�S�C���c5'r��:yyS�"�\`�� ��.},���&������Ҝ��*��렪a��ѫ���0�P��_#��V��+�bt���e�e!���N1��dzړ_2�����c�V�7�B*�c���aM�7l0l����$�,<>�;Z2CW��Dxq_!ñ��P��ڣ��B�؂���n�hc�����l�����m���ڏU\�A].��)�i`6���2���D�d�]���
<�ݡ��D|	��DFz)=���7j
�]�D�׹݀9J�UPc�Lg�a,}rBH�ӕ lR�"WGϬ�)_��P����qO��*�����"�؛��m4g�v�a�d��F�
��W�m�x�2��	�WZP���F 3�p�E�V� ��?@\(��Y��JNߧu�1�:�9��"J�Ȋ�"d��Z�++���!?�tF�F�&�t3�+]��9���:r9@�nլ&O��}��ؑ�X����A���Fwyj�	����q�-<$P}��[�x����*i�'�G,6��#i+�g2�d*?:"�ݹ�UӅq�Ǭqv�Ĥ�k�E8p��V��K2�����.2-q��>E�Ib761I�M���KN
]+S!=T���Q�j*,�]�e��y���hMo]��X�G1qP.@�@� �)�`K"�1�6�NOՏcNۡ�������Y���U��W��F��.wr�/9�|�u�42���!�ɞZ��X,+�K]]:����o��H/�$._��M�>KЇ��u���ءZ���A�;˷ ���c��P�k= b�j�q��1��|���)"��Q�?�#ɖ�]ž�Fڰ��"��S
�%�5-��ķp��-8mV'��P3d��oh#��<�m�M@�:�����͵)B������ot�}�ci���>j�ǰ"O\gRQQ-��������F����C�7���M8��4A1)�w�$]����;�W'���պ�9߉�V/mӮ��% FP��r��RL��D�]�憥�?N���)���T�a�euX5`9D�CP��"�â�H��X#ܠ�;�l@���oI��}�e�.��4)�b0�� �4󊸔i��6
QYs36���{����Ն뺆�6Z�ԘRlƻS�������7��ߋ+�.�����ӥr�����E&�gt �2S��fl�pF@�	�[����Oٲ^��R���c�l�`�$Θ��lZ}:����u�nkr���UzP��d0�J�d����>�yH�]��˸J��"o�7���T S��g�%���妕5�h��
G,!vj�sB���K7��[��A��8`	M�'C;Sx�w�^yy] 7d���e>K��U��	��G��W��Z녓��R�����nvW͔�Tdj�6{[#�gyQ��l���1I��AC+b�z�����֓��Hdw����1N��t�EPt��nU<��Ar�n
f&��KÂ�a;UDCB,\��l9
���S�'ڳ�k�РWDg��0 �����8"	����45a�
C�j��Wu�S���6f@�j�FZȬ�鰎q;�0%�?Hݜej�=V�y���X	��j������T��x�ɐ��/�ZG���ᬁP�/�clBN�D��M��E�����ճ@ѯ�0qT����Y��'��]�0�w�� �k�)Qȵ�g���g�h,�����-Q�!I��tU&��R�2���{$��Ek'�P�1�{r��i�7(+��:�aw\ol�\��S�2h�sp�����b>Tg��M��St�Ѳ�*&����brE�7D4�t��D%ys���],���H�)B�M=��h&�A١�b��3�nip>��fzUDT���-x�/���+o�*_������#�X8�F��cE6��u���������uA�=�*�=�O�����t�*;�+p��$�$1�G��������i�i�����ܛ
Z�Ղs�|s��t]":L�]��B��W5�!�!9�ro�ο��������E1�
�9���]�Eü�6H#���?��Fw�Ƅ�e�&Id,�����
R
�ad�ԑ�z��X�L��N�<�J|��!)�=�$/�js���e�[c����� �hL��Mc/�{b�7�0��=�%Q��P�!�bʦ�x��Q�nߜ��:/��|�X9!Մp�S��M,����G@��znI�{��t�O&F^w^�]�ѱx`O_}̮~�Jק(o]}����k�b1���`9��:�q5�Ґ;d6���nwp%���ܕ=�kf:��=&"���]4=!���Vߜ��r�p��F����[���pT)��M�6I��@��1���ʦ1�s=E�b��`�T0�]��[g��*��3O>187'�ɖT[o��M4WY)G���F���K��״�iG���]�l[��9�]�K������%��`I��@�E��Ē���͊׵���8N5v�<�>{�����n�~B�;��ŃTkq����lQ�E���S��gs"L���$�t��:o��X$��7�8:�
���u��������|pG�`o���� 35e�]��"i��.ʹ� ��w�A���T�B�L�#5 >�{>�pR2'���,�̓�]1�2
ÿ�c!U9��.Yl��0��{���`A@�޾@_�=F��eC�~���bp7�aP�����)�9��3���Q�h�V/B$�P���c��.���w[�#D��!43uePn��Y����+����G\�-��� ��e�j�G+�'�d<�J �'hC�������V��o���e 1��}Q��(u!$ ;w�We��iA�Trm	[t�*4��h��������������H��=�Ä_��BK(�Cx��>�OJ-|$=�D���UL%Z;����+���^�d�h���QT�uk���-��KJj<�E�J���G��n-��M*-�:��o��G��Z�oEkA��
�@��N&��Xj��Q|׻�b���Dr��>�>�NG�Jm�e$������<�>a�^�G�il��={M�K��<��@�vd��Aͥ��h�~�)(��X=�%��4\�����ԕ��*: ��W߀f᭭�1&�ê]��~���,+�3N�19_LI��HɐG
z�Nv��o΄3[���F%���E��w�5�߷�N��r��4rJ[��S����Ԃ9�4%��o�~�������`�f�(�X�[�JW�w?�05XK!��y�$�4J߲�[��.�����me��eč�k��'-�B߃u�˘X�a���&����i��[��	���;%���5��aeX���L/d�{M���6p�le�� �D	���Xf/5\yn�RM�> A�(���~�ĺ���0�A;1�+?kxe�,j�n�C�?�Q�mEp�[iD6
ݿ��=�W�M�;l�_$&�Q�^�#t����TK��f�d�HA��� f�Z�����H�А?Mg��E,q���z	1B��{��Bv|z-���811��3�h"��	�)Iـ;��c-&�u}��L_{����h�w��zv@p�t�Y�|��n�yi�a�k��I���λ��i]߅��ÝkҦQ���Ɩ�SS�f���
�%:>��٠��*���F��z���vX��On��	 �M�V,�� �)�D�{�'��i�n7o�;���Y��W��I]0fQ3dL� ��`=Xࠎ�����2l��t�3���V�u:I��S�����oB4iǽj�
|Y/IXf*��Wq�{�z���?N��[�JR�u0y�mT]}N�~w�AJ�U�M�]=�N���]�)2`�<�� ��k��J��Ӷ�i��e��)"�,� �K0T92���\9_�@���&�lޟ]p5-¨�̜x��l��UO-#ܭ�sB�1�S0�ғ��G1*4\�?1OиRUgZ���������W��j�7Lh��^Q\3���Cҋx���b�W%��(��~Tnk����0���@ �N���S�&�H��Fn�m�a5Ɣ�.�k6݁��w���%1�,����Ǡ���
�R�qU�F�9�]uD�bS�m ����}��������5�`�6I�j���{�=�C��@�.����?�����}ڨ�h��S��Z�}�f��Wz�g���_${��K�o[y	����dL8Cx"AY���q$4�*{N����9�JRxsr�D>¦�!�Q��M0����\����JLu��M��ca�ĉ� -�Mh�۱c괫t�[���K��`�2_?�`��'d[�T_/+�TYX��ц��!��=�&�����z^���:D|�����iľ������e">�]k$~��;��� 8�!=8H��]�]��W�˱o�֋�(��[�+�xg�$�1�/����%������
�0��׭o�\���l�H4����f�C��1}��UR��3������Bc�d��+#�Rc�����e�ܸ��uȃAη��٘{���%l�9뇵w'; �+.�n��6�%#��s C�4*�5-�&��E���30s�6牚��&�E`A��q������#A-3g��\����0�{���g���\�Z!��v⻸���L��`��n�7�RR�f6�je���̄~a��]K���N�Ce:/
v�"i�oi�h=��|�f�f-���߃\�]��:�lԉV�W�l���NK!�nK<��)a�$����c��z��1�5y���P�nX3�M>�#A�&�O��ôl{��Dj���g�-��?72* u���1��y�:�y۱�|���M-S^��Wcq]�3VI9c�ɩ��wf�y�0Wl�Ya�#���#4������D�jX%���zYY�6L����y�B��>��^Վͦ�������/x?��r� �Gހ����ݴg��*�_z���@Z�Lk3���\�	.�<+R0�6+*өPr"�NghA�t>�h�T.�]��_I�ČW�)H
n���l	)��顄��Y�<���UR2�E�n.�`U�gԳ�D���j���t"vp7�(�?���g���p��e����_�9�1O�%(�v� a�"��Jl��Y(�%��-\�����ظ�JՙB#��v��v��|Rv։�7@wz�I�=��*����'\d���IS��W���S�R]jh+���~IR�Ʈ��@�6��W(Ƒn�S|j�\o*�Q���Rj����P)_��?8{𦱁���A�.��#�.����E�v4�cj/�<ȏ脇�F��	��6�����#n��9�S^7Konu�XS�������u^��"�l
��gQ�W�BH������D��c���+є��)�_���G���'�ٱ^߳���md�Ms��8Sa���-�m���_�A���}d��L���,�j����304�Cb�3\���h�����C�s�b��l_*�m=�V&�����P(�sT�K�?A`D	�ݎ㾙}�N�DI��Q�0D�/��cv=��!�ݞ��M����꿉�P�fOHR0v9i�.�b`Y����������v�n��?���XU�>�0�Us�{a4FT�����۽¢�O ���)~�vp٤k[r=�wsĆU$nÕ��ߪ�}A�Q��f
.�r����p&�r��0G�u��\L�S#�����\!E+,����*wK:4��1�,���B�$D�gjR�B��'�o.N�~�v9�S	]BS�X��'�\s�}��/��c�C���x�)���/��_L5� xDX |2��O��NE�(����H�iQ6��eϧPfπ;��ؿ���;�]���/C9�y�;%p���1	���������]c)ԩM�B��M�a��(����E;�Qf���|�k���EDs��4= 	;p�ۥ��.�`�`HN����C��Ij�[~:��f�(W)�[�)��N���b�d�	�J:z�1���5�����N Z��`� ���t/P��wa�7\H��lM-r����i{B^/r}[���u$ �����8|=;����5Ej�-,
}��IqMXa�@��U��FX�E�"�T�mp��9@B҄?"�x�����&S��L���������Cxn��m���*�|�?�f��g��]�!����M�aNd��V��]H�]D2A�Z��q��]G[�m�9�-�"�cz��ЛS%N��mq5�4�GC��H���iV$��?��}_����w��.�Zidt�>�6sK�jk(�ޠ�n(�µ�Y�NU26l��B��yg3��ij"c2߉ܠ�($  = ��),��N�-�\o������;��a'�W�-����eu���+�e��_��r�tp)�J�����i�SYuW��iR�1��NK��߁���B�~������I��$�y��^��hٟ��Ѕ7����I��˭��5:���o�����9�vm���ڋ9���^��|�����S��E0 �yPtPCH��D�N�uɬ�	;r��}�9Җ�������:�x�I����UK���ݛm� r��Í��27����'.y�\̮�T����;�y��#4T.s��/��ح_�^-�Bz��YC���LY^J���-L�0�/_c��m�jU��M����*�`��jĩ.u�w���8i���&�I�%����!��b����߇���r�Iլs@��U|����8R�c@�R��G�NL-p�ݬ1➸>��s����eh=`�B�N��VoU,.��0A1	�,���f?rr��A2��+�-��h��w��@H����o�P���(�$���d��Sߤ�@�%n�1�����3��쎞���2�.�j렺M,� �s,�ex)A�Yt=����29�z�7��а@�_���c�(.�m&�����/}��:	q��\������O�ÓE���9i����e�d����x�Q�v%��l����V�6D�4��P~�ʶ�N�B>�&�Ν��5¿���P��=���Tm�*� jW	Cd�PX`i�������MH53E��8�tP򠘏V=�@!I=���[�������C߱�c��������5���8�qӜS�,���"Ӗ���,ݾ�
��d�o�KF���p � ��qP{^��B�{��Wn�֏��.���D�5̉����Oe;?��<��pm�̗�վ�w�U�3����٠�L��t�E��)��1y�����Z���~�]8��ض�@�cEq����N�B(�N"�c(B��H�
&P1���n��o��k~�h\6�
��,�����S����=G�X�5%���y�@���&���g� ��;[��c3{��/9���|> ��O�=�&}5K�����zN�o#VS��R*j�#��kC܄T"��[ʵU����ft��|h�&!X�6�~�����nT�eH�&a޸�jr�U{�1m� U���^��������K�H��X�/F�hB#Oy.J�\�J�\Y
�;[n��+k;K2�X7@[��Z�c{s��_|%#�[���j���Ү�Gi��6,��XC,:	�G��3�g=p�7 s�HҮ���Y�� �pҫ�Y�x����- ��۸�s���Xi6�W~6����:�Q>U��l=�JȖζq���̤��x&V�t���
aA�Ah�o��ֻX�2��i+&}_I"��)=������g��+45M"B1r��(��U�f� �(*�]����}L���-�2�|��^)7I��y����-1KHϛܗq�$9�~�/6`�(��������._���^��P��2�Iָ���Inr��ۓ�$b^\�,�L��m�-�Mu�T���+��֤��S����4�Y��'2�=�`Z4A�i�H�?-qpo�h?;p@RC��aѼ��Ϣj��9�+z�IU
��d���(m�����]{Wr�ֺ�!jJ+���j���p����I^Ս�m���L�����x,=Cy%����]��P���шG��!
~�bե�V^��渿�	�{)нp��D(/v���)���f#Iރ%���5�x�ĝ^�C�\��N�켮�y����&���y+�]:�D��	k(��C+���Q�D3(..�F�	vE�[������C�4���J�Q�W|��b��5�u������ÕP����ӱ(��wȏIV��֓^�-I�M����:i��.̲^�p�$=�J0b�Ć�n9�r+H�0�|}MC�f���{^��{�b��SB�喈jא#�.Az�K���6T~O�f����Ƌ'��,쬽���Le��N	�?��
�a�w����P��,F�Ρ昏���V	�m#"T��I��.��6�L��1�Q�u_�!w��B���s��T6acSq�
�l{;'��|�{��J�(e���h=mB�����1�LT�zɮ���%P��̎׏������u�����K0Z�y��IS�bk�H6!B/���K�L���+��Կ[��e�Vd�'��\:����		��@��˜H�2)�؅��YD��B_(����Ӛ��˭����}��!s����#�9�u�(�0��<D<����P�JgI~AEyh��dt��NW��V �v���*G�����3W��R�[n:��)yI&C@k��j���a�%[ЋB�����v�T"�_�{��H�ȑ%l�j��8.��&��M��,l_9i��?F?���k[��_|=i1�	T�tuh��#��D뀺��,41x�~�~�&�8J�ƕ|��5�
yns:��?�E`��n$��B�"�_�6��cT���B;�̲��5w�e�l,��h�|/3�^!d����&��l��'C^
I7���+N��7�~�#@������tu~=�a��_8�mmo<\����� L�\�<	��5fV�B������&I�\���4D�η���Tc�񓷇����b�t}jHSˆ��,�����p����-e�WN������'d֌M�#q�� ��G�mwq����2"�UX��F�H�����S�I2�6;�jd�(|R�47����#�M�8eC��o(��T��`N�qԯ,6{�g�;y��ds�RP!9�O�Z��2K�j��91~?��;�^��r��u��VEt�[�����ݪ��/gf3�$I��]b �8������cIF�/��oIA���b��k�d3�ԝ{R2��׌7e��RoeM&��\8[�~��j�1Vz5$�*,;�A��7tB�yPhc�.5����
��k��d☪E��:��4�1��8 ����9b�T�?�Ia��6.��bEyw�t��J����$����
���9j���4f��!7X�A�n�j<1��A$g3�0�K���Y;� M�pZ��xs�ػf.�N�m��{���0~���،U��J��0oY~kZ�TZj�W��+�a�V-��������g�+KdL�r��p��^lR�$� �Å�؏	8��͈������T
����gs���V
Ha#a���9��_�c���X>+Xj�U�|�L2��V� +�¬������P|-�3jq.���U�s�5W?�`���Jk�3p��k8F�w�<1��?Z[�������\v��=-��	oV� �E�N3�����δ: �޶e�$%|��������C��
f�6}���q�Q�������z��\���{t�;�����H��;���{�xqȤ*��Jh�ٕǚJ~j[/�����Cq[F��|�t�%۟���a$���C�\%�>mך2E����~��p��ao���$m!Y�H�5w���س�-oL�2ă�kn��+��g�`B���v"[ւ��?|�/��kёrv��ӟ`�T�!��C�����b�0�<���S�����uH|`mp�_�뫶��G�F�"�>���a�����g���n]b�cWF �1O���lKz�[��U�l���]Kȼ~d�
S�T���+r
��;���K)�ɼ177U�ܓ����s��l^�����L�40f���`����_��;������q��-q�1���Lc��K��F���i"�F�ٗ�E+Q�k��yݜ��y���p'&�;�@�$
�#1"jgɴ�d��3���b�>x�&6�	�9�
	�� zsƫdI����Kv��D:�j�:0�&m�7�S�8�KE�NQQ@��Xٲ��Շ��~�Z�R��#�\��lwD|���LE%���������p�{]^�V0]v�u��
�W���,I*�+SX���(�V~.�:~fC���A��tE[���:2�D�z�+{�bg��f]LmH��i.W�|�î��p���I��V�'�̛޽1�F�g%|ݥw����'&��tзndش��o�o,�f �9OF��K=���,DL�ͅ��eLfD��Y��$w_ H	�� tuJ'K'Hp!P�bN�V4��㥃h�5�щ���-T4m�3�u�J�ؕ����jD�w���V�����r�ߑ9<QT��;�I��\<Pnk�&l�*c�F��uS���&�-��Q%�:��oCർb��,��vˬX���<�9͗;�&O����5A�\e]?�u�oU3�.FndЛ���j�f��zw?8[1yf��K�"aރ[�sL�LLj�q�3٠��-X�W�;�R$4�&�~��b)B�l�@e��9n��YYS�d�(6���͟-��@�Cv@�����4�4�Ǣ��}?�������	;��Jn�&��8 �:���ٛ��XHB���mQ��{��S��mo�V��x�����r4䝏̭����~!�Y�.6�"�IM���`��E!�A�)a}����★C4�7��bs��"� 0T�x��̈=,�N�}�\ֆ�0e�;̻��;$�\G.�.=^��o�R�u���KG!��I�?����wU��>��	�b>q�݅`���V�����I�E�������L{�D�=�d�|VF�T�2,�ܳ2�/�]G��EՈ�8	������� ����59�L�޻���MbC�*�˙E#	L(�q�a
,�X6��fy�6 ~H۬�\T����K$�kE�,���1�����P���ݳ��ѩ`{��j���7�p.�t
;_���:T�+"�D�푎\�E��zod*��f���o��ǵe#qV ��á��@ ��ܿ@��f�8fO��|_M���J�H���&��K9HI�c&�˽�������}��K�4	��1�`��?UI=N
��Y"���P/�>3C8(�^��A,��$s,Ƶ�}߲Sx����V���ӝ�B�|��ȕ̙���Ͱq�"���&:+��RO�C�"�u".(l�|lW�����/�u�V��ǝ��s	����]1練��^V�7u ��"p`
Lۧ�֜�_�ө۰�Tx�-C�c{Μc=+�粑ͤ|���#��`�?Gbn{�U�c|	�q˲7k{�HZ���J9��`�����	�����(a~F�~op�0�\�Zy��v|fH�^��� ȒB��=�Vx��Ƨ�$����j�/��i������n� O]�O�ȵ����1d't�pҁ���A�[�F�ubzy��_���@鶛�i.�.h���jt���|\�!�N�U�[�;��4%5t6<�p�0���m��*�d���
�t�K�[�0�L4���g��5xz��+�ct��mp���7A����ʉH����6����흰����|K��F��Y�'~���E��^ӹ@�B"�y�a��	��*�t�������F��f����M<��x9�dU@���"T۪��� ����f���7(LR!����P'�ȁ��Q�HTJ��9!W%�y������	:� �>�8T�"�Z6�;��(Ҕ��Q�J@df�:;���Z櫈�]��ܽ�9@1w&���}]�<}7�+�2���1Nt��hٍh�D�k6*}v B�5��U�9�jN����ף�-y�U�ǿ)�����Σ�M�_b�#����C4M�(Y��3��JV���[�d���O�����'�<�=�K��Q^o�~mjﹸ��1B�5"�>#�(��z���������/7�x��.䖲j����8��@WH5I�iK3�薵�t��E��t����SwP�3�a�3����잪�
���/I�%z����w�~�_g������շ�q�|IzL�a�,���ߓ���N��~����{9�뵌3����3\=@%�:���e�=G
J��^����C�`�����@�fm�zV
��4���o�����mn)���A���m�:҄ڧC&0���?@֫J����G���`�p���_ߣ,��$�t6����0�ƙ[4|P ��V\�@�|�����X+B-�ӕZnM��i�e�Sg<ȯ�T�ρ�!�S����T��.�¡��q���̻����!�y��>�@�-ܬ|�q'�4��ϧ�G���^-Ǧ{��1O_?~8�m�8/|��^�	{; ��3{H�H�\褈�V�+�d!��!�G���7��f��ֆH��J�;�h�4��j[�sW�{0���o�|��6��B���q/�l)h�Y+k�'loDڰ����=�P��s����д^&a'�o-��Od!��}}S�σ�O�bk\��Y���]�8_~Pj����q������`ݼ�U�a�,T'��(g�1ӣ6C�g!�g�0��<^
E\�d�^���,��fo�TN��m�O�0��fR:���"E*�,Qp��P;�AzB����u#a)�LH�+N�W+�P���]���2��H
+���֫(�
�.<�h9}������S���mV�=؍�\�L1�� ���#L N���HT�;�P�V�3R�@��}��x�=����蘤�]�a�PZ�q��8/MGZ�g��+ya!�O�ee-,*Vg�����
�Ν��fg��<֩˒�:6ߩ^���?;�"��G�%#H�ҏ�U���f�#��3�$S?��S�av�]#֏Q5���ěM"-E@�1g�j��y���-xg�} ��ؤyݾ��t1̋8��M|������~�9��Z�b���ֵ/�[0�2��?����u��[��p�{O��{{�?B�ܽB�/��㨊0���\zO�������;���J��nW�ugy1�a~����Az5��S$yЩ3��p�<ߣ��}?e�����v^�r�V�)�bZ���pAijȓe�	��<e�� w�P^މˤ�ɾنd/}O<	�*�!�<P�S�ί��Ն��4(Y�[��e#���k������cb'g�e�M��PC{h���0��7���?����vz<�vOz�_���k8> �L�j�����!py�GmC-H��Nu��A�������d\Fd�)��1����)�w�cE�IĚ�l�0�	|�[�XvFg��Ph����p��|�yo���,��������^��n�7�e|0ӳ���_�-t�~�_}��B{�7�}��Y_�������k��\>�����s��&��c-�ޓ�}U�����=��� s�����ػu@�I����p8��5�V�܎C�`��&h4���%*,�u+#�J�.!��l���.��q����`'�M
�bMC�iP�W��<�B�O���|X�KeZ�=���U��t�.d��R@�n��lmK�;h+�4�T8���������"���o0=�+�dh��!��̆�	�y�-lL��F���4v�s����OV��9M_�������Ó[��Y?���@G��*�E48q\����hՀ�:%rX\����>p���")#�X�D�+�b\;�L�u@6ܜ�OR��C 0����Ä��+�t>�"�c�.��%Y#�] ��R����5^������?qj�ל��H�Lᤔ+� W���ƨҬc�dŔ����?���$��]��G��׹1�V�Sò���>�-܏�j���7tƈ:z�m`����b~0ڡ�▨�B%{�`_�E`-��@鿿�4V
�DIb��� �Iv�st`�����,W_���x�wfۀ�CRq�2}Ƹ�(�ʎ��}c��{����Y��kJ�zy���!A~�;AcSGTC>�)�3��?��jm`� V��}}��C����WF�O��tS���`����`7U_i����Iyg�����L�����p�|,�+�v���G]���R3z
6�;f��^��b�j����&o���!�(yeߦ���A*��[9�1�/µU�/�M��RԤ�ٹO��V?X~���*�]���d�w��`m���p�&�0��AB�~0���j�V���"�8��E���S0
��<; ʼk�((ᅮ�@�[��<�}ԋ��6�g��%��>��yU�Հ'��ٻd�+w���f��ok��I$�@��P=D^Z?��гt&�U\����sf��6�t+]��0[*2���ma�k�"6|�^1�4�l���k�A�e�æ���#+fT���J����&�Y$jΔL��#kۉ;�=~����<�8F��1[���J�R�a�}���}��Ŝ�kޤ��]l���&���c�����`��OZ��m�3���������6�ڻƧ�c���%	�@a��
u$������i��_Cs\k�T���(d�V��#�#�;R*�:�*�#��j���.��߰y�#��F�Fo��
�H:2ݦ�d���m�h�c����@c���?�g\�����-��0�{�E�4�F�x;�&��5�Jp�#�u~�Vl�$YН��9Q�4����.ŭf�C�ϱ%o����L!���A���,�ث�Q��)>|��TNy��jų���{�+IJ�}��羄i�>0`3�E�7/��Ny;:1`����D�$�`��~�E�E? �������ewA@t?Ģ��f��H��%��.Y�%�jZ=VH�?��G�%�k��#3o��6�p�'�\l�Y	O;3�n��(6՜�$�+Z���/�,��zEwysN�j�q@Dt(ˬ�*Id�;����t�5��4���}�Q�j�N�A��=33qB��v��F���ڂq6��*$��Ό���sYϬ��J�P�X�}������>����\4��y��-���1�L%0h�M!3���' �eF �~�ASg*�MjU��S�,lDMv��Չ��j�%ח4�E�@*��1z��~��_:�i��/�-�b7��:s��gk&}g�2�&��6F҈��c��?��	^�[P�1������rW�}`m��{�,:����8�EP_��m�Ao�aZ����ϻ]}7
Y�0���]�i�0�����J��	�^�q8�����~畨��n��.GU��`#����9SD[�ʑr2d�/v��E$Ve&,K�?V�Y���q	^x.�̮�;S�<�'z�r�F-����n�b�=�"�?&2{�|i)w�a�h�@�z������꫋�:��дk:a��0y��c����@�Ei7"U�E��Bf���_߭%\ф?����t�ɋ'G�i	~תH>c�b0`ݮ�3dוk}�	�l�|?4��Gy�7+.���b.����3�?^�~�&�9�JF-�^/�/�J˶PfUȮ�_,��'�p��)ͱ�ٽ��FV �T@�>j��蛍m��)X�:�t��x�;�P������ȶ�|s�}�2��q�0�r8���5��1�Z�(�B�0R���Rv�ĕ��ځ��l���w�ay'8���%�iG�)��`�M��;�/D,��0�jE�X/e*�/F�H��P�$���U��H�0���������k/��M�(.��9�pҠ���<�)��v���.�qQWlS2�K_�VӅ�9vߓ�LC������R��tNB���x��~��I�r�#��p����E=Y�o�N�t爭a�Cb�#�Jݾ�ǀ)8�tx&�B�֙0����i޹�4�:q���{M>�[mqU��U͢m�n �#[F�%s)S�[��y���j�vv�$b�N�w��O��
K2��#��u��?����z����C�Y�.8�F��O0<�"j�GNVV��̈́�B�B���Q΅V�yH�����5"C!>�Xɻ�G� �h�i.�̌�N��jAT��jv������d['�>���o���/G��B��Monf�G�̻К�;d?0mv�׌��a$�vh�׏� �a>M��1o�ojfܑ��O��E��Z�ġ��u쑷:�a�ia����}��vc���P(�9>&f�Η���;����>DN�?��hg�v�2��$S�9;�V%�{4����-L��]�wZ�I��Ah�Pv��C�W�
а�=(g�3��o��Y��W!U}�[B�҅W�O�4ٌ�~jA��5��@�a��9"H�/�*V�o�����\9J
��w�<o�w9��/{$��N�0����ӧZ]O|�I6A��`Ď|~b
 јd���H��w�Ԥ�|&锗�=5���Jv y���t�@����.Ĳ!�Q�����(��E8Gܡ�l������}�v��m;D�x2_5��fR˪"]˛oK�E�	L	�X2YNbDk�?	&3<����n��
"�Ʋd�bI��7�@3���t$��J�֊L�6F����<��P������mV�"~�Bjh_���b�o�씤C�g�w��ӀƌS=�9χ���g*]D�dL%�S������}l����oi�54�+���vn4o��cA.���~��3h�*�ekCm�Zsm�fA	���+.)^��bo#,nX�"���ҝE�NEze"S��]��
�a������\�>%���NÕ?��.i,��w���zy���^�$��JzB-9��ġ��H(Z�0�����\�'��zw�;�^�/0D�ԕ{���&Mժ���e��
�0������	�r[����P��I=�e:{"-�3�0Em��\�D�pv�)�]�q(�׃Ή��Qē"�Xt�F7�X;90��[�Y��m{�O�ݐz��~�+���l']�|*�eh�~�K*��Fd�\I�<�8���AA���o�lA��߰���Z�6*�V�-��ǀ��U#�!�2p��Lö��auA�`�7�d)���Xq��O,���nՃ���0��],<�x��2^��j��[3�B��f����O�N5��;�pxp�	 ;�Q���#�D-8��( �'1	��d?�JJ�����/��K�%��hk��kV�w��za��6ef���3dW+É%�
u����g��a��Hw��#V&*rk��MF3�U,v�ks@Qm��^�m�6Հ��<����ܝ����_Ԟ@HSua�7��!��ruB���Zf�p_��i!(�a"��eL���i�t$n_�A�w��1�T�,哟4^~9����p��v�{�����Tc�"���N�z��~�QZEH����uL���M�b����FN;H���s���9U7�E��7F L]�|��&[��\#�tĤ�Z��S��d�����O4��v��+Q� ��#G!��&��"z!��,/[�zl���U��%Ѧ��;�%��
��E!��J3F��I �ǀ]��ѷ������d��fؗCPĵ�7$���D>)���y)�/�W�����$&�C&a��6��9�F�U,(��Ww����qtd��y�\Y>	�f�"�at�7��7�g��9�D1(ͥy�psj�������w��l旆ಠ�h.��	�P�Ko�,�&�Vi�<���M�m�ڢ�����R$%ǾxU��Ivsܰ
�s7���u5�,��i��ah=�$�Km���i}���J�؄5���_��ڤ����PP�鷖R������T������k-9�h_Lp��롷@\UT���6,��O���Wi��V�u�g��=*��[k�m���Nh��9�2�0X���W��ba�Z;6����5���D��KJ��2�|��.���ll���3���.d�װ�э�2~���b%܀s<FK@s贖��_ߨb&�X�J�_������3mG�����B�R����]ڙfn�"���N� �\c��Π#�`1�`!�5ܘ2;F��C!�-P�u{A+���L4�����Q��.��A�;��%���u���7����֫�,yb����o�Nf�\�4��"�^�Cj�߲W�8����;��=�`�$e���eAo)i�p�ƐFY� (����k�I�vA�2�qUv``������e20eD���L���4��G^�$T�����JRl���QR�rg|Ѯ�#�/��O�{�,PO��u�"�x��un��Pkm��C���Ғj�]��
�^�O!-��%H����_p���ӬV.�L�)Z1\ҁ�x�=\*�7���MJ�%�۫��Ώ�gU�c�	o3�
��M�zX��5S��8Y��(5�:���%���Q���l�c2�U�3�9�hҹ��[��?\��1�&~�r>�t#�I�ˎ��N8��,�nɪ{�Dq�j)���?.�qH)l���wr'W�ն5�7�H�=T�GG�	��nރZ�'���9��%�3������e��tLzx��U��XTЛ�GvMG&:~�+`r��p#�\5����5
JuAmj�H�WݸF���t�����a�36ƻ}�~y���=d`�t�I%�'|"5�'�1f��9e�e��0m��^��h#��>u��}}ȢCF���*�V�(���:x��C~H�v1���A%ǌ6J�[9\,��J�M��#��C���q�!�R�NӘ�p�K>�.�{��/߳=#��c�Y��O�4R@B�9��~zj��R��'V�Ќ�_}j-��pAL�T�b����@,�R�@h���wÄB��ziC�V�{�:g ᤩmyC7���p��a�\�Dڮ�+��᡼�7��.��_���Iu��y��W���1C�␆����)�	y?o��
���6�1����o?�/�ŝ;�B0���/�|ܬ"FuΛM�5�f��C�u�a����e�/��4���������/'_ZX��Kp�Ǵ8���w�rl�s�(�l�������J�v�u$��6������[�=4	բ�:�M��K�݉p���O�B�`N:��Xz�$CV��|!�f�ʴNr/_8��1�^[��٩���X>tgi��D<��~�u�`lr��j�**��܏9��ѕ{���ew�������Ϙ��)����ss[�9�N���]�2��f�v������r��
�nTnc%~�˧�e��=���%�q�"����8j�+�mq>,�9�]G[%e���&߬���N|��]7'�x�%�fA�%f�)�'v��x�7���G'���tl�BsG��A=O#�}���?]�~z`���31Irh�j�Ɛ����T	�'!�h�:���3�tTn�z{�+����1��q�#� �Qe{�Ƭ��Y�o��\ɣ�f��6����?�ؙ�B��A��a��d0��K���SA`ל9e����ʾ��q[Ȳac���R��m���)I~Nu�"��(:ч pQ臨�Wl�UYLa����>~T��8� 6=IH�YRL���F�#��Lk��Zaߜ���Y<���X��f��xT�rP��5!
I���I��Eҵ��M�#@o��><6-Ah}�i2#.�KX�h(��밌� �=#�%�AaR?Xb��`��m��]�b�ǃʒ}�s30��J$<*I�_�]d�Y����J�6�p��>��v����6�:�W^&hѩ���#B�u�A��U���F�$Լ�3��~l�\��(��SJΎ9jW��7.��GYX���L�+E�T^L^>���m~L&i�oޗ-���k����n�j�Q��T�R�#q����s�i_ɥ�#Wid��2�C7+W�3e{]	�zO�k�u-�i�T�J�Bz^�z��F����@�	�T�-�- ��u�e�_��\w�7a�C�g']�w]��1B�:�,��K^'NQ.��$�����I��Z��j ��8PR���b����[�2EM�JqCZ�к)�S���[F��ݞ���I�vBCi���jLҶ�dQv��l�~��;��٧�|�AX�̘���Is�ƛn]�XJ����O�1L�b燄"-���3�EXB�f�"���	��S|�&�a�l㔴Xe=SE%�g�v��`�y	d�p�|CR�o��Ѡj��wL����PA8�f�Y��ZBZ�yR��Įy
r򉯢��!J�+�� 6c��G��*΍
;�с�zȮf����v���T��K��!\0ο��qY�|��;�$�;��:)�icFh�?i��vѷ��[�X�a�~��S)XWN8�b�)-=ݽN�#�Ѫ��q#����b�{R��\�32�N��{��+�Hi�]\NJ=5��n�8̝���,�\��̞�ㆾo�?�0*>��wH$۠Á�@V�u���{��<0��=����v@��C�x�HR5����l)���t8�E�J�k�u�����@�ձ!gi�t��^�\W��ec�#?/�
���Q4m,($?�vj��a�Ɨ%��͢�V��)�2��Q���`���x�.����{�#��HW����`�HY4���>(��� fU�,��5���������'���%�K��=f�)
j�Fטd��?������,^`Lnֱ�b�說����紵: <�ޥW{�a_��G%�[�/�Ϣ��ns�u�*�Q˰��풼��i�GkO�e��}I�i����F�OpR���(��K؉�����,Y~�l�x��S��6W��^��[��m���"�p+�M��O����'�r��4]��)����[�VE�y�V���(�x��Vk��o�w���h�l�c��h��[��~�P�`?����7��7�X~� 	 ��c��T4�c��nΰ��%t�l�� �B9�S�>y��{��2�L�3�� ?�k��Ո�M!��`�����k�%���K���f�;�Yb�C�0�){~�.�߫E���	u�><w�Ã�[���(����Èc3����\?R�ri-d�Z��u'���ϩಎz/`vv`��BJ6�^d|^т���������@J��!N.N�XLA�>��L%x�[�c�8�uu
��ҲLwfD��'~�Y�'[���9�D�NJ�t
�/��7+�� ��D��(�`��(I��P=�6��@��
3�9��R$;>zD��MQ.N�U5���ѓ��2B�BO�}�?��2��[
�q�8d��HM��	(I�d�^(�?1Q��c�RV:��+2���쁝:ĽK^��9��<�ğ��,�3���6L���n�VL���e����m���t���[j��WEm���0�f��dd�|�Q�O�K����Y̊I{(J�dL����-Ȫ�R
�W-o�e��{\�P�P��\�vq��e]�By�B|: ��`�ʶ�����8��׭1��.�Nm�D�|J�����G����CY���m=��wd�HԾ/VT��I�P�D:E�`�:�5�-�o�����Ӟ~aywK�u��+�Z��9(�'���՜���6�ڕ�ic��}�OrF%Ӻ���m1d�?�o{�u�yZ,�)yM̰:5��Q�W �
����¤O�,�#�C�1Q���*E) ����?Q�DS�jn^�>g�܎�A#|�*0�J?�o�1\ ��$5�ە])k�)0E���!C�ұC��]Qӎ��A�y��?]�4S�s%�>��Q��G�[��H�;�7��'�W���c	qv1����6P���._��v����⼋_��:;\��Ǆ�9�=�1�8Y�N'����@~ۯ_��lo�G6Aa�G�i�����@B��jg�$�H����mL���0�$5_R�9e��qA�vp/�P�"�E�F�w���z�`�b�m��^0��e��9J<����f7f����<�u&��fv��=�n搔K@�0C�ï�)Zˬ�� ?]�I�c�o�}�"7�%���.'����yj�40���4�Z)���ݵ�Y� -x��}d��l@��g���6�6x���_�ae�c��D^9�<��N��'�@����8�]@X���@�+���+0ꨘBs��ׂ�ed��G�E~ʵ� �8r	�te�X*�\�hŪ3����aI���H���]4��_�=X����4��Iz�#Ej��)y��L�d�_��I�\�y�j�[�UP�V��U��K ]euG���K�'���t�Y_���7�����!nS����s����mq��#��+����Үކ�J��p�pU,��b��x����>h�1|;RjG6���	�P�Ҝ]���!��	�ån�Xu�g|� 6X�������
#�<$�M,��@��1׈ �!miJO�Q�z�
\�j�{�v��|��Y�y��mU=4�!�ڰ\'�2o�	H\�*�]�b�1�M�fM�RƝ#�+G��fkM��.����u�@w��\��!�+�<:�=��0�rv/��j���(;E&ƈ��'*a���Fi�^��H��YS�P	��"�9۴�w�!'l�m"��$�ܳ�z�19nI&����[��,9�^����g ��s� 5�oM�ʬ�+|=��y*௡�m�}5V�4�
�����.d�G_�B��{�U��=�}%g���Q�N��)�9�m�7`9�"�\~���cU���,��o7��WQ���������1
̩4� p�l>S�c���Qoc/�]�Èo��BR5
r�����(~H�A�P�o��
q�,��`��0Eꠒ�AO~O?\��?�LP0�n�g=�D���e%����<�0\�iL�O�/,����\�1�	�<�q��8�.v���5gr�Dmf�a����n��Yx��}��}�@9.�=�g u$7�:Vo@��X������qW���ن��g/�g�k�=`�F�u��d,��l+��a���p��}ƅv��'�W�EB�X�D�d���@<^�B�7��چ��A��v�H��"e"'�4���k���t�3a@���3�8��m�Tyv(ہ��P�Xߞ�r�<�V�׳g�_��+� �S�椸	eL܈o�����q	����:�3�0��H�.O����4�D}��d��:_I5�+o�����9����SQ.w����8.��drL)~�+� ~@����6"
B� ��������!�G��B�����'���g�6��ڦh�Yd����_`p��n��o ��UOH �]8W¦x%��Y�:�-�l�������e|uL� �Đ��؉?��o�J��O�1�[f*�on+on�h
�#/$�������)@��ڿ�4����($GH�'*9z��s#��H!��cG�u<�I܍dY!s��n��H%`�$��[��j��Atr-[��H�g����lpU3��ޒ�i\�L��p	&�/a���.���(]~�Zx�[)�h>���]�C"�n)����_�[d��/��B��;�Y��_�=�r��n���5��}!0>�4�}��2��"�!E�-�O�e�BSϤa��S���pI�Itd���iwz�=�!�d;�������^*$<���]$ONs<��g7�+7K�4�t`��OljH-!P*{�O��Em�C���ó�$���]�������g#tn��T�������j˖�]��M8�1a�i!���i�X"O�`��?'}�Ιg�hu/A+`2�,�S�a���M!�G`T���l��ٕ�>":�v|���W���7��,ʠ�QH����I���%z�Òf���P7��ɜ@Q�9��)a�V�+4�.ֹj`K��K���P���}����\w׏;d���Ҥ���T�-k?wu> ˢm�:D�Q�,�oPI��~��]e�q�DR���e��"�-7��c�N�%�;�~�������Au樉��l/�|��p�F+?��L���;-T[3�c0�*���>�����b�F��~c��w�	��Q=�DT琗��Tgk}�&������${���'|^&<eby<�<�IYr�Yx���%��O&,L��1��'z��`T���>��8`��Ҁ�=/7���m��"C��AZf����V� ��\1
���#8L��9fQsMx�6�+�!�(ﲀRK�t2g�8P�K��8Q��rh�7�Bv�s���SD��K܌�� ���L�8c�E��\Y[��ܰ�<i��@�6G:�08��)u� �㕐��,yq� ݀�&p����޴	�!4R�;����ޘl,��d��X��,Q��Đ�f��Z���Y��XW�7p;ݮӼv���wq0��\���KY.cOň�lT���rٳ�#�n��AYĊj)ۑ7��^�%G����,�2�}9D��psS��Z�/�ƕ�eZ��v���z�O勒4����M+-z��N^t�#�݂V7j�ٗ�����o/���2Vz�w��� �Q���x&���]^�OԀ�2'oI�]y�:��C4�[� ��u-�[<n��x�8WXқ#�]�R�F}�l�:���?�x!{G82�?��s�6v0d��k2T*�gP������s/���M��IuO��,�BVOc��{���k<,���/tֈ�P����jo��:�9U�t̽y�st�Go
�h0�0/��wӲ� ��ra� 3?1��D�?�����݂��6���G&j��KҰU���/K�ab��3��>���/k�Ă�X����s#]��F�~����A^ǖ���?RF�&�c&f&,_93cx���nuM���UO;M��oxr������xe���N8C])�p0X�n����\�(M�7b�S�iC�0
�I��oن�黧;^S�T8�,M��f���h�>����7��x�se %s.p��PZ>��st��BF�]��U`d�����Q������Q�=�ߜ����@����[��.Bn���+#N�L}<s�jK?�E�
=Z�m&�Q���V���RB����
���ڴC?�������9}��I�R3/�������6�#��a�r�d��J� W�V�>���瓫A�+q�3S����=�-���/�����S^c"7���DI��ޥA#rB}�����8���K_��Ϭ�^���GϣO+�?�F����~$!_�������@�j8�������R�9�Ή�Ȕ�:��Fp\cn���"	Ia}x%�.�u��dQc�b$6ik��AM�i������~Wz��
BV����.m-8��[�9ȦmN�F�#�/- ��1<[z�����/s�;��i �����ڗ�����"��]�_��~KG��pE�����M%��M��[�@O���\f�ڴkͭq% ����!|���(�:�Q_����swu
����!�\���x����ۓ��cr�l��@X��iK�AjɣK�3rP�;_3�l�9�+Ǚ7C0?g<#������̠o6�?%WG�o��Z�-�/Mf<R,ֳ�2�ٞ�n6�Bڟј�&v�Y��i��		e�h�;I�o��Wz*	�k��ę�raUr�Fu�6�M[� w�%��?��������<�ƒ؉t�}ˮ٦�pm���AN�ܹ�GZ�,����.�c�Ԋl�8!S�Z�������/����:a�C<4�ۚ�l��Od嗅l6Qr��S�L�R��@�7r����}=����d�W�n���l����z����v�N��s�1���ڄ<Ҏ��٭ٹ��F��/�j�䅙��,�i��C�co�hi�/{�7�r%��Ja\  ���	_�ƙ��p�??I �ω�:�p�����i�s�_r+�7UUmE���
���f�BY-���Ȁv���P��dv)d���OL�.0��;��kSz�C@�<:� �����������{}���#x5E@�as6ޅ�[]�P�Z'���>�?���F�-��x��id-GH�3�:B�C7���Z&'1T0�M�iY)��Yt�KU��g���ܸ���s�������HL��}{�ؗb��Q1h¨G�-j��(I���f�X���_���a�ZV� ]�G	�|u��E��bJ�d0�H_��A������ֽG;�9No���ϩ���d����
��Z<S�R/���AW�->��D��]����
K�7Yo��W�}8�&�ͱ��9�r��I:su�F�F�hޣ�E�p��
�Ds��������3�ҥ�nh�3��
5��DO�M�6����4m�s$z�I�U�\�6���d���8(�=Ym�}WI����d6��IY�8|"�w9�2H\`�RF6?��Ճ����;9�\<M�=���CI3��j�����D9���c�5N�+]Rˎ����j���}4��ZL)7���7��e��p����}5`�3���I�C	V(f1K��b����&��n�C��&V�������ق�2`�vV�[0�v�������O��������Z$�k���NI�����E�)����˻s��/n��Y��O� �`Z���sʳU���5r���cWxx=�����?�Y�sd����Gh�� ���?e>�0Y� 
���nBrf0v���#��Dm5��l�	[9�����z���ƭ��b��I��6���|�6G�`
\6�m��OΆ��{�š�n�D,��f���^K̄<����@�t��
z��	f�K���V�-�OhtAopn���ֲNN\��������B_%$�X8\��A�v�V�/|e���.e%P5��_n+��S�B�͊UIo�>�c����G�J(ͤ=%V^T�� ƶ$2*S�p���%`.]�G�\��$�ЛQQ/ B)5�"!��;T�:�����>^�hé.�4h��s�9�gHFc��r���?ה�LӸd����X���|�Bŏ�B����)��'�/@��V>.��&�r��>1�2u�e}��	���J�U��7y�I��Z�3��v.-�
��l���"�N�7��<���T�����g� =<.�mQ%��Ϸ�g� �9t{���o�P%@q&1�z͗Id�Q��&|g�[�|���s�d�A��8rh]#6T�+cF�J�8L	�X��풔-P�� y���ieK�w�P~��]�{�~M9��Bow������hZk	*�n�rW��R�dM�����u4�\#�@���=P�\X�3�����@��8�a�Ys��W��-=[��m��C��]0&�.t���kԿ�k�i�&��Sv�;�RWB�X5�F���� %oH�9�VV�I�<C,\d��A(��8��Y���� *K5~$[f�a�K]�."�+;�p��t3i-
� <0Ӗ����g=^���AP�+���_E���_S��T���)d�%���X:��)�i���=�=���&�:�_R�5���~��Z����� �5��ǭ`�=�ɻ�������Z6L����9�u^3�ɟ���Li��cH%9��� 19;�2 n��\��Z�����.wɝSâY���b�>�دl����A(�Q7���Tn��͍���s�Ⱥ���̋֞��v�	�Tz?�E#�<��o�q�yX�����d��7�к��0C�)���󹐯ܜ�I1tV�2I���z:���fC�69�R�J�lY�o�P����-Gd�\wjZ��ĔR���gkԨ���6�}s0U��,�R��<1��/Z�@�i=�����vf/��|0�;�z<�CGj@�6.]���F@�o�pbk�\3�덬��T&Z�� nQ6����O�[v�����)��/��^V�|B�H?Ϊ#E��:�h� V��	N�C��/��3&�x�T�$���H?�23��J^����Xd`�_P����"�%���J
u��؛�����L��� ��_�i_�.��<�4p�퀐��h�NQ�NU\U渷�*Qq�
���5o���������-��B��E�X~���6��|XU���N��x e���ֿ��@���x�f)Y�譅�o}�|
�YP��1�W��P�U��.1(9�tB���V~�� -��oC=R]��r����R��{#uzK��ږ�}���K��	ޛ���ф_b�t�<������))���ދGѷH���Fz�9b��"�k�G`?�~��;�-L�������͋8C�q ě��P�d�ZKs�%oʭ;�ͧN�*����p]�N�v}��gsB2 )}��l��Z(��{4 e1����v�ߓ��b��V�J�@Y�u�����y��"`(a^����z�b_����g]��!���Ҍ���GF�
6�(���d��̗y{����_¬�BDj\_���{��"�1�'��I��S��Ժ�O9�V�:T�1��(���{�R�V��e|ݚ�E�(�U��l���ݥO��E��E:��1�nUԫ�7q������륨?��Ƅ�w�IL�Ր���T���0{��u�f�?�N�w.q�<
(�,~'~V0P���i���� �"��JTn��!]i�Е��w�ȫ�s��J�t��U ��%ެ3��� �Rq@��oU��B�u�b!�pS���w�bIsΟ�Q�5��Y��-sFf�E2��
�I����ЄI�P�F�9n:���x:��g�΢X~��$c��8+mYu:�c*۪��^R�s�w����AT�e��^-�>Ց=��厀 ��o�R-Y|W��A|CE�%�J��V�z�(���pG��	2�n&6xjX��<xP��W`���a�M���jM�o���C��\��?�R�E�]t�Od0}.>
��\U��A]� !+k"�%]��3��HP��QKq^qUAQ#%��BĻ,���<o�|��jz~ڨ̌uº�P��Jy�b����_YN�:T4�±$��F�qM�K�q���0@pu��/V�A ��l�p�hLx�T}�y�3s����
�v�ML�V�������>�v��/i���m�(��;l�n<9����X-�r�*�ã�  j_����#�!�˄�>�U\5�@%��yg��_��#�F	���Ũ�����ٰ�l�5��I�H"�Hjw�v�7�\�\	s�\p��B*�x�T̔�W�ʼ>���ì�&y��G�+gw��ä����fW���,��,�����QiK�=ϟ]m���9�$�8��4���q�'g;p��Pʊ��;N���{��Ta�DTO�љ�o�5�A�ǒ�7��L�[����ș^��4�i��{AJ��N�7[18}&9CK���uZ針�/��"�q�[�J�V�\�B���QNd6�N��1I̧�Γ)����:ăKZ<��A�=��A������3/m����H*,�>+�����~��?G4wbt�M��rn\Y�S��E��v�&%Y{K�D��o�Bj2����,A[�H����Ǖ�2�ؠsɉ<����Dq/"&�YK�����3�*5�U���B~\T��K,N�U� ��f�ZZ\�q�d��u��8���l����n�&U+�'���n��>y�#Y�.Y��ї�b`��a'ؒUoJR>��&�@L]����������G�5�'��g󒲢�~�Lm9cܛg�j���=)v[2Ј,J2��N�P{��v�2�.(�4�7b?�}4���"!rW=5��x�.��Ϊ�v�	�ddVk�ھ[2�&��0�f��Ҽ�
��ͅQG�_=7��	hC�t�<7:ߓ���h��s�9#�.�KՋ�PZ�L���7�ͫn@����o�T�R#���Lq�*P d�;U��ў!�"��Z��&Q6*�}t����S���겧��^4��I���:w-��4����<~��7�(�����bΛmo�n+�$
�'P��'e~�W�����M��}d�hRkb:�r�
�xH�]I����?��K�%��޴��F��[���
�s�i�Y�j�x!��`~y�i����$� %bE�3����+:xR%�����41��}�2V������-Ou��	<W�.�3���2����>{]��8��cM�L�VV���ڭQ�v"=F�qZ,�#�`�f@V�L�f�m 6|�!�
L�����1�+3zD����5Fږ̅�/1"b�W⟐��ы��6�Tڪv���#����
�6	`�r������Q�[��L` R�e�W�����|v�[��ܲ�̓��\e����ᢍ7>�x��uC�c���
z�˔ �@����w��Aq�>��F$���%3�m���AF��u�/�0i�I��L�&���R�������E�����g�[Ȭ��aOxu�OLM%{ܲ��!!�W�*q����8���&�5 h>��B:���뉰�0�eEJ���qn�uY���ӌ2�� �	�>����Ħ����_�'�b�0`U�l��~�_�2j����o��{�8w��ۖlU	@�~��P@}�x8}�ֈ��z�=R
)�}�u^UZ���(B_ϘYl�BK�}�M�����C������AD���	���/��O��)V�l��)�o��s��U�1�Ȗʅ��͜��
�~<�ÂL���,�yܖ��||�M� f��|� V�{+b'Zl�o~J�!�ǿZ��(e��8��ӭ�!c��3[Vj?��ғ�K���zɆ!��<I��)��/"�_RT�g�:�^ݿ5�w~[�ʑ�t��ޘZ�W��2��%��2�uC:�����W�K����Z�)�O9���64��o-�%7#k�mX����EX^�CL��[��$�w��ݼy�"I��T��X�L�e{�m`ƪ�'{Ua�y� �0J��YMy#`�^�����:�EQ�%ڛ���Vz�@�Z]���0�|�;���w�t�<��<�ڊY��-�6���l[x�l��'�C ��j7{���a���!#�$Ϥ4i�`�ȼq�b�4 �	0˚�W]8�������3�Q�:B�_:��E�(SJ��Ϳ����;�]UɈ�2�!���IO)*s�G���ӭ1C�r��Ó��턁w}�_$e�5���t��EDo����l�D�W�bw�U�!$J�;P�⤽pJ�`w,A��� h4��[��P�����E&��]_��A�i�P���Sy�)�����Z,���胖��m`�~x���j���X��;��v��@���,i4���L,��X����+A��|�RB�N�a��ƽ��P#��C~���,)���p]�rr���ƜF+��if�W�Ȝ1qs{�)]�+a�4�3�����q7�Ĳ�F�46������]�x�S�uq�P�JX-U�=��|��O��OI�W������B��o���^��r�=�l49�����N�r
5u��֭{���-�t���!Ğv���b�}(ᛛ�j<I�Hn��"ȥ ��Y��ՑE��n.!2,y��}��fM����reA�����{���(�[m�`_D�u��[����D�Q�Z����E�䋈��[臹bK�`�8��[#;P%㼹^ܚ��R�oڤ�r��z��O��{ر�~N�<WH��>���Z"1]���f�-�K&�w�����|B n�8 �:4�Q;�G�F"�i��1�=��66	~4�dki&���X��%9, DV]��n˨k
tܞ��g��}������ ��
�����0�t�h�d�6�P��"���D�y����.�T�\����aGW�u?����T�ڐ_4L���^�,U �Ki���4EZ�ÝV�oZ�'��9n׹3�=;�B�6A~�9��c�)��ru*̼��b�Z�*0BS��2/B?��'�!�����!}Nd�;n��66Ha-4d�ӿ[?\�=�l����o��������5{G���g�9-{�ٳt�����U����)�O�%��v��'F4N�Z�b2Zف�S��c^�$V��Lx�ZS�(''h���7z�9�^v����k�V�qì;��d�����>�ե����jO�%����c`���ޝ�b�,��IP�S���k��e�ˏQ-���ch
�Q���r�cr�e9���R���6���%��w2�SS���gteN��\�S���&�c�V�\���yy�7-�]zl��ؗ�������#0R'��{��:��x�q��� �I�?���x�
�R�8r~Jm�ʲܱ��W�#��ޭ,#�Pܽ&,�@�����mT��ݕ�8�<��_����=<��x�C��h9N��r�����c�5Mز��ċ3S �<>��QmI��	ޥh[3�/c�.���r�x���V�Dp[��(v+=GN����{�>��Li��9����2�/�%�6�.Ok��8&�U+���P,��̻��L��,R�ȑ4+X�奁,[p�@����S#M��P��-��f�2��V�|3�w����'gA��ڽ����LQ7'�#挒�f��_̢�4G�\�I�6��`:T{�4��N���z��8����_!���JT?��Y�	1��G6�|Oƚ9j���m��MA;��ٰ���l���*���b�4�!�![�y�q�)�_:o0�/�&�1���0k�a�es1H~�X�lÐ�e���]0�������i\�� ��B��r����&��?�˸�˼����C\TӐ� $o��歫�F԰b�3�7%�������9���D@|U�!X*�s��z@P$�sJ���1D�w[Z-Fw�k�;��q���9��i�z$�`�o=��c����Cw>���J���Y1xIQ��mL��(]6.1���5�����3���Խ|ڗ�]{�y&*i��������<��e����x���Z5��Ū,���,Rz��p�k��s��!oa�hH���pA�Ŗ��9�8�AE˙�D^��z�(��逈�����ۼ���{��\��:킛���
!��X5��L�U�Y뻒�v ���.(���8���d>=�ˇC�5���\����s�K��kv�a��p�vB62,�=
'a��^K�LR-�y ,��6d��a2�k�|�+g��~��o>qt#�<���D�k�%�� ;:��o�ԼX8m`���9������k��`�g���wFU��ˣ~��M�Բ�s��z��9ऻɔB���`���ыHL��7��JM>J��ߤ�P+ksY��W*��_סq�)b�u@��HOl݁��_���t�Cm��<�_�}�?���U�qe���E����z��=b���h:��KqۄB��K+v��z}J�1h6]�	��h���1q�J��������:u�Z�Y��ϖ}�� �/�S�sgDo�J��O����B$�ҝi�Hꤧ�l��}��2٤ldY���q^����|��w��r`4Jdڧ�
�蠭�����!7Z	9��F#,���U9���D�v# ��@D�)�1;7���a:��5F;V���˸$p���4�9����Z�gs �������>=�T�G��l���5�lV�4��<S]�����-Vf8���H:�B!��w��o���gZh�$�p�A�:p���%�$�6"�U�����̞@�Q?�aZ�[N�<�I���QU�=W���L��9����2FC�I�s�<��k��"���̂��090���"T{����D��o���g9���F�#�c'*��V��~O�>�d�TCv�CB�.)��������n�" A������-����r$B��J��e�E�%a�rG	����Z�?$xbz3,�h��>?�ꇛÓ�������cݡ�\GY�q��s��XG)@�{,Gv�k����,�߈u���zV%p�ȎEETĐs[g3D�{McB�ћ��w���D���c�5#?���u�[�=h��F>h�! +u��)F5�7�1͢ӼqI����.h���9A��֞�&u��	)���S'�g�m�|9. !ԯ�{���)�{��R��umQ��c�5�Uo�x44g���K�?�,F��S!�mۣՕL��ݢt;��gy�,wIґ����9
���ai�ufX�&J����|x����m~������<;N��~E�
h�O&��؆VyAxs�8�i��X�h|>uK7�y��Y��XI�X��G�����v�IL�+v���v�g�R����=cs��E��B������ܧO��>�U�d���WQ%��-�A� .b��O�����d�{���D��cȨ���>	�8��4�0��!�;g4�����g�,`�S��g*43��-���M1�k�[D"�N��g!F��W��TUR؃".�����f�*Q��G(?w6YvR59�IW�{���Y\�f�m	Oc�?�]�B���iY$Z=4)|��:�&"�_)S)״�(Z}M;j/x��X�K9��}!F�6E�Mʤ��m��#�����*GY���r�3o=��y�RWJꖟH��{+��1��Py�Ξ���{�����:�.���$nͶ���FT�g�k��/�*7Ԧ.�Q����Bm�����T�=- �
���aà�R�V5Ȁw�KAƴ~������;_��;�e����)�Y�BV|�-��6]�ڏ$��Pک��U�ֲ
qd�1М������S:b��}���g��������2�O�R�N忳��sZ�F�^d�Y��ۙ($E)E������ρ�=kG�M�$�����e�8������Xj���U&�����,@�D�z�Yň�?�,{o�����;~�s�"QH/�5>dg��| ��`[gC֯��@Mj��R�Ht���1>{']L��!+��Ds:�%"b�$���{�ML�s���̂K���>���8�W@-��nz�-~�(�p�t������ $+	 I�14�l�[�1&������͹���"^gḟ���Jz�P~���v%\k�C�e�h=Fj[[����xT��*Ӥ��|�0ȅӽ���@)!9�������;z��A�����0���U���M��ae�K��dǣ�g,&��򜅀@�1��&N1
F�� ��Q���7�v�;�:�%F�ø��r\�n�Κe�np�ڦn�~������vt4m�c�+���(�+y˭�9��W�[Y?ic��:m0�uP�/)�4��!TI�wB��E7g�:���)a�L���R�i[1�w�or1i�/��=yTꁜ��t�j�B2B�wM��yU��� 7�U�G��I��Aa�z�����AFi�	Mjd� ���pq��i�p�B� �KC��Ұ��	�2M\n}w�l+��q��/sO�����y����p���Na[i�pS�=���]��w��IJ�*p$�V{'�pg�G�^�4���j<��6��5���(���;oO�o�z����HIV�<�Z�ʄ̷U�P�ٖ���lt,aЧؚlNQ&����N�h������}9I�h��LkXoޫ&#�w���@!��hO���=��	��Z9�1��4R�޼]�_R��\l�j\�T���A�~��JȯB���VaS�p�� X��-f�E�V1�9�������^#��..+97m�!:aA��I} A�꾡�{��;�w��+�[�]���B]�4Q�y����%j1��n��*��<"W�x�Cƍ8B���s�s-���^D�Ld��5�!9bH�a<����c�F1���9�5�^0�<j���=���DC�h����]�R�a��'�;^r�a��X�=�a]�p��*Uoz>ϒ7���&��+�]O8+R��O�F�g_��v�x�8��9vPT�H��JL|�Cmm"h7eDr�X^��A���w��]��e��m�����<�p%��(�xa[4�g��!�Bɍ�p���D�5��K:�3�T���d�X�Ԏ���G�$� �a>,�L{F@�L��>�!^��-�m~��"w�Wܳ �M�h~��N.@agc���I�b]��e,��R"#y�%����A�������j+^�Oѷ�x]@z�+���� ���M��[�D�����G����|���+�4?վ��]�?CqL��B�!5}�h����X��BQ/���t����P�1�H�B�2�K�n�cv?c!��-0	c��21��g�ɎMȲ'8d9Ӝ9���QAn�ھ��m��:�'
�<E·C*P��C���C~ky��7G�.-$h�,��¤�Ow^���9�	T�ǟ��(�gQ>lDu�����ص��b'?�NBA�v�$�we�:C�c ���1DJ�i�]B{t�w� ��םͮ�~�U��/F�l���:簬�z����g �0�9&Gj$VB`����쾯,�ޏ��{S��`��k~��v\L
�L[��o��1�M1��Q6�`Jq��OX冃Ɍ���]\L���fi�&*U"��/(
�8/*���JR~m�Z�+�2�����&8V�C�&7�4M��t��;�I��/�H �pɒt�>�T} v|"m��]�x8h�H�}Ϣ%L���W�i�E�W�e���C�����Ö"'|ϻ5ۢ����9���j���J�E(΢��J�C8S�������C�B����{Y�LTA����Ȫ8��\~-7Г����[r����2�6�*~
Qt�F�!�u$A|O��>�9S�Gw��������P�(�Iw.-��\�����?�	�v	j'o3������'�Nq1e�H��nt�d7���|���N�r���V��ĝе�8:���i:�Sp٩r|�s�5ۏb"X�V��_G8w�v�S7��q�`>eM����>�.�;�JHڔJ ��)�1��ˍ��M�s|���_k�〇� .��R	�'�Q�����M�,BP�,��_��l�#{�A��)���,��*��s�iZ��+`�agH6¨N9�q$Y7n,r�9�ɤ��g'�튷oe�)�*��K�j�1�5�anъW���5��S�T#��P`H�_�����_љ���}Dy��5�Z [��MEf���L�N�VS$Sa�~E����4͛C�w�g���-��T��	 ���5��μ��og��ٳ��)�4<����ԯ�S9�>��՟|l<$���.�V��'z�Ѹ�B��@�����50�2�+����A���8�_D��u��!a�d/i�oAC+�{ɜ��A a�B�b[���k������4.Z��*�����\NӖ\�]g��_w�:�%ź�~�7*a/��AC��&Dd<�٘�H�m�
��>@)~�	���	C@�Z����Ȝ�a6�O�U�m�,鵍 �Q,� N����s�O��1�E8M���0�<��պ�� =������Sh;��C+s�~��g h/
��쾴@�*��q;6�ݑY���[s�~��O�t���a�/N�<Gb�>��9������^DƖ�@��zͻX�� ��}�c$"q�zB���;�����5\��-��ډI�X���f��W�]X@�f�.�c�����&>�&5�&*}!	%�Yٴه��H�B�?v]-��X��U�p����;8����ؑ)���/�iC���x)gͅ��zܫlTq>��?bn� `Q��g_��ѩ6�#�im_Z%�]���,���,���F����IKi�A���K�2�"V����ᴑ;���sw9���aRh����.OGڄ�D����ٯ��3F��^c�q"�.!5A���4R�]I��m[��2$g��w6���p�@�fci:"�|g�i�KD'�&\�Ł
+���3�p�@�m�ZG*>C���qP�� �}N+;�թ@Ir�0�2�i|b鱭���ǁ[π�h�7X||���@��[��s����[i��x���
:�jUX~�m���[������3��	����8�P��@O�La���bAn3�*���4���_�c�Y����6��yK��\�Fm\�Qb�g)�*�u�Oaq[΅$
;DwĦ��;�i�����ƴ%��(v ����xPj3��x�In����=�4s=`��Zjn�Z ����C0����]զ��Q�a�VK�e���lW˗۾.2� ��P� ����#f*N�PX�U�'�(4�,|=��QD��[|��2l�^�(�8g�T�����\�(��%fcx�a�h�2";��L C6��CV��plR��6�1,�,���.S���"��J��M��#ڍ�Y:�*���?��3�P*���Q��"�ʑ�y4,�Jf R��J31���Aa4�dH�kF�a�Z�UU�.u�fZpC9�Og�9}���TȾ��3ĊВEl	�c
r�xڊ��BF9Y��U��|�i��R�H�4�@���DWgD�)aй�: (Ӕ��򵳩��b>e�r�H��,R���F�Q������7mꠦ�W�ɚZC�6��ok�a�|������$p������̣c� Gk<�A�}a�v����tߺ�2�-^��VO��SN���\k0F	,�"��/ژ�k�9���K���Z�"㕾�=��Ȟ7��n�qJ
���.�}]k���q�k�Ǖ��¬ڬ~��(�x�x+��To��8���&�A��f�d(�w3�"���EV��f��c�׏s��u�0�zK��[dZ}�g�N�������)cA�;s��C=!�_�|b�F�N���#��)��p��?�:���3�LH��/v��ƾo11
�U~���i���{�׼�Ѵq'}���;Zs��MG�4�4���v+���)����E���,k�=��,}ȶ��o��?��<P��oߪZ(Hug���7�ϝ�e�*��� �r�Kz��i7P��P*#�j�ct��b���o:������*����EQ2�����Wr�@)�0^�O�$4{g�������GG�~Lf���VCgG���O[A��*�=_]����h�P
�����(
�_e��*�y;�wXe.��K�2��դ��r���fq�=�ŷ2�ȏ�
���3]kL_����/vC2�c�t*y�;�#m%�� þ!kOz	�v��+L�HP1 ����&7(.��\��֤��L
�(D�f�[�~,���ՙzS������0O�}<�s�k9�G@�j����/<�~d�|�[��A���{34��X��L��|%Z^K��d���=� �����V�����B5���j��Y-F�'TVN�H�>��=Ԓ8bjc��SI&�f7��|�� �8��ۧo��m.J�Xӈu�D���M��7'�e�8�)�œ�Q�ψSg(�����;��fu�r���vȞQ�H����T�XTd�v�v~ �0ǭ�D�b��O��t�Gx0^ �E����wt����ޔJ���j�.Z�jGo+D�1��u���HѳT����kiJ�gn��k���#��C�޺�9	�,g(Dk����/���_�W���߮�{m '�}��=x��(p)]sBf*����M����ĮU���U�oxē*{5�n�0A΍�D�O�S�Y��w�����L�J��nJ5Pq����6Th��A��K��2[G�<�t�N�C%<I3���6f+]vnf���T��&��pB]�
7��q���F��޴=G9_�6��Z$:�c�����/[��
�5��U�����ym��$٘c�{Q��0~Y����|A�$;$�5�iG�"�\���]��W�� 5P�]r�njG��]cJ�kc���G���@��f�~)����c`���&I�vh�l��-
�3������^�>Ą���j���^�wɭ�m�t��\u͔��/E%��с��H<K�`e# ���;�r:�Kc*���B+�N=����)B}~�c�e�#��ov�2��d��?����|�ow��sr��-�{� Z��J,�5i���;R���k�kQ��J�Q��7<<�tL���<#�;��F�|���T������ ���2>��KA�-��2D����WI��*Mk �V�@��w�jBz���<da�ʵrk������֮#�lI+X�*���� d8,���ɞ�)���V��ͺ�� Ov����4?����ZX���s,�)�����Eqj�.>DC�a5D�ƙA��~�JY�C�gV���M��{Ӳ[Hi�Ѕ����&��Og&$F*'�v�+�fS�@%߃��ڞ|��a)�k��f{=(���R;�*��]�U��=��.�@*��J�Pj�U��~e�!��j�w���|U��˛��<]�3����j��F����C�[����G�Sm]������o���_`���	��i"�?<�3�4�"��p�r���`��m�`�Cv3f+��-v�^�L|gbP)���	��8G�(�%�3���A�=���G.�m6���f����m�����jl��xW�������Rg�T���JN ��LnV(�g�R��T�{��$Zb ���N(��A��HL��U
�i��>)�/�����p~��,!.���q��� 
b���C0�Ĉ.ޖ	ٖr[5�_�������FL!ߊ�J�{wS̅��� |�0�/�H^|p�mu�y��������:j�D��9k���8��~!o��Gɢܳm��}0횑��q�]�{Qc���I��
	 u��?�df}�@N�{E�#KV)(��x�cu�ɞ=���8���r����C]�)}�f�J x�jc��	�$y��P�r�c5	R5LQ[A�-��]$�	򚹅��U���.��=ežiw�^ܴ:�/�*K��D�e�( KtXN:��y������s��D��k]���f%�O���P�c`	z�I\�w��?=��f,�J,)F�u:�V��{�c7�m�{��a�����	���=Q�i9�%yl�W����(<���i�]�\���=\ڇ�x �BZ+�X��`���kb���]ъY�c0�W}7�z��8�����Hٷ+�b�����N�zKjL(oQ�n�g1����t�0՘�Xp��j7���
��3�!<G׼�,�5-Q!�<[~� b�K|�M���2��`�'��o+1�l�[�<R,��P�9�˓�rͱ>uj=yU���FF4�m��fL!���h��a�mJaw�$��=A=�9���*��n��d�/�����4Ov0��D˼@��i��N��L#~[��
��/1y %�!#��9&�əg��'kXB��&M���yʃ�I0��Pʔ�S�'�n�xsd�?^��\}�	�T���d��Ze'����k;9V���j�Lr���̚�e.���ւ+�W�{C��5��g����c�-�ϊ�� F 3g�#V
��5�[�b.���b��M�e����$�M��ۊ�h԰��3����Ƒ�r�6�⫔���6eS�?��塱���4����+u�0�\ٮ�ޮ0�K���3�>�}����P`��?�g��%��Aά ub}�W��{ν8p{���P���X��$�8)�:�Fx ���XG���m{�ҕ�!����b!8����L������t�4o��qF�g����#(;����_�S�$��1��Ma^|֦�sOL7�M>�J)�`<ZS�e@�I����񦹷�K��U�$�{ʲ�X���Q�ڽy���ީ��_���r��G������Z��s�%���D�l�~�=�P�.�
zޗ}�b�C��T�/�[��71�=��6����/Y���L6��}�{*a��MS(��w�S�.6zׁ��w�M�9$��		L|ЮCc����	ʲ z�+���N��A�0�	�����o�6wpƗ��On{�v"��+?uM=�7�����9��D^�f\MfUu��X��KT�嘿d�&p�E�`�0�S��41'�zSQ�O!&"��� ��g'��	�E���(\����usV��H�6VK��F��+�Q��T��Jp�A��i\�9���C׉S؏g�,P�ͲZf���=xfi�j�?��B��%�_�k�{RfBЯ�JV�!��9�j�"�u�cV��xh/��S��k��1i�F[��q5�1t10Z?j��ʄ6���� ,�N��dbv���KM�nE�Xz��])>)��cߕ�4h�aj+ۜXa�l
��,C��M����(�}�/�]g��i#��H8��A�����g1��i_����o۽2.�-� 5J�Zx�n��B�I)�6&,H	d$�>7��\l��핞�r|*���h��h��}��/P����sP�P��	 ޒ�1fN��[���-E{7_��,C���/��b인�A�����Ǳ2�8f������� �/�m%���Jr|��9��l�����>�d)�E��IT��b�8�!i��F�Nb:�¹LM�g�W�c�����",�픤Ź.�����s���^AC�$��6�b�QI7�/IFؠ���{w����g��.����|2�j��ug�����B9�xմ��H%D�*�� )��T,�5������*rR�����2⃽�In��7�F
�E��_b���pS�d��Yo/}���V���l8\�h�B41g�hk�}m��[�$eXƼ켮��Mp���a:mǖ��8X���lu�����o.���<j�|�bV�E���]U:5�^����שP���H��'�I/{O]�X����G��*��ۙ��|�v^�g��
���ΔP��bL����s�:�Zt~��a�j~%С�r����7�	����e��8:D��	�x�)il�7w�6-���Ga)���'t�dD�_����;���C#FA�����0�r r�n����x�yr�'l�◪5�l'��4����
�����g{AP�-�
�`��:�-����(/���ﳥNDI�g��ˣ���O6�7��j8����U3���X���,)���e&t4#���?׮������Z��r���l��*��Ef⢡��Sd����Ѕ|~٬��9w/}���*�q} {��m%�tr�śc`-�'3n�c���8�/�@,]
KƧi)��ۑ2,r�X?���ǋ �F~��6>�s�^g������$6�&�[5�s)�H��jV�;K
ӫJ���F����J�llFS@k{�{�c�ٱ�(q�pe�R�� `�f�Ϫ�Z��v�z*�'���Eʎ׫;��9ب��p�����`{O�8��V� .�����;X�&(Cңd�
�WT�ʛ��e1�*hV<���w�%7��,�y-�ot���JL[�A�Q�#���Y�g���w0GR����6��KK}1T�*�N����_ӻ���|a���2��v���q/h�z����N��z��*��u��^?����ٲW�j<tj5�6��d�2*6���#��Ap�P���8H�=r��;>3�43���F���W_��N�/f͂��� <Y��]�/����(U!Ȯ�QNs	��F�=�Q�鼫l4� �N&uڟ���tb��#�z���؃_n>�S#{~W
Pr��>��6:��B$������)a�r#� �-� /SqF�3Q�
hU�-���{IWS�M��kIǅ��Tګ��[A1*�s|��l+Bx�:k�"�~�҉�yz�c�[���"�#*�;����=C���b���v:`gS	�f�5�>��KS=�O�	�?$|	=�9��1��ML��eo����53	.;ΪN;
����Zw�֪�^ ��<׼�@�mPD �!}\�n!�Z%�ު{���7^��ě�OU'�MEbA~��
r:p��.|G�2��"*H�1�z;�G]a����C��� !È��n��/��Y�����u`)\��h�����[�G�����/�0^;|.8��Wp�۸	?;x��}�N���u��b�מ����I����fgq8~ܢ-�h�b6D,���o>�w3�#h���9�g��P�a��0|�o��Pf�v�s=����P�Mv�����v�²n��H&ǺSdҸ�ڄ��y�CPр�,@*eDꉵ���,[��$^�͕l]�`�;�Qg/X�Jn!� �g	�︼���\8_�N���R.�p@�
r��D|��]���Q����\�����������yVz�E�Si!���Q��]���u0�L5 �ۯ��&�(�[ ];5���cpx8�q��a��nBʯ0�l,@}���N�9+'�A�[-��3A
E�9�!HԄ#_�
%��=��]����;�m�9���5�Ӏ}"�B� 81�I��-,�g->C�ےr%��<�1e��s$XXμ��7����F*X=4�4svG���]�'7��:Y��Iu#��契1�Ԉ����d_L����y���@�</��?e)��!���~1��f�h���Y��c��]���m	��=�\��XQ��q<-z�B;x��0������$r����l�۪�&K�#U���|��k[�$��b~s�v<G���`�Ts��2�Z7P��.�_e�٢�7D�D��N��i�O@ax���/��$,R)ʓ�f3�?�N	Ս��}׳�߿�䘼@& Z��v�<<o���[݋�����${�f��5$��T��&bD���,.�&h��ͲB�v)�K�S�_U�^�s�"6�N	Rd�QR��_�67��ܑv'��Æ��f��2-�l�6�qhQ�6�0��h>�y��%׼�J�̳�@F�e豤�M=*G� �O;؇;�e,M��S����1*���Jyh�����a���0�;�pxߔ�,%��P9�B*#��������ty�k�T�� �)�ܮ-����Ҙ���Ks�Y����K�$;��M�[���kZ�ߊB󔸧��k3gv>��F�����5!2�ln�54����
�2K@�:��O�iCK,^��n\]���_�;5BF��]��}����C��I�K�W�Ci\�Q�)�5���m~	�Q�lcmX���2��ͅ�A�`Ԣ5(���[�=��G���u�1��'l>|��H�����qtxѲ��rU�(��6���d�1�R��u�D�V(h�+r���e���SN��]R����͓m֦W5��}�Ѭ��14w!�,��J��<Z����ƨ��&�Y��n��g���$�RjQ��#_�l�hU�q���-��"�0�W��IH��q7S����Ɣ���;��S�1�f�����7�#PSd����G#���<�OMK4�#I���c�u 9靨�\xy����0/���m����֍�W��@�����An��|6x�u1_�;J��EH�N�킈�׳�J����|w	y�QDU�*����AĀǱG�rI�C��u�H���-i�: ܻ���}z�D7��0�$��
�IDyN���C�������=��jg��E�\Ѿ�2�J���b�n���4�]k}�����3���@#213�<!�̥�8�-oΜg[ܒ`�N���Ը�������$��Ȇ,u6��
����{�z� 4>���x��H��>F)~��HC�����ಷ������ҥ��E) ��{��y{ H�eE�qZ��
(�
U^��H�g�3���j��Q��bW1ߺ$e�a���u��6�~���kqRyf�o��ƍ��>�����Fr3޺c�뤈	]�9�b��d(Ḳ�����&�d%L�����"��F>vU9�S�1�h�T�Ϛݖ9�u�a�^���"�V*��ֻҔ#�� .10`&Kf�C.u9�ɩ3���#�t*�iLК ٯGR�D��O�0��/r�|�֕�_��0��B����mO�����MT�{�TX?���S�1��E}�h��r��	X(r����m�����8�3��\�.L�W�w ��r9�Yv�;���ѽ�aD{��kq��E9J~�9�	q��zf{��Z���{�.�N�'�D' |\o[%?w"����>{�r��t�x֠[TO��k�; �0$��i���wF����΂6
!��v���ؘ�2c�°'��v{[��#I�Pc�����)�j��p��*k4��JM�uW���+�l{?r؂�:Q4��p����V~m�`��&pN�|mZ�䠤iEy�ȸ��w�CJ��۷�0�y�O�2$�#�饙:͓�����2�o��\Ǹq���Njo�7��%q��՚�)����;�,^D>��tW�����Z�/G���X�ro��I*Σ��2i��4m� �eP;��!���m|�?�'���x|�Jі|��(]�C����^��xh�=�}9`iEΦ�E�Yi. Ik����4'g�y��g1��B�/3aXAeI���E���,�meRf��&��[䬸g���յ��Jc�� �p���~��n{�V��??/��ܘ���)}�L�ᅋ�@z\{�=��W�wa�W��"b��8��iem��O�5Ci���	�|����PǮM�ZC5�w������3��=���y*R �ZW���5?���3u��Ru��9�sK��/�HWcj��p�w��cֺC/���S+od��5�To�t�IY�*Dt~�"�"��RMճ,��/�R�/#�*�P@x��s��濉$tq�4kR��/��W
Fו��3*����z%)����9n� �J:�טp��o��*�gkMV[��F(��m|w
�nTb0�v�ݎ���I�{���ך����|��wDYWq��
���!z�7V�'��{Y��PT��b�.x�D��E<���Ʌ5�׶��랥�0qF�!l�ڇկ���qmw3���99��+�E��	&��G�ɨك�w�h�p3�	*�f���"�Y�3���G��e9��ZE6h0\#X��B���/�� �n<���T.�eR��b� �:?S�T�WƩ���a�Ѳ�VR_��2���o�#��1_�B@5��w�vf�Uhъ�#/FY(��g��y'M��K�.�2ya�{�(N��ouԮ9�*KHVV��,�0����(���b1@���[v�1�9�{?{[{e��HGH��1-�$-�N����W�C���qq���s*�4}��4ŕ���?m�&
}�O
X!%��IFׂ������b���J/���fu��XBKPH�B��	�TBj\b,V�И��;n�jV7�FѠ�4�N� �|��+�<HR��f��o��<�B!nC�o��$�A�R��'Z��n
)ږc���f�b�	8��3�!�+�Z+YL����/�jNV��GE&�AWǳ���7���%�h��(�[W5|X\Oh�y�� �������J�/�s����_g-`�w�$!�����V�C,���w[��xn7��i�)8��P���v��G�X�L����q0��Cӣe������5u	V����ځI�P�0X
�F����8΍E+��ڈ' 2�����	�(h�َ�~�{�u�k�൴cfK�T�v���qï��Z���N��7퐍���>Cam�Š��t��I����|��5 �������B����_��8R3�c1�6'���kR�w���Ev�񿈚;��Il�|p� �?<��ؔz����\�?�r��t�)���9ħ��^	T���������K�<VW��[��j�:�~����*��j��9�IqcE�Z�S_��~��z�y�~�r{G�Q5O��:���N"~�q���D�){n���0���H��@��$'?jr�1�V���]��|��� ��?���L4~���~��t������5���aUz��ˑi�pY'�?�O@��=�}����zz΅_T�8���x��L:�yDc�� W���^��6��U�Y�)|
ű�D)-m'�m�t����o��;���-���M�
自B\�V��+ ��G�>[��`�h' ƛ�o}�4fА��h�^�(%�.޾T*����uF�?�;YZ�m?��~���-v��X�(Fp,!&~���)�9�����њ���� ��q7P�$�	�*E_1
^]}0F(���ae�lqG��y��i�~�5�����5�M�W昽1�^���Kd n<����a���wO�P��Iї%�*�:@[�������U����]x�d���ݼ��|t��]T�&��q��Պ^�5�!ԋW٭EAk�6Q^���?��ܤ�����wPQ�.+��6	P��ܲ�uw!ux�D�O^C�XBu�������Q����}Dlx/����"����Y�F��+_#�F)Hl�(��0�_�Opg�	mL­[�T���/����;��OtQ[r܆:�`7h�a(�-P(X!x�a%Jd�gNB��Ad��@�Y�QgOG]�ټ�sƻ
 %S�`1�_'-ee�����k��7�6��wDU�,� .A���hk�947����d~�E�/�!���X��l�j9��1����c9�q�G��,w�̹�/x���v��#'�7�5eQ��f�w(��Ɩ�����~a��e/��.��o-�Џ�e'}0�R�P� �B��VWQ����H��%�M7y\d��f�L�;��Ċ��en��o��Sɫ����3�)��B,EUia����Q� E4f͠~ ��^�J�!����ӆ���%Ӆ���J��/`Ǣ^b�:"	���&8X���,��3�*7��c���G�Ƭg'h�p�=Ò���+�|P�*�B�
P{W����!��;e���Q�u�rI
J2f�mi3?�Y��5�Z�ʌvT�YF�k��?�)T�g�@0҅��F!�P���������l���w$f�|	G�s�~�͟X[gX�eA8��)�j��?@ħ)�?AG�j�5S��
il�@�R��%�Hæ�K:z$��`k�<�ӿr�N��#���.8�Lsb5V�h�4�rx#�&cIH�B�U � ���C�~������BE�,�f�
@�<���Y�����M�!�\i����Y�ɯ�C�b�푎hNL/���<�z;�ZeC�mG�F����`%P�6Y�����nvYpe4�Fl�k�~B��M��ݳ�:l��P���ѰF�-��q�ݖ����P��ٗ��P�*Zu����t6F
������[@�G��e՛j�j��@�.	��Q��n�n�6�+c害�Ny�(}����q|Z�� �#(e��<G�����v���<����gDK��A�_�����&�͜�<?y'��l�@���z�Z�S*ߍ�9 ��?���2�ǳ%�Q}ݍ�T����KL�ww�$���{�8��t�|��&�Kw�/��c��g�ؽ�Qg;�piI&�J�3��!�F�?(Ur-r�;�1;{E�Q�y���r��:����F\ʺlo�7I��e4q9h�I��_�8�F��M�Ы�t<:Z��p����(j�@��(2���:(vK��O���ӯ��2�Q�m�^�x�M5F{�u3
S�N�"�o���C�l�� Qr�0.�p���0Pe����F�P��q��}�P��'��o;�
�%��yct�4^�YǷyHl���>���/��Ň�=-��!��>���w �OR�!�5qkH�f��y��S��Pbw�	����~J��]K?n$[��P��ZO__���Z6���
�z�uw�v&�/,Hm>�F��|8~�?ܱP�8#%đ�Ʈ���s�}�g�������7K�D҆5�B�%�y�E�y����y�)h�_bv��e�Kp������(���`7]��2��]��Ri':�X"R9��u���5�"7$�~�j�+VqG@Gg:I,=��ݢ��^	�\fU������}����00{q��)/��3��e��"�����>���r{k2��!����j��5z��(>2��k�Rj@�\�۶e`�,�=�F1��e�V����²7���^��G}�`I8�$��{?�]|�ft���2}pQq606��3�)r�/��򪲮O�h�&A\�!�G���r���0��A(	�9}����y�be�qي��o��K�t_�n���r1+s1�A�s�[w����'J]��?��ZX��-T�A��6�g�Rv�>�2&d�"8���(�����������t�P�Go{ڛ��6Q.6;{�Ҙ��-����K�:t���)
�+��&��7�B���2%����n�I@�O��2�Ʊ�y��4�c�*�!�6�0ظxw'c�V�!k&~�b	<Џ(���F��;�>&�fvרD�_&��$v��[Z��;�V�K�M��e����V�m��x�T#��+�ĕa�[>;�_�xf��_6Ud�̦�!��:��/�j��Y�M��԰Oxgt1_(G����un^�&�g�U?��}o8Ϸʞtd���c]��X�c�Jˉg�ؒRpßJB5@8���
V����H�F�)pi�UV�G@�f�A92���yjI����X7i��В�x�/}a��G|�:��f����`a]���*�G��o?B�/�	k�}i�Rn�,��y�F�8d��P�>�ơ�}E�4�/󤝰��.Z�(V3sZ�	�0^.a���U��2��\>�L�ċEه:��R��R�1*�'��9؜P��\��6��^�z,2�{�f8�?���H�����n��J�f���u�6�Z)��䢂�ޱ�U L��/(��.�����u�v7��~W��T�መ�p^�총A�}&E3�J�Ϋ��pf2%uki}9o��:y۳�*�R�҂��+�p�#����<+@"������[1[��D��=��A�Ǐ������ `w�.�!��e�'��aX?M�U`ݶ^�����l�Qǹ�K�b,��?�R6��熸�_�O��Ǎf���)��W=���`긭&"������y��ک�+�"��ĥc>�8@u��:
΅��M��ƶE&6���d�e6��HF��g��Nk1;�M>�@���w.��ݺd�e:ϊ�?����4Q��J��~�����8�d68*��4~�����F�K�Jm��Ylt7�������O19����Qw���i	G݄FT2��>�ؐ�+�)�ܥ<����,*$��ji�)"��O%<o��g�u�I$�-"��z��-`��A���|�P�S}�bh-�_�t��5���]���A��a�q� n�vwI�������	��W6_�i���,�Y>��4'~����;���F�7ե�ŢKw1m�m��$�(���N��f7����/vc�o�O>�.5TF=N�b0�lS��5;E��|A�2JXW<�h{c�Nη��l?`��Pq���yW����X�0�]�I�:g�*��c�F�❀���=��2Ό�&&f��#�����@G}����j�+�b@X(U'���&vB��sM��Ι��<�;&�L�]5���zƞ��͋����2`+\Z3x�d�M�����8&���Ӌ���%ɚ� �!�]SEjK9��|D�0n�7L�X����hh��ł]`��\Z��XivA�cvtc����p/��l��{_ȣ�,z��g^>P顭���]��RX��{���\��)	�g�>�{v*�p���h��e1Ds�0�{k�����*�Ik��z���ַrm�~��
�c��5YrÖ�sei�}��%��ʬ�݌�8�N��p��&���j4.�a�0���?��q�%۞s<hS����6L�j $J[O�4��U�U@=N����M
<`�����QZ�������ۙkhAB�Te�6qkwb��@�D|����Y��:	�Z}��gC]�33J��r65@t7�h�_���SHJl���;,dܦDu����'���J��*��嫄�u(�L�~�78ή��q���
��FG_b�&(~5�)P~�	(�96n���	,�@�$�ǯ�����e�W���$z��.xT!)��*q���ҫ0�5��\m��ٺ9��.z��#��v�R~s
ۨ�(U�G��̼2���$l��׮�I�8�`ȋFy����B�����H����������FDEBp]����$h���|xI�>�r��
Х'��u�j7#��=�mD�G"�����	w�0�E�^-��&��Z�޼E��w�zB�,��.X�(��D�]�ǥ�T���,�qd��Y6FF����L,��X"�����;3�ӹ���a�7lpV9]n����[k�,�it��s�-�
}6�O��S�>"L�x�"!ұ��l&'�g?�'�T=U�dA9�:�0�=�!���^��(_���lK�F��x�1&��'O]J��F�2y/��/�DhL���1�AQ(��BU���Q��{�u��8�M5��ɣB��n�T�`uK)�k�b<��p��dJ����~\�5��h>����}i<�]��R��,ÿ�p�B�k�?�*m\�#+�W�v<�]���D����9BA��Ȫ�%"Xg+����R��Z�oS��g��չ�R��i� Ӌ���Ntj�3aQY��v�3loy��A,��#����`
t&�-r����>""Q�A�_,}7�wI^.��p`���VؤfU���eWw�����0�/2HGӹI.ӷu#JZ%|�틛�����������i�pH#�&t��	m7ɄS���gKm���s��m�!Š�h9!R�'���aK��x�<�f�����%��p��0ByL������1�f^�ѤF��^C�i��I��m{��V�I�`�����g�������o��=�)a��Z�[M��IFC�#P=��;� a�՞�ÒЄ��mN|���>Xx2�5^ S@�h	�����C j�9���s�&���*��T�afF����~��.;8�;H�vqS��9�!�!Fg+Bvn-ǘ�t'�����IW�1偭���� 3�S�����1NᕔƩ>Fh]5;���l��d^����X�~�A��ZÈ�B:�����#�n�b�n����\k�L�h��ȺNs&:t002��BGs.u.���(�zƤ�_�@���X=i���R 1���6JMb%ɺ�g�\�<}�E[� �E !t/5K�9Q �#�C}�E�n�\a�ᒤQ�i�vi#f��/�±������PN݋� �@��G|��M��O��rv (5�2"��'6�8K��jZ�E�����(Fަ8)k+����K�k��wZ�7_��swM���'5G�H��������2�8�YַҌy}xz���!��Y��������L����,yQr5GnhRE('��|�d#���R����!�;O�#J����{s�����<
�<g�k����!�lщw
�riE4���3����� 	�сV�����<a>Ï�V�$e��6�t����%Ps��g���½��#�uSb%N���W�bB�h�i��Sy�lH��'?F3���п��_�j"��d���r�S=���'�@l�!YX��1��!������Nxp"���k��?�TG�7���*#N�B��%���D}��e��;}��2�7��r$8�sq��ˏjp�zT�D�i�S#�U/�wy��.=b��J�-��2��Iy�ҩ�}R6.wK;�\�-��^���0٣yW+u��.*������鬒�(�f�N9�a��2~ֈK"��v�k�}S9�������t�c����8�Hτ��f�J��.ӊ�2�>ww�R�We�e႕j}�յBw���BjĬ��Q�?�:,��[ �H�I�:�;ϭQת��"ī�~�J��T���w]r�Jn/.�cB(wD+��>��I�i^*�i�r��̎!��z;�C=��6���}��و��/2t�NwKG�E��м�a�b� ��dİڢf�!�[���8}�[<>� r-�~�s����,zou�Uɶ1܄7ͮa[B�;ݰ�=6h��t��)��ݬП9�� ��_.�2���T��ƞ�=|�ט�I��ğ),P�w4X'/�d�S]�N+oE����x+����m��V�~˄u�B��%�/S=�Q����]�7��B�]�����-�#uM�!&����Z�#�G����15 ҳ�VԨ&.ia�J�B�v[��i/��Ոz�����ٟ��.9��n���	'���G���?��j��y#�G;�;�Q��\�S�q��0���s�阬U	��.�k�U�Xa1��+�Zq$v���E[�E��^��'�`�C|I�h�*�A��;���0�R��n@^��UX�M�Z�^f|��~�NcOt�+�������*�˄�-�z��r�x�:��ek��SW:�,
P�茕�ɜ��=І뼆�
�����0~�t�!V���7(�i�=O9��z��0�B�Ah�J�S��H�ԟ�h���_��~�Ci�8p��pqj�Ft���ë?��<NH�r��;r-������*ǡ�v�ʥ�����[��꣖�F��C���fޗo�'���3<�*3~�V����?RU���H�@��r�u���\��2_�Q|����X��%��8_<>���D�8��Q�Ή��rT参ƪ��7���^��1�*��O���fk<]:*����0q &���< }!&t%\��f�p��{����_�������\	��d8-sϣ���Ă9t���p�@�g�8���>��l9A%vm9�� 3H :�~@�ڳ��ƛ�v1�;S"$���Q�'��ݪJg�K�㝶��Z����_&�CvH�w[�0}�Hz
�j��M��G�ꍝh�o�i�%-ܵ��!Wb�s���ۤ�Y���E	3mi���48��$�Ҳt���9 Fl ����Y��2�f��lj�R�������!.b��|�]��qW��dfy"T���Af.�ai��٨d��Vp4�~(��H�� ՄI/�� ��o�Ϻ�n��31�
'�� ��P�4���E�ڬ�!����#q.8�,�����"K7;�T��x��;��*��>k��K��Y�&�f|�ř�������`��<kW�;MnG�j��2BĄ~cҹ�؆K�ԯlH_*��%���g{a`�'�6z˿�Y��\L0�N���5c�&ݦ,^T��lk][�����$k�e�?���E�h��F���Nh�EI`!Ɵ��V�MO\�����:Y'nED���*���vl�ĴM�Sc6u�!UԢE��jЏ��F鳰5,~�!��c���X��b��/�&���|�73
Ot
�����_�(m����@�re�k� �ɕ�]����\vebok���� zL��`͚4�;R6j� ����,s�,�sJԭ�+2z�i��Yp�z��h֩TX�9�n��FzI��j�j��=��f>�R�B�$��5��#�IM܅�Z�$,����3I�1�	Ȇ%Y�A��C�>g�v��/�+ΰ�R��K�go��V�,�:ӱ����?�+2�:�}(��V4��lƍ5�Td�@�B?nP��D!����Ls��G���j�xϜFԦ��`<`���~�%W۽:&
���Kh���?���e�����v��&Bq�X��e��Y�c�*�Q}1_իʿ�D���->ȯ����;��ɉw�U�#�xӈ��A�ʞ�7�tṫ��$���a*��"�3P�^�Iݮ�T��P�zdi���a��/�]�u2j�YPO}02�@��fIq���t̸�4����B��'��_�^�8�_)h%WtO��I?�.8�ꊜn,�U��R����ˈ#Y�>o�댄��R�$YJ��q��[�r���9X�Tޑ0]&��_L�[CŚ�~�$̔���ϗdz/���(믦V9̚Ps�n�Q��ⴓ&Ǯ�Ԏ|��&��s�_G�ȸ���w�"�J�/�T�}���I��G}��%st�,������<�hƔXZ�9��q�o~�w��D��}�%�̏	�@�W��w��UbTk�0���Kb?SN����o2J������Y|�7�忓�.Hmw�e'��>�a{�j����ï�ڣ�"jF��p���p��|���3��,8U��##�ү���V����'H&� �U4ԣ��l
΂P�vH+C�4fRz�6	@sF櫲]�0���+�0�rΜ�ABa���Tr6s���Rma���}��jY��ftBwk=H,�F�	ET
�N^Ԝw�r���?���L{�~��:dr��c�s���N� �f�|[��Ԙ��]�$�gG����p��&�}�S�&;�PK������?6M�o�yF_��nW4M�sU-�����Q�OC-����Р)ܟ���F��Fˊ�{�(��YPcG�ɯ�e��	����{H�PR�W��ܮ�k>|UZ�^��>]S�;w���H\s��M�:��Š�����nҟ����|�z3�F�+���2�byJwP�GIA��'E��m�aQX��/�Kϗf,xA+���IM�!����:a]�%�y�r`�>�S��ꛌB���F>�h%����gA\[�P�)8
�g�����AA�x2J�}T �k,�U�	�ȃ�k�/�o.F�%p���`�|���F��j˺�M�����#�'UF��j�F�'-�vdB�U
$���!�Ț�w�6��T�8)����!߾m�amX��x��g�Ɏ�y�y�	���?l&�6Q��";�5��ź� �x�%�;�7,0�q@�1�g�/�%܅pݪ-��."e��&o�~�~hF8y$?�"TF��@�����
������:f��_��i�<#V�B-�c���'�`����ڜ���=�5�*F�(�xX�U:�f�o�S%�����X��~D��کry�BǹO�@4[U�zXL�0�G1�9~�ap�=V"!% �6G�U�������FV\��+�=K8ަ�n��眖���^�K^EYu��Rv�`����� �w1��`(����� �*d�g�ȋv�ë\t:fBlӗ�h�2������1G}�X;��4o$%�b7~�
;�����1N&�ג�k��N0�JK@��G2Ĭ�z��V,rJ�(�����Q߀O$1p���g�ai�\W����� ๅ�`ȯ򊚙��4?�4Jh�~��pW9�Ê�k��#���M���V�E��Z�Fuӽi��P��=������iM�R��^W����p�GÂ��@�c��[.@�B��^�^�����%������AKLx2"T����✄���o�����,�܊�����zиf>:Z�Kܼo��R��j�)p�YyU�@�Wc�Qt��ta�Q��5�pq>N��0�D�҇�r�����)J8L4���l�����>K.گ���7!6K�+	��Iř�{D>��iI췹J;��ƭX�T�"(Lȭk�/�� 6{_@��0�ﳪ�Dx�&Mڟ�s��-2/'���D��D( )܃��*�	`<�+C�ak�`�������
��5Z�γ*.�>��|�������{�h����3�r]��UׇD�vYA|�s2��o��̷
H�m�H<(A�L���UL*�l��������LRG��z���KF*D�7�ymoiup]C�18W,����XlӄY�r"����k�a<x���o�}P�c&�wx����(-�"t_�_3]ĩ��>j��'#�s�س���\\I�!G0r�������5���ӕ�'�vt ���Kcy���>���)���Mr��eZ�n��_���]4�Q�7��H�ˁt�%T|��w��5�	|�*���g.,���%���KOt���]�F�H>ܝ�%��Z	?�6�2�m'��wx��"�x��0�]�^�u���E����]w�V�"R��gn�J-q�h�6hQ1$�췏ͅ/��]ހ����<�t�h o��BbG��+^"#R��w�H%�&VC�V� ��(���(���#V�>w�⎢#f�r�c}�J}������X�Lq=Y����0��������Z3H��,�$��+zBd�B�ֽ�Ȍ{�¤ǖ�ER�Cfu�{�Hb�ͨ	�s(�a_���>k�6s ��.~�ӵ�0g�^W{mLy��I���:�S��}������Rz ��$�>�D瀠-�t�;i�pצ�:m�S>�[��[�	�ձ�L4�,kI~��"��z�?t�	%���R���ƣ�_(m{�A���o�ǁ�/�+�7`�0I��q�#�{Gm�&��v�.�F
���s/�kTw��64L,{�M6ñdu��i_�4lB�z^�A/D�����c���`�CU�FE���[��JH��cޗ�%����T����e�s���� �-�������YV\��~;8������Q�:�h;3NtV�
e���Y�ʎ)��Ty:u�z�:��NW�6�8� E��̵�	��q�b]K�����.�;���	�R)��K�]�e����OD2R�ZG?�! ���v�1Wz0<�"3�<*'��Wmǎ1��?��5 �P��l��,��TZ,m�i-�B,1K��&*�/ �ʢ�V��kD�0���D��Q��kL��Ee�Koј�J��C��O���u�R{����G�5�5��PWyٞog\Κ
�ߏ� 
����Q1s�0�̝�lé7dQOW��Q�D��<5�\���:q�O�����<^T�ʬD���O���/�(�g��0����V����ޖ�;���}��y-����oJ��f��?aV�z^?�'�H%���qx���þ�<[��x�6̷A�:���G��Wb�Eۘ2P�4�w�`�RR7Zb��	c_���Ω!(E��Ye����5C�M�Id
�䙿o� `�Y	��ԞމS㉶�2`��\b>V�T�w��?�#��Ti�y�ԭ[�b�E{�iy}�%m1ʌ��G��q����f�2G-w����xKU$�ll�6��5�>��FR�]%;�Hƽ�#��ꕴcU'�3����������:���Ĝ���>��A"�익؆���b��Ay���r����D���3�SAǏxe6�|�5�>�֑�6:O�u��u�v�[��yO��i��R�\d�KJ�TΓ�aW�R��a������?�e�ހ���m�Ǒ�:�A����6�G~�B����+Wz��4B^�Q]9Y����>�]	��;��̩񠕩xW��h7�PV�O\��4^uL����~_���V!<�c���$�|���6�ף		��e�H�B$JL��̗�H�5#M��a���u�p^̡�u��)q7z0f�X�����V���u�Pv�4}3{b��&v̏��ź0���Th�5൹��vop&�#�O��5Y>~�_�, ����{�)sZ�2�#ʖX��˯�I����ȟۼ�e09�޷�>�m�������e���]�è��ς#���a�f�����D{����܁3z~J�z�}���Wg�y@Qk	s�rkihH�ߝ���_��o�bv�tG�"���~��j���Ì,�%&��������Mu:�.O�=�]?��#1�fT%�G\���x�i��x�����F~-^l��0���P,#[���|�S�P���J`]�GK�}7d���C"h$]@���8�z {}1Wm�x�I#�ۤ5x���2�3F�D��N�dZ�.���k$��=�_Vs4����a}#��#���.��}O��oC)������e�D7ke�{(B��\�k�j�7��WC��L����t�(����Qw�~��{{�)��J0��d��Aj6d-��o�\�I�iB���͐��� 1��]���dq�����H��3�ۡB��C`2�C��
Ɇ�6��%I��	�J���'�� w�"z��o2�����$���4��%ǶW��:�^#Sj�@�7�}L݈��!�kHlHvg&P:�G =M���_�ȭ��l���a�(�)TI=���6>�=~�˄���a��+V�l8E�-@�D\[D4��i?~k����]�����
���(��@G��.���Zj�V4�A�jO��VN����$>D�'N�����_U?�vpH�s�H�p�]��u:�C���@��Cf���u�Ћ�������&�2;�AH�[l=u�ckS�QC����M%�������ȋ<�1y��U�U��ja�^؁vG��D��f�u�K���(ՙ����m�C��º�~�������������y���%1��d������R{P��>��X]�B��G�^_~�{MA?9&��RU��Pc�^��.s�b�ݦ�$, �O T��t�����4�AS?~�j���{��']%�G�@�Fg��%�W�x=9Z�����\��*��_1���+�@P�C;Ks�5>+�$��Z���&H���[�4�}�﷧ ��}��\�ҺD��p@m|���Ǻ����ɦ�7V=�)��*�;qQ��"E���ĊF���B��d�ڢ��n\E�Qx���>86 ����H��;"�pVV��?��q�Ӱ������Φz��1�����A�h��D��ǀz`~.���1wzM-0d�#�bQn�C1�^�7�r�Sx��;C?�@45Э��ϩ;�߈)���@���D 9-���<��"����c���"��y�i�	"�����a���D��K���ȵ។��R����o�̸D~�-k+gO0�欋���!@ė��3Pɞ	���l$�����M�;��P�&��E�f��^f���k�Hq��@Լ�4_5۫x!�jX�UHR�U)�)���. 	�D2H��ӡA�Eߕ~��S�4������W:{�/I�w�$����c"��lQ�?�Pĺ2�!�!�7�m���D:X�Ԩ�`@<{�|��g�-�핉n_�V�?���L���{���3ӎ7�
f	�½}Kc=�8hߞ��>^:�0�WʩӀ�wg2}�y%� ��k}�3���@GCO| |��`���l��(�y�J��Xŝ�8t���F���� W��=��)��6�`�|
e�0����������94`��c]�`ra+�+rB�3Xb��
�u�X���u,U_s��U��I���%1A�\i|�V�;:�r+d���Հ7�Ö�\��u劆[�g饇�}.zA��%�t��SW[�hB��_5M�2-��"���:��j���PJ١�0��K����I��h`9�w�ȁ�������:�M���1ԕ��i17`*�x��^v����i;����cB$F֬j)�-�Hɓ�^�M��CN�A$�N5�{ޫ{�mNLRsܶ#NX6]x8ݔ']Z��/�������1��r�D�V�^�A�N����o��Gg��M���ϋ̷���G��\�Քqa�0i�kj�
�C�Y����=�-mP�����w�PV�A"�;��HC����R���ƾ��.��k�OugN'fA<{X�<S�`ϭ�#��9�P)u�)p4�'"�hApS7���L)��P��G�.�Z��NV�Rn��κx���y��Eu���z��M�X�a�U���ωQ�G��ٮ��/����Z.)P���{K�ȻQF:XաMP�r�s�r�N��H��]��#�����p��.Y�����D�{�d#��D�N�+<;4"������Q�k43_�}�-�Gҫm��%������_;������u=_1��/gldqpS��G��.WIg.��}Ǹ�Ԋ��o|�JYx5o�5����#*RZ��4�EW~��Ŋ��!��rܵ�
��rs�cwR�e�y�aKK�&���F\GA�Ek	>*������ FJy���Cs΅t���1ד�e�vt�x���?�mb\�x����43h��X��=t􍯇R羻=�o�R���O=�B) ��Ngq�l��r�z{�l_m�	YA�e{�@"�VUfR�C,��Q(�3��.�+�d���Q��d�/w�x�e�{DUO���}��������E�#�fc=!���ϭr�N�.?�H��3<*˾2�0#��>��Q�Q$?T�<^�,$�[��аЦO;�xǁY&fAL{�����.OH�s]�F�lWZd�:7�T
�S2�`��+Nx�׍s��jծI�����dG���L/���#�*x�#��k�g;k_��ͯ�t8HX]��[��zҋ;gj�^ڥ�Xd��s[<	���R煶��u0�9&�M���Q����\s������b���!J<p�o��|�"�����6�4gx ���׽��MQ�c;Q=P� H+>���M�yԉ�l���������3%iaC'��J'g�xՈ���)�77���j:Ҁ�M �����H�뿽k9�j$��7h�W�}�0B"�-�t���I0f�P,�7���Ti�X�i'��A
V�:�bRY��S��18��V[�M��n�o2�2F��6��}hR��s����	���.FGT���,Ԃ�%x�z�v̝K,KF�Z��*�}é���@�,���XG�HS,��1��1Ya5�:Ǯs8Rַ@����y|N�X�/x��><˫1�u�$n��r(.���1���6�2��j�b@)�gF�z��g���ru��A/�g�li���w2��|ic� ��\Gď.ֱΩk4��Ĺ3Q���{M�֬�GoE�R¼�٪�����uj �FV5q��AW/g�z2��o3��G��-����.22f#�t�UNMw��ц#�Da6�D��3�g���"4x!N�J���Sp�Q���K�R�Ƒ��D����"
�j��Ir�K5'��P���n���C�i��a8�ɘb�kirӹγT˘�;�l���*G{� !��w�CQ�l�A�_�Q>
�a��x4�ה�
k�RP�2*S�'e:2��?�hMs���"����fw}{�h4Ho&��A���FĶ|����Y
قy��xQz���Q�.'�����
����ϔ�ҁ��p��z<ap���k.�1�☙v4�d�˞�Ql/�ԫh>�}�\/�K�x�6��Hp�� ��}~�P��9�l)�r���ϯ��(!F��:sX��tZ2���F�>̄͵���޵�{��}��*�˞d�T(hl�n�;E����xBH�8�h�v�`ߕؼ@,�V3�n����5ʿ��B��b N����	�ܷqC�~���k�i������m 1Uq��Q˪�@YN�N���������<^^ӛ^��@������C���;�͏��ݢ��V{(MㄡJ��YjZAi�3�H��D`�׿�a� ���S֕�B/�!M=��-�{�l�݃Fn4'�Z-N�]�X���l<�?Q��t�����01BI�[���_C��HMT���E�:��6��_c�����"�=�痝�煙r��/]��3� X���H�w�p�0�銥x��>	�����ꔢ���[ŏ�a�GS����XyJ]ދ �� 3ϙ�a�B�Aug��s jz�rQ�#B���N�پ�e�2Ք�
˭ѝ�1������vba�{�t�H���� w� $�MՀ����)6�v��vd�.Zq)n��ēi�ݙ|��&�z�tktL� ���s5�I�Q�@?��/O$�zaj���L҂Eݠ:�����Pݳ!��l�e�����G5���[g>2���T�����*��J��h�K��p��"�\�����+:7�b���F�s��`�K�G���h��mT��21������:O���$����ן�L��v�*���<߷��)6��5! ?��aꀗcL�1AO1~	Ԉ�)�O��NH� @l�ԋAW�� ��ܨ�g��n�Tu	^����&������Fe�X�����1�b�� �(�R8���c� ��Kl\r�N�?;�N��z³��Z��KQ@�g��pUp@چ���hdo�QEZ=Q�+#�q�ܑ*�3�5�n�H�cf}�w��;�˜�2��V���=�j�W�/%h��$s�?�y�V��sXחL��_��+�����~u���,���L��df2<����p[�	/?�آ�@��L��_˟�&G��C�����	a�!j,�i%���R���{De_Z8>��`��^0�w�9���+|�,+���z8�u �H@]r�oP8�".uӯ��b��������W��l�Ω��S�M�r��)pU��Ӝ��_頋@�ʂ^���p�&f�63���/[��	!x����)^l����ܧ,� �m~��ğ�gY���Yx��Ʈ^��sQy�:�Y_���'�83A�K�`=1%��@�[��~;-�93Ɠ:y;>;���ʂc�f����v%R��=O�1��m�s,��	\#����z�'ӂ-NK��7�n��Q@��@O!�O�?��D��Ӱ'�Jx�.��|��m�&���Q+����om7v�snk��ɺf�˜x��!�}jO+z�WVlU(���kH�}Lc�܋�mw;1�ȍT�NH�阓�L����G|�m�'�t�J���;�l8�0�6������"(�'j��� Ѩ\	��IU�3L���P�d���ws��c뽎٦�
��f�֢��m�e$t]2�3��hb��0<=x���B��a���NB�9��=���"�m�D�\��%���vW�)v�.�¶�����-xՓ]�<~g��c��kЉ�(�$�8Ɯ�?�6�l������ʉ5A ���z�	�^��u0�J}���0���%_�@[�Q'���)w�V�z�X�jD���[8җ��"s���=_c,;hΘ&DT�e|�ػ�0A�:�8��N%qꋱ\Q�=��1�S�
y�������n�C5+���MVXjc������۔�GV�c��Gv�S��b�� #�Y�Hf�8�s,q���A���s>o!�L���&4�hI�S]�HNw�@�[�
'���\�Z��Q��{�6�M�3b�빲Z�Z�i������:��F~y�<����dk�K���l�v��Ǟ6}�Ӽ����|��q�D�?��>�(żnqg�ˮ$��9F�1��&�헚y���ɠ61/W��L�^�Xg�?���w��kh���p~����!�֞'�������%�P��Z�a�%w�Ӟ9�bP�-]7p����
K��D�?�O��u��ՙ��(�i��~�J�6#�ڹ>91�UF���T@8Z�KX��kL{�q,o��iqkM#��f��;旄�a��Z۠Ju79�W�R�Z�3p��P�#ؾ����FHM��z��:k���1��*8T��R�֟R"}��\w�����oх煲W�.��=�R� �b�9G�'�q���F�xR	9p:Q����3G��� ��p��5�
�p���
��"'zm��}^�}b>:AYGB���m'��z���zP�T�R$N\�(Μy�a�Mxϭ˕����R���|�.h�����Z ���R����@z��o�0��Q��Dk�� \��N�����bp/��slw���f��EN��)g����O��u��Uޒ�mmR�����)�5��9!��U���Ϟ���WV��ŧ�=�X��
H����г�̙9S�h���w˥�^HPb�1�J,yڧ�ÿ��J��=�r��P�eHս��p�
�e�����^��X�N���zB�[>��y�������ǡ�K�0�	L�6Bs(�p	��z�oY@g���a�էp8M�DW��q�{W&� ����t��;"<��v���6nU�'i�wp�y� W��C�G���r��/�a�%��I0�*Hm �eX�Og�������y��.`�H��1�j>5.���s{��`�L���SL�c�Y�kv~�G�2=���Wx�	�;D�*�`�j�,E�>z��}�D����0��8��x�S�]&��/�G��\U�ھ�c����l��o:&,<uХ�����D��&usTR�b�@u���Ho�O{�\���U^���l�Z�$҄�v����9]�$MR׿��F�yc�a�� g�<~��[^fD�C��t�x�� +������d nT��Y�e󅴠���:����H6����L$4��^!H���Pp&�w��͢��Z��/m#.|
:tZs�� %��p=��f<M
0��O��
-Q�F1��V�����#p�|�zE��R�o�x��}&Eh��ƌEV-O���όQ��;��0�:��N���X��۹2�J:�
Ҳ�4���)S�^Qk��/���9B"�BYFB�R��]���o.�<-	�"hea<?o��#F6ط�JJA���m�B5�; ���J}��Oo*A�f;���j�9�Q�\��\�U�k_�By��\d_9`t&*�|>�
��>�i����j�
TWt�h�����cO�'��W��;�Hʅ�DJd���_�2�� ������j
�桇��D�`Ip�Ȉ�����zIK�I9b�݌��� ���W@m�Ew�TH��!*7��aO��C;�}��M�z�/���;ٜ �,�LW��� 9
�.E�M�x.b�����}&������'t��L9D]iu0dnf#�YJ��z0G�k��;�)�_[Ap�[b��@��YU��:�H��zϓ4�e��.%m��/��9��&W0�@q��.���;���|2�;�;��f�R�]���f��R�����>k�R9; n�d'UU�	]BF�,6�ꇰG:�7�Qj�L����ŋX�g����b*s������.��@*���7ߊ����׶D(E0��v�"�;�ڹ�{XTHY�)b=��a��O+; ���j����d�<Z@ �dT�F���ܮ'�M�XHjNC�S{��0��>Q��a-��P�5��p�ƻ/�_ �Y��T�<���W�={��RƖ3A����Vv�4nʗD߽F��S�VB����lq�%��� ck
�`��c"њ�n�N �so,�u���lhJxH���y�49"�;��%�:!t�f�}��3�d 6 ]��d�e��T��Z�c�-MZ�}"�X��S��s ��W���r"�U|�i��[@4��H��D�����,%0]"���O.�雩��jH��%�@eb�̚mʥ�RX�gX�Ƥ� v៽�g�Fl�����{;8��R��)�+ �/Rl͋�i��rGiEF��y�Kڻ&�q� ,˕ ���@��Ԏ��7�%�o��!���1�;Zrl��d�ϕs�kk�Q7kH��c�Nb�YV�v�WG�_���)�%��H���@�)���*��N������oi�N�{�$�E��vH�������
�������7�:WI��uDi�l�+�ȍY�iy!g�Ʌ�|���b +�]���!Z�/q7����&���?�X�.k�n�%�A�I���f]56�Ŋ6{��u##Vw�5�ڟn#;4r��j�2�[�_J�Xʎ��$�v1�2J��u���$T��: wҟ����w�W��I�i%���	b���� Ka���G|jx	Kxn�M�$*�hJ�F������:��B��H�'-����a���G>ڗ��u5���������)�S����]��<\�}[�V0�V�sg����~�\��39�ŕ(�ϵ U�k���V��T�7_�� �%w'8��2��i*&��^�1O��]��n��]մ���B���l*`�N&̩o�Y�\=	k`�Nc��S���3j�9n�s�ڊ���ɚe��s�$Ӵ蛳��  ϝ�`d1 ��)�UE	�1�([#@��1��T� %3&���+=v����Ǉ?Glg$ȁ�]�[PӃU5V����1-;���>��D�lkj�ԃ�u�� e���8S �E�a�S��j>���T&|dwf�: ̧J;@����yY��_��q�|��5��c.�yZ�p~7�����6��s ��Q*�&J�gj���-4��Wx��)��Pp^<S�{<ط��DM*���ǧ.sN6Xr�v�w� �rsh�����)�=������,��l@���!��q,-�#ds�Gۨ�����g�*ܞs[�ںy
��}��C��:������Q ��Qh.-.V�Q��hB��5E���\`C�ڥ��^P�yb�ҷC}gG�^t�
hq�=��}���ם�������c�)��?�B���z���������U�[�`y����Ƈ����7,�C�g����^q!m焘�}�¾�=?](����]�"G�ҥ�h,>p���2�@������y2Z���~���m(�wO������c�k���xo_-��He�Ԁ�X�w�BnW�T��S�Zu�v*!�����f����Y�Y�N%ߩel_��&�W�vY�����r9Ky�ɐ��[k��r����ͩ_¥����L�C�G��)���k&{��AvW�!Vhe��������u-�􄑔�dob�&_]ݕ�8�K�'�{�Xz�o}�g��({M��RyX�=�� ΃����it�v L��R3C>�\q��α���&�)���<���vy����9��''���<�Z2�w���P٠W�%b^i�άH"��V���
�.t����0E8z�t��Td�YTǲ��u4a$���9�󖊌��e���Bnr�h2���8Eeѯ�H��	�sF20�n�����쵭�qss���"����V�#-���@=j�Q�@JE��	,w��WGP����%�c��,\>�m�v�fآ�b�s�g�TN s�=�� .�H#|��#��?Cw`�h��c=����߼����z���OE�M�lo[I�����=)H�Y���/:d������]=��W):��(1�98 n�͸6"�j����e����&�9�5��`&�>`��9�_���D���"��zY��W��)5R⡎<z5>0JOD|�7n��0�0Ok�{����XT��Y�A��.f�T����t��?���Ef3��~J�,����ܥ��&�c��I>䬛IR�ǉ᩽�Z�JX��6�ʂx�h�m�����E���u��<�B�����TDI�\�.�A�T��or�m7�@=@�����s�L�����ʶ�b#��*�������� )�/4j!O\zēM6p9*bЉ:��#o�����9���&#�Z+tt���2��v�,�8���ۘ��	�Uի��������{�YV�0j�����ޢ=H�u�g����S�P��S�[{J�;ly`
�:@ڲt»OTN
����4Z�K�wK�]��7-�a:%~fh@K%�kd>�!��Uz�Ѱ,�k�%�Ͻ��5y�������`��p�`���� 	��C�/���h�!D��n�P2+�J�C�Q�=Rj��B��iV<�P�S %�:�?zH��M�*���;־K�~@C��b����>�B�Jz����l��}b�~����^�����J�S�?4d܀�����4�_��N�B'�3�6m`������8�,N��9
FW�(T"E1�I*�yC��&��
<�P)
����e�L���N�M��C���~G���D�c���HrH��,Z��z�c��{E`c�{���Т�tm��Ly݀jO����~=K�X5�	�d��)ɇj����D�3.3^�+�SR�]߈��\�*_b�g����@nh��lh���_��/�{N _�"�����5#Q�4,�}\�� �(�L!gL1��<��e+���1�)	��ƨ��Sp��� �be���yy!�}��5�Л4?G�� 	.ۚ_p�,8@	�x�e8�EƻF�t6���RsSa�ُ�[J��i̡2q�9Su�yW��0[�.eb��-\��CW�����&L+�^�J�=�`rO9pn�l�����2�V�5����wi�f�v��{���y��UZ5�%|��ECy/�>8�+�(��q]v��Y}{̯D2���뙔>HA
���!�́M��ȃ�{�8XF�ka���4�^����2aM)�
�ǔ�N�*GH����ez����/�8z@1��~|��h�F�Ap��Eߪ�7fU ��ɏ���"�&�=�����Ө��L.��?����
�ń�@q��˒�����h��,���HőXp,���(�=J��[��������c����
��%�zc�%M'�o����d�n/m`�ʈl����-輘�kS�˜ɗ�Ƅ��f�l����_D��Vÿa0,\��%$����ToNk��Y�{���'�8xl���`ВPR<dr(��?䯑�fj���y����9
�jE6�m�H0�p�51��ie��$ @��lm��ԫc�K�y��6��!�c���[2��i�n-���8�#�����j�c3��g.��<bE�e&�식b�f`������m���O���>�.��:w�"Ռ#܍����K�N����i�#H` �WȨ�+��P�c%�_�0C����l��	����D�?��*P�Q��� �0���d�~-h1���S�L~R�w3gz7R0�г0�Vv���Ԙ?�K<[�-��p�)�:0:7�65����oI#g��/D͑�m5�� �A�\�SE���Š���,@3k����Bڴ�I��;T>eBg�H����?�?���5���4���6Z_���~I��.�_|���Z�o�%9���9o�bR�� ���q ��2��T-�����4�����扂����{^�2���C��-l�[��F�@�.��[������`�&l� ���Z�A�1\�ќl�B^�W�7���W�[D�<q��!�ѵ�u�_�`��ׁ~~>ٯ�E$���R�Z!vVO3jo����7�]a����q���Te��d����Jy��gj�8�<q���Ϲ�T<.V�FƷ��I޻B���0�×l8���݅����>��f쯃�?�"�Ƈ��H� �(�{d����A�m�T}�ώ�R*d>9F�k�Ѭ�5>hs��1�]EnhX���U"}�Q� �ڃ���a����� �]�/����Ij���U��'�(b��Z�QQk,^ש*x��[��~r6����G�y�c���K��ݭTB���z,�e���U�w�������M�#��7z����i_�'����N�����$
�$��f�̟�p���-�PH(������;�� R�-����.{�*t^8���f]�s �}'���6���t��m���p��3�?�DRZG,�Q%zT���-��o�Q#	�X�r#;�wkSo7;c�<b�'��k�9f���Kb�K��)2i���������S��9M��7�>��*W�|�O� �=r�s�����t欽�b���t�N�I��@�/b���%X<�����*�~�"�s�r��߇L�qP�cO���7�qyJ'}�"�KP<h��ǒ�,�]��MeB�P.����9*���ɟ�p�Y��GTj)�t�I/kfۣ,�+�"LYC���g�2� b�=����rV�ҟ�d���e��wB�ߥ��E�T���1�?1�b���[T�r�^�șv}��Яa���4�E��ib� �x��P��t��] �5��£�دC��ґ�Mr���C�{��`{>�^_����Ja�!o	��9��ќ�m���4�S��<b�Rm�C��o�����^u�u럎�Z�F�ý��M�$ ;���ͤ��*������i���"o�!�3XI����`6,5>\�������LJ��gc6�ki:�k�/�t���L���˵(�zH�o�_�BzՓ�2q �ώ���}�ů��P���'��--��evsG�hh�������Җu�nip�I�Q�k�=�i�rFb!Uw�;�p�VV(�ywe5X�Ѯ~�;v����n:};:��E�K�w��c�=���9����p|�p�GB`,���{^��8�Z�.Sx۩L�)�a��k%�����\��	Ƌ�Ӣ�Z^����F�o�$��[��Emލ���y����1-w�N0����1r��*ڴ���TjJ��������߭�D�^�m��;�2���Sz��䄛�}��_�
��	��Iߏ�9x�"��<���w�Rm`G(K�3�]R���)@=���j���QliwU_q-Uj��	�ּc6"���0��1��2���1I�[����z��g��LPǩZ�Ȁl�i�1Xrn6`ujD�]M�xd�|�3c�����C��+�]~�S�=}B�WI.T�D�ѥ
jf�������z�>&e��c�����8�N��f�Y�L��&�n©��mk�	^�`O� j7˭ԋ����PsFi����Ѕ���6���2��<])��ĴSUـ7�nަ:D���<���@�d�6P���kl���w(Q F��M�H���30��#�-ά��7�n����;�1��{5�E��q�+O����g� �T� $IG>D�(ܿ_����.��1w��Sd��\-Ռ�{�Z��g�?�폄6�q�*�yq}��<Q^XV#�����sU��#�X��$O�S?���c/�{�"�vU�J��Vp���[&}4$)��f����ns	����מl�9���Ǫ`	�n�nN:xؙ6����bPbr_-Pw�'�V>G�NS�~h��o����r����A9r�Uƒ������s��)��~W�u[���:^f�a��)yp82�N�e� �x��\ߩ�b�3�+z	�R'�����X��&�S�������$�r8~���4ڶy����rI��u��>֙�ǌ�8i���QH#=:.[Lwd�~��I|�j��"#��?�4%�����;#'>zBI�nj �A9�����86��7B}50V!��I1ۯ�ɊH|!�"������T�Պ/���'�{z8�TI����{kH<�������?�-s�ĩs%�ú����H�_՞AU��ffI�W�B0n�����!J�]1|��/;,oK�1�/O��\�f��]w���K�Y 4Tws����Ǩ�hv@u�1�i9���]���L	�T��JH]ڍTI�w����KE��/�{��]��-b8.��N'ُ�߳�~��5s�n#����^fgɌd
g�q�
�<�n���)�	mW?��]�	���l��Zt��r���U�ĉ�P��EH��:Ȫ�]������ѭ���`�"��ff�S��H�6޸�g�V�3��)g�/P>퇹�%8��̈W��vÅYb�Q �U��E������9��l�+�k�X��De����y�UQ9yY�C����]��o�#�
I����2JQǖm��}ȼw~�ԉP�Bl$:?rKZ�bIf�h��C
�Z
?1MIsR����@/�C�pbc�o_˟�[��w<o������+~>Vuݬ�bHq-y��-�@���ĕ��V�m�O_؏��$�&��PuC�OѢ>[i,8ȟ����߹�21�P<9?��~�����A�$0�crY�������r��)�R��0$IR3�'���n�2c���4�Q�*�v	E�F_��Ӛ{۷������`oz?eb�����0��A���is8�ټf��J�� ӆ�0>�,���m	Ŵ�,�G�\�a��|�̠s��$�f���PN���KHK�	8�o�(� j�4!A�ioD���~�s�;j��Iv�͚8�L@�a+�.S�V��`x��c]���>C4]R�nњr�� ��dC˙��Y��>��%�PxV�[�0in����a�ZD��@�J���[��5�˒�ʻ@�y��E���+���l�oj�ʘ5?L%���Ć��7B�	��)c�����;��C��z�<�i�.0��MO(h&�A;u�a��I��J+�W7����qʐn��^/jM�(Z�����-�w�5ь���)v���쬸��\��1=z�0u�o.9�tsr~�(����m���}�g�I�5� �3ҖwK�\�`�n��\T�.,��{��.��#�'֐w���3�Phl��贈H��՝Z�:u��QN��P}-�oe3���w�L;���Ѻ�_(�7�Y+A�u�8S�]jc����<�w�e?�>m�,��Ն�o��Ȅ?(���3.�y��5�Uwh����$��#�%8�!N��D}������<�JA��5]��'�1�H��}�}�ݟ���5YW贑��W&�#�!:j���1���iƲ�0�U��}�1f�y��<��&���f�w��S��-1�� �F�&n1&@,u�%�Q���*�WO�+�����fƮ�#����0��x�&B��?YK�9�G�"��H��Ǐ�sFTW6�놀���sN�AS