��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��s������\�Ἡl-�y�f�����f� �ѕ:�nA�kb-q��_���ѹ(4�dê*���7��N2�ɐ��+ٞ�4Y6Mx�ejǴ�y9�����=���D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6��\\�l�����r9s��@'�k~�{�<���y�#���i6`#Ɉh:^[����*`��Z��|���z���N?`q_���ר�Z���FLe���Et *�mk��:�2�|��S��1�L{��:�;��?)��/os����$I�G��S�Y�a�.ڌ �|\�E�7��RH�����w[��`�d@�<�S�쇦��y~����췔ڤ�8��p�%M� �;�.?���EJߒ=6���o7jr����SG�C��,��)������ݍ,�aj�� m?N�L趎�i�eb�>��Æ��򲃁Z�7�	E�͓��rH�s�&��7��_��
e�F��H���)�W�g�l���[��燸TɆҭ�V�{�Σ��G�kx(�}L}j��"���*���A������s!ɑt�`z��t�ۣ@��� �f�wA�4��A2��rx�Y���C+���:Ѿ	w��i���5p�-�� ��Q�tMd�ei�oX:���}�\�C �\o�r��Dr�����dF��]�t���+�!��D�Kw 3�ػ-]ų^��g���������)X����Q��zo�c����*���ݍ��[���� �6<u��m������p�T��K�Q;IL��G�ߛĔk�������K^����Hź+l�O�[�	���tb)l��\�J%�NPM�N��J��Dh������z��{�{�j�p��U����5�2�%5����O���~h����RʗDZ�$A��#_��5/�O��w�ŌC�=���_���2�Ի��pŗ@�{J��JP��>O׼4��e�����w�+�z��jr����;Xi�/�w�p�h"��ġ<h-���d��`����P�t��R:޾$����B�L�w]9
5���he|����Y��i��
uz�h"����g��
���i-_0�p-*�������	�6旲k+�F�Q�S�6[���E�pl�۸p���YP�*#���z�(�S��u@��f�6��W�n'����g�K���3���Fm&C*�ҡ���I�nJK;�{��W��a�"4|�ND��B������M�?t�妹x�%ކ��d�e�0����zɍĐ?Zqs���x�KȣУM=�����~Υ{,����UV��j���g �ڈ�sh�Y5�ͽ���p�~�����W��	��6\T((�C��"rȪM� t^n��X:N���Y�*�1�k�ӗ����E�jds���6R]f`�����t�L>��4W������ʲy9X�M��ciw�`�Q!�#�nx�:c�m	Yr]�����eb;q]��Ǧg)�@�=]�(h�������{�.g2ؽmy�<R�R�&J�E�TN��h>N� ��\�������V���Yn��u1�[V���=�a;��If�һ�R`�t�q�}�X��&�F�ʈ��L��:���	D�a�����.�p�{&�N$��'�aǖ��Ѯ�"�΀X���y�6')� �دK%����)9�a��ۡ���5t�!]���S (���XH_@I��ߓ��K�7���7wy���y~�H�!�V�v�h�y~�޳8�U���iG㸥�f�%E�ʳZs��C��<c6�@_�b��i8��>�G�Ҩ6�5پI�S�� =����j�;�gC89/�X+�Eq����=$��d��y����;�N�i��l�����v_V�@����^瘏���*��x��>C֪XȂ���G�1�Vb�x��.]ی�r�K������?�s�ٻ�!˶��Ľ��u�)(@"h-��-D0�$��'�8>��	�H���0K�|��"~i�\Yx�ڦW)�����jO�z�hn��`qGۘ���+�Ǖ�j�_t����E�1}�}L�j�ePOF��?�'
Z�enH#���t�%�#�O��8����B�P�Ϙ���I�p�E�m��%��l��">1��?#Q3��qie%��6T�y�
R[�0Ez�V��a��e��n�Z��8�")���fi����
����>\���%��2_��D�:�3'���m�*�y�Xb}��g�����������M&�6�,(��~W7����k˯��e�8�o��]��o�S4��U����P V�Nw&2��q�):<'i쀼�4���5T�䴋[+,�K�p&�ގl����?XRd�P��^�^u�Ov`���J>c}m�yT=�C����G�h��L�\줦��#�i]����~�x���$+(xv[;(/Q�8d_s}Gv�Ĭ>��+"����`��+�uC#S+�omnWsA�4����S16�.��9ጡ���BqQ1�]�\�A8��gB�?�th8��Y/��5���F
̭�e�쭑���Qd�eWަEݸ��Z-՟�<�{�3��
Ʋ�Z��dRHb�	�M.׌^#�����I�2�+���DJ��qr����-e��&A?5L;�iF�%k⯿��1�G���_���:�g3֜K`�_�F⹦�MÚ���!RWB)s^�8��<!�`��R�8��;Ƈ�� d��Nh�ƃj����H^H��°
2qn��
#�Lԁ�^���5O.~N
Gi��v�,:�vȨ�wa��$��"<2��d	�4��T�2�^�y�������+����Au�¦�U
+��$I�˺b�K]�r�˔!�����tM�q:<fQ�������]�����jV�#|;` n}c�� r��{8��d��}`pU���!3�|)���9�'��98Θ��o?�u�_��67T��yZ���6SK������CC��;�鼍���E�T�˫0Q��G{V)�����6�ۭe��dN�;FzWf�ZLX�Wm�|�/x�y��Ij��Ҁ�.��g��ݜ��9%�g�:Ǝt*v�;)���~hJ�M�x�婖����M��,�H�W	S�_U���S�� ���H�W����o���n#��ܽ�.���n�7>7�f4�(���H��B����I�\!_B�˨��nݜ��_���[��\XXGq��ea+�������89��� {����/�)�74 ��9nM��5���'b!�5��~[b���t�,e ����&:�B�>z�H}Y�YHW?GI�V,WJN�n;i�������du噪��E@R��X>��./i����% ^�uw�2-����`,���\r^�R��;�K���M��/�8�J��= ��A����^�����O�ϕ��X������с�ԇ��dI��c}�yVp'}�����w;�@��<��3�0U���SK-�gd_v��Ec>ƚ���7T]$�Q��I"[�㭬P�#.�S��^��}<�
$�����K߫�=�dT��i�i��e
W����۱y��$AVXr�һ��`�?��^7�5`q�}t��w�+�E��bkC�g��Qƌ\N��xnJ!�;�k2����/���Qv~�x���hPU�7gs�!�y�0 ���{P�~�L�����mp���R��C(��?�:3��O�8h�>E�%"��2���)�_��A��X#�_�� #."�k���:X,»AT�Q%]S�����h���B��)w��F:!�l�x�ԭ ��1�i��E���а�)�0eHoe3�aȣ�m�)
�z�x�f{�⺅�Ƹ���WQ�Y�t�@X�|���_4�ھp�(2#��Xʋ�L���j��A8�K��i��3� G=n���l#�H����x����Ht!�xQ=?��~�{bf��vv �ƶ#Q_/��R-%��8�+���~C�\���w���6��eViN\�.���<@k��h����]Ɗ��GbW�����Td� ���6p��?l��Q�C��.N4U���ҧ�ٟ?���[l���w�9�i<��SL�R�2��L8k;h^v�m1u47%�S�/v�ث6B���9$6�ߕ-쨺T��g8h�jӊ#)k���,v�>q[_�b�4������ݚ�|-u
d�h��"@[�/�J��dFGM� z��8�n˙�o&�1f!ٓ�}e��(�@�����c�A�~�t�e0��g�Ad�l� �@Z����iL���o��I��:�u���r
�[<\?ƿe{�O�r���&��D��:�����dٻ���SVd�{��B��k�nqθ�Fur��5�W��՗��E0���ۄG��p��	3XI�������ViKb��~��BY�ñ���n�8ݱ��=��:P��O���'O��El��@�G)�1��/��'��#�J݌��� X����q���u��At7&�S��H�nI1� Z����.8������K�D�C ʹ|,`x~$L��Վ��{�����ħ�R�lh�=����:h��-�$�"S��_� F \E����H�q�������(cmyhҫ�&���AfRs-��i�C�����"�P��k$������b��.'��7G�܋����Ă�������8AD~Fy ��w��ܧ\\�ח��"���~:�o�ܴ�!E��ؑWdI_��2V���+�HO $Q�Jv�Ƭ�[���rȮ��v��L�|���ٍ��v۪��l�,����+�$��W�^� `�M~��Ǔq�$�z1��ۃ�>�Z5ܿ�f��f6O+HU^�!���X����rsf�����@!���L�������=�V{,��T�������7��Ӵ�[	wp�v�Y��<�W�Ƞ���l�2�P����@�~#r�瞏ǉ�� ��xav��om����P8*��_ЂJdP�U�*O��͢H���|J��`���t(��҇v�v^�ت6��h_���ځ�����x����C�dd��sE��af0��f*N�����NmpF1�삳Pd���W��	L��|��F�W"/��eP�����i,�ʜ�b���C�Si�*m>��(��&�y��<G��:�ɀ�h�m�g���z"�� ���c���A�?�
�K,j=�T~�vI�b��6�1*	�ڶ���ȳʒ�
ˇ��?���to��#�i���1Q����V��a���_�Ɍ��Y���e;���)���y���OzϜqn�)��R��~��It�t/�J�x#��(h��D��}�9iOS:��:�-����-�\�(�px̳����Lܗ��ƙ(��0�ԡs`F*�a���n�!^�^P�z(D����j���(g�₍6����B��Ǻk|����G�s���gc}R����P�r �.�*:�&n���k34����������Z��d��2�ߒ����p��rXr�F�4f�H�ťWmz �/�%X,zd��8%7�x�V�.ɕ@��2Q� �~����qT�H؃�0�Xg�{MYzl�YS�8�$���6�B!b��C�Vk;0/VE@��¸�r��b�|ݜx�8��Fr�[�&�m�2*?S�]��k%.��_��2y xc���E���V?\�� ���5�iQ=��� @�q��B���N��U0������^r�k�����CP8[<�p���0%j|��9򱡳�5�#u�$���+����7�����vŵ�C=��/"
�@.�,�5�s������-9(-�b�����`�\l��}�Q{�Jr �x�yBx	���[�H��cg��<tm�<M~�z��q$���nǚؘ7�V�k.��q,��o�s �K�_�nW~�;ԫY��AT� ����)+]��� q_���l��� 2k�g����}Q���)/��������va7��rt��J����f�"ZN�:�n�v�&�h��3:W@"�>�VcR�ɕ�rd`3��%9�?%��H��I�s�Ѥ7}5��ۙ9�q������g�ꣲ��׿��!�Kt�n��§P)8�-|���D�巅����� �sm�)6�X�!��.A�p9���\�⯮�ZB�����&���X?��5]m�����0p�h�f�%9vp�Q�AE�C[檻;A�B��Юu�( �%�L*Í�gPY�UT�����b�z���fa҆��S�t���W&>(c�/�x�zD��u@�l�^�>������R�b�7����)��\�Fa�k�m[�y�͉����.��x�D��M���ێH�����sn����0��|H�/�>�/Ī��V5�����LC-�J������N�v*�#q�l�&0�;�z�z�p���vbq�D��J������xr����>�8�� {��M���5��-�rL1#-�vܗ<��ý�&6:'�s9~��C�[*2���S}Os(��"�E�{��9��2ZV�o&��6�
-�a�țd�|�ֳ��JyrB�B٪�׉���3��Z�x�M�E������/��-��	ڛ x��a�Vx�'�ȟ�G�8ڋ�XCI�T��
+	Jń�-\�hm��z���L8����;'��ųka����3�nC���)��\&X�gv���CK_E,�dy����� ԔG`4=��N�4ǀ�2�*-IN��sS���m`���P'ۧ���W�~��������ư��-'�EM�0�^��a��r�����M�\�DL�&����΢��+�s(A�m���/4�7�\�E4�e^�rʳM	�I=/`e����L ���aa�����q�a^��&��3*�Y���CsK����+،�N����
�ų�tZ�$�Zǂ�����<����v�3�������iž��s�+�9�>n?kD�9�EI�f�?���_�(�ŚS~��nu�<%��-x\����_Z��+���@��w[��ײ.�~3|$�ª#��5	;��[Z߉��ߏ��@̅u�e>�S�� �:�W\iҚ+	(�!5S�Bp�1���1"�a��:8��i@�C/��I���͕	l,�F����uКh�I�kor�����-�i1���LEH����[)�к�#�7�5s�5ܖ�
�7�|�������_����M���� ;�唝�8`��l���jY_�6(6z�If���*�� 6���6�AU�C*��+��L��������A��cW�W��2}\�;���HGS48�S��T��_V(����r��t��ݡꆃ~�K`a�q �R�h d�O���i���\��E'���~<e,%��ȵ�+����P�"-�A�@C,�R�[z}U&wG�n�9����~����J0���"�L1���*hcN�QAF�x�U��@D�b�F:!��Z@�uq��Y%"����i�N�L̆
��No$�T��\�����OuU��/����9��5��;�!SB�D���y�<� ��������L�{ZCi5�N���s�mKlH/�X �L�R��}�!JGA��a9�Fƭ�n�7�$`@��Y�-&¡֯n����A�K����"2�%X�i��=�����b��F��{���@7Z���h6&��s|�]�B�J�B:�q^��3:�z���y�t��|���8eBB��a��]�lxq�C����\Ȣ�0p�@����#��J𸕿�[|=VH��Y�J+�u�ס��1�
� ��MX��� ��F�뾮���>sr�o�В����kҒ�/׊-^p���A�ȔG֑X5t��>�U�Q�p>�@��Z�r���A��$j���rM��~�Gzk���N��P@t)����n$������T���]�t��Ho�e獂��UC/��h�N�O��X킐��kc�M��|'�Ypc�'�:�U�՞�� Ma�!:��{�K[�6��9�0DB���Lw� ���6L�C�'�j�>/�&��CT��)�N6������П!L�3u�7������ߵ朮��1�c��hQ�^��sY'	�G�/��wn��t5P��޻gk}?e�/�5�{坤��iQ�aƲ�UN2�t��	^a�R_�9pHd��Ƃg�1�%C��Ꜧ�A�TO�es!�A��ە!���3z�,2��ܓ	x��u�L��𡖫��!8��A�E
�e�pJ��L'dQ�ӣ������g�K�!�D��-�����@rI�;ђ����
v�z�$@��α�j��6��h��і��_؞�@ߙc�Qh�TO��v���2T"��w��2��89�'����Z3瑤�c�5�6S<_z�J��;]����	@�Z�w�����"�	{����V^�Nɠa����q�;�*Zs���|�]6h]E^Ô�.�on�y6_ܫ|Ǿ#�bq"i�<����?$}�;
�� �o�(y��(w�`J;}�8��/'C���e�m�ƥ����z��L� z��iz�!%s����Z�ٌ�qY)���C,9D�Uvg�Q�⣁��ʢ�d�o_�G��lh��v��,�
�F�o�_�Ձ���ڜ�C��������66�R����^1$��h�QX@�8r���u�@�ׯ��*�XF������T������jSߝ�6���L?up���->l�9��k�O�`�&C�Ϙf.͵{�Do9J�����K��:��Ʋ�䒴�����������	��
����3�����3?�d�,�u9�h��M)z�o^a���b�4�sչz~�z�r�����V�� �X�;��A����`���*�<&1Zz;|y���;ý�W�����4����Y"�;�+98D�`�#�h]������u/�����oWˌ��s�����xif4�YA��Φk��oH�"�́;DVx��3ު��z���YCB/������,�?%x섉L} V�1���%�|a�Ϙ4��.��/�!���C�H�Z6�݋� ����M������C	�R!�������1O����L��q�2��"�S8�k�v2	t(��}��[S�4���#�_��>��hX�w�N��礐��Z�e�C��}�^Z�U��N�F:��������bD�mQ�Ԏ��6i����;��Z$԰`���za޴����l�Ӛ"b6�c4�^��gLVο�z���7]��2M�iW ��oq-	%ą������h��EN4�];�'�@'z<�GH#�Adش��<��S��~�[�A���푚b�y�ɭ�J�*Jfo*M>���l���0?$5u�һ75�5��q�,ܹx��\IG3�;�:�|� �$��1��x@�@�������h�0�e+�M�x8�P\o�j�WPpf֗
���)��x�����D�2�"�n%~�P'���Sw|�����������W����0ߕV}	�;P�����j�x�g��P�=/!�^�o�a�%��0<FY\���N9��q��2^��,�p�i!� ������8�&����Ӏþً扦9��B2��	Q��7�A��g�5#���M�9�!E���SԛR�c�r/����k-�	��6Q��z3Ng�3~@�8��'�8]U�r�p��]�^�5���8���UZc�o]�^�GI6�F��	������Y�bIc��Mo|h�AաA�'���������u3�D�ɴ�2?6��+B�O�W�k������J��3M��{xj��q�*x9L�8M�.U� .�a����nmY8oQ�Nf��9�@�<��j}] �����ą��R���V��%��Q[��S���\1��+ps��;z����y0�d��p�s���.����K=3��T�>�"xtl�4Fc�����ʂ>=P��j���]5f�l�\��܃p~	#�n�r@�������;��<�v�cmv�CA�1���S�I?�$�(l���+z"�B8�6�/�׷.���~�I.��g�G�b�w�:qC���I�Q�1���>-ip�t�����0ì�ۋ0M�����Q�:w��*랃�#�PH猀���ic�p�U\B�ȣ�q�A?3�V�Ǌj��P�!�E υJ�nB7�^�OS�";蓬��ݞq�0Ё��T�@�T�54u���$)��RSom�ǭg���z�p�!"���m�6�eZ;P�2�����B��ϱNԋ�����ܿ�I��jz[/���	<��;N��|��S_�~���%_-�zg��/bq�5;aƬ�qTfF���A�!�[>�7ʏ?�x�9_YH_����Ο����%F^�NHp�p�y!TJ'�V>�D	n��ܷ����o&哋�0�{w�u�h��B0���c���*=N����>;TVD�I�y�g�od�.	
7����"�jʌ`�4G�?���5ٽ?;���5u�>�S;��R����NS,`j�,�HN�h�����hn�������!<Z��[�l��,Kfl���;����/��6�̰ `�@�U ���t��8�x�ѣr
��[m6�J*o��J�'�jE����!�rH�����e4g���)'��#-Qd������{���Ԙ��H�.�h��Y���KF��%���p���ӀƎ [7�A(\��Rgh91�i�����u��$fF^I�Ԍ��I�ux�Ͻ�9��ƽ�w��ؤNS����Av�Lg���G���EG��<�*9�Wo��Ï̈��䊒�$=G03�]�����ۃ?:�eNˎ�~��G)�%�P�&�)#���w]PK�ؖ�ƨ"4�
��r/�FX����C���.s���@�F?���䫬�$	� ��3�,�'�"��T��i��y�X2�V�N��T�UòK����1�*�l�!��qS�*��%o���ɱ�	��NJ�T�Y�)�vT�g,SA�w� ʈ!jV�x�8�o���o�,=f��Ք��,���8�Hk�6�l��bvs�ی8A���*�n[Ϲ�.hS��3��B<��-P��m�[�zEUh���r�$ h�M![�w�m� ŭN\��Q����?S̻��C�V8��I�h�t����n�����]�2����E��n�<^G#��.o ��O�U����T�!��2_Ք�p�}�)r�����&�����ܤc��9q���]�� ��S��3n�����]�ZW����|!�۝�G6 7�[;�AAJ����";嘡 ��-�u�z2V�+OI�58*#���p/���̺̩�R�������o��z�F���[3����Kz9���~p�py�ݠ��6� Z�hӫ�������\m��	���K'<��v̴�y�v��M�ь�*�r"��oW|�/�K���8��4W�P���]��1}mclLŊ���������z���Gs�\�!ނ��P�+yP�d1��:5����!�m.�XS����X�Z��D��r#v�(����1���S�&[�Aaf���Ga�,Ky[[����R�	���S�)zR;U��ex�&r��cYgћHIo�_~Γ�R�+��M���ׄ�>���p=Xew:O}{���fd��4嶯7��1Qm+���i[���IF5�1��9CS�k����E�aC��Bn�t�5砓��-��#G�U����N���H��,W2��앺t���z�"�U�kC���L<��ּ|e�?k�4��Ne �r"���x�y8�㰧n�8}R��+y���,�|G���_��>�P���V��'a�CF���B����<�bӌ��?yx��`�.>�v�0ǵ��i;j�p5w�]��u�l5C*zgY�(��58������k�ө74��O�����m���HG�=9]��ėR�K*�7sv(d�����,��Po�A�ѝ���E���,���
��?f���W�"t�Vgq�o�g�E�����V���'@��@��������Ho+�� y+�5R���Ɩ�>@C�pe&�(aӓʕ'���;"+�O㈍ #�F= ={!m,�zP�"Yy�+���3���	9�&���,䤢�s=��h�eK�OV��؜���A��&�t{�nһ	Gb7<hT�"�\>5��}<r��nуtTq�pź�̻��.r)%pɆ~P��J�&�ɭ��v��؍�z�ZwU�"P�v4-}�7�<V��(-�Qڐ�!u�S�0N�;�1m�怰A��]���K��F�
�#��]�L��d�jI�I��;y ���ϱ3��%*�x۬нr6�5��}�y����Gñ��o�OWx��^"w�v�o���Iu`��d����b�B��3*���{�Ȗ0��}J�t�,E���]M�Ŭu�"�>�b�s��N�~�M����=��b�Ev��P� 	��P��S,���T;ff������VH��W;#���I>��%}U��U{L�"�5��Ƶ��!�)ڳp}*?�QOuaWq���Рw2X��U\Q�G)b?dᣄ++B�y���o��I�X����8�����{��~�[%�y����Ѵ+P�Yj�����5O��	b�=+~���w_-+-y�	��*_*1S<�➭�g|E�ͦ@��T�R45�����0;<&i{]YSei	�:����f�!�}��0
'7O�I��\�r��I���F}n����Lk�Wca+%��n2�X�4b��##��;�~ef�}�`�;����/�%���2���H$9�� \zpr�����D�v-�R��ֶ��%6��F�oLБ�^b[��y4�C9DZT��(Z����PԘ&h����)��59u�7<Ce�]��s�筝(�8��U�N�w����63X�^�7�Han��=��� �*���WM&��"�4N�1�-�ZXx���rX���2�چH�_�JX�Ydb�~wǎ�G���a�����Is҉�1]w���t��L��u�_���������.��Z,ծ�Č>B�&��|���9��H�9�AA9\��	��������9tP<�Wj�ܬ�)U����	T��D�JE��9ڲ!�r��hS3HPL�=�@a�-!�6-��o��F�X�X�\O>�V�7�Q&��E?�>U����@�����l��
[�5�MS��g"/���*ؾ�f>@~�#\x�U�?F��[�@W#j	����hN緡8�K��+�E}�h  &*,��ɑ�R�Ѵrg3��{/Q�L�>S;N*)��|�Ы�Hz$*�����B��]?�2�K�y2�u��I��]�i��\�~&w(_Y��G?�<����eփn
� ���Jnb_UL�"i���
��!�Xs?E|�����u�9q��o��l��t;w�� �����UT��
���T�:�kX�e�e���>6�	['Ɔ�Mq����d�ʾ�ﲉjy����,x|�+�|�@i��7}Uzjv?n����x4�<$��A�=���h`�y�Ԗ��qZEa�IIW65�F]�Pk�+'}�`�f�o�]��͖�ؙ۸!4m���c�3���m�HP�"��X�8��,N���?aO<L�xH(���)��	SѬ�B{����l!���j�k���򗱺pM�� ���j�:��#�����Z�$fKGz��<Z~������t8u���b����pn���1j�I�����E���.������M�4�ʄ�d�`6����]���:0M[;9�v^p��mCo<��߸q4����\S�	�$H%��1��]����]8��Q}l��r��ZG���1\J�Zyl_��S �0=P�@�w�ݯ��(v
�ʕ=]#��V��2�%�n׆׆�����f��	��Ԣ����8u:ó��C�5���T��>�V��O�o{�r�0�:x�Q��j�{H�c~��9���\N�n��fv�v����ے(���5��ĉ/)����_$�B�	o��y�/(�Q��ȎðԐ�u�
�љ{M�r�k ���#�
�ۥ3��ьaf\v�l{zw���tz�m��ب圇�`>t���T���ޔ���[zw�Ҁ"��"����h�P�	�T�!�N%b�����Bm ���g�*v�9%���?FO� |�k���3�s�:�'�����C��JZ��� ��ED�P�)�V�C �9�2DǎHW�g�c &��7Q��Ʊ���8�_.�� ��
{���D+��6c�@�U���r�*1��w�>0����J���땤Ɗ[KPu��ȱk���������w���/`��	�wS�F))2ʹ�/��>&�o��_�2`W����*{|�������7!����&������+Ҫ�G�v�=�p^]��4n�EݴąZ0^�PC�D���u�"Ç�#kx�U(���x<��]^r�[�ݫBX>�'ҋJ}�����S�&��Pi��a���&�����˖�
���e�9[�*���l��4-�|�;���oBX)/IJ��H`����\<�[㗛<>�F�Q��Vʔ���'j(:��KO9������p�:ƣ�nWj'29��$�s�>�1.�.V�����#�:y�fz:|i�.O��y��K�u9ْ�?g��q%Z����ܭ��f�_����s���u4���[�� EZ(�||��n|����������Y�Gc��.(���xu'cuv�����\�+ki97�?[ދ�?��V71~*��pP�a ���,��{w�oS���iD��Kq�4Yj�A��.�{�`�p����rK:��CosfT&G?AQ��
�`-�;�<���x�A��x������b��X��P�
ς�N$#�0��}攠)P�_p����O��5�2|���G>�	=�E�M������j�UV9���}VV���39{�Rw��]%�������7$S������d��};5c�l4�xT�C��̂��\�ۡ��f�#+s�S3z7�N+������_\�M����wKb�M����=B��A��Sz�����������1�dd�riZ�6���A���'39��.�f�Ƨ���){����w�	0j�w�I���z7.��Y�ZXk̡�VяH�YT�e�Y�Me%��8Q%=?V���,'��c)�1C*�T>����(�����
؅%���!E����h�}|��|r��x�  &���WRi�$�9�ӥY`6���@�8�O�w+�RD��Z���P��b�� ��ߋc�P�������VĔ	}���LsΖڏ�-���;�
3����s-_�J�7���(�j�B	��0g��^�w7Vy(A`�F�����'8������'D�&�Kd}�F���QO�_�y�SzحTHs�9IE\�s�:u�2<��Y]:��4�w�hW�6�r��V�ɰ6�x(���lC^�b׫�R���ʞӑ\��Xu�*+�s$�t���2�&��Zm*�EGӆ�]��%G�s�J�nR+�`��o�����j��U�8�I�+l�J~��[��3L%��
��v�r��e�OHѥ���)�[����}3�I+��h�)5�m����8>\��k�ģ�B�L*r��C�$�1��(�}���|(%� �)w=nЩ���=hv�X�>�c�e֌o�e==�>( ���Y�D,����6+�h:��QˊOx�'�T�!�r�a���S��M�0SvT.KQ�~Z[ȳ�<��p��G��2��2�C�2���i�Scc>l�M�.Ө%^ ��̭�us�H.�뭼f
�����ò
�cXU_7j�r��q~LvB�ݗW�5[������.�.��O)��7*�MX�{��ROK���@KY �T��]�B��'�P�Mv 4�E(��$N��kd��5?ʊ�> �J��ܪ���KE�G����j��/W�o�����";��uw�8�`ڌCo	�5�sC/� �q����NR`�c�����X����A"���|�@��L�	Z������'�P��'Jk�ɏL7��rr���`���v��U�#�b;�X��Yn�����"���ܯ����fV6N��p�X�*|����Fz�eԘF8cN;K��]���j)�1o�X�r�m��9�C���0[?Ց<c;fk���� ȫ��|�[���t�)c%"�g�:_�Y{��Tu
c��Vz��7��8Tih��QB?��{��J���>32*��hH~���s9��͗%�7��'�aW:�hb}�8@��8�5 _t�I�����F��:�A�S��Yx�~X���a�(R٫@����2��-`�B�[�D*�u��L�T��i�\ޒ�ʵ4�]!�u0 SC���%�kk�`�'nc]hi~�}�(Ƃ��g��=|�b�< c��ɍy�@-`hZ�sd\�vt�S	!	E����"ק�@���6�5�{��.=�<<)��sآ�W~�#P�4޽���ĭ؂�S+S��3��7|��Tz?�wp&)D��R���� �^��3�r,�XS�9�"�=���<7�`:��t�|��'`�2���L�Gn��_2A�V��.��6��@Qb-�H�0c�,z��U�"�2в#g�O��+6��#���>a\��鸐f�ӶB���upu�/�� �c�*8:����T{���cF< �d�OAp:�A�\¥�A�E��YD�6���n����D~�X,ލ��b�~��8��^�G�� �b,����!��@SF��g�vj���A�]ն!SH���^'�F��Z29d3;_A��Z�tB
�����{@��$)[��Ö��X�գ��8�a����Mz�/i��^�N �	����Cndt	��7��I�\��+,��u���&B��A�Ȋ99{�Z	>�}*q/���VpG�Ƽ�6
]�H
�뱥-j��ӕf,LYc����3�)�C�kCC�E��(�Ĵ��z�?�@LZEL��RPlȅ���ٶ�~ҝ���Ug��%����5
ʙ4���ыUx���P�AK�A[BZ��b~x �L�K�k4��L󤻏�I�e�)�LZC����4s�>T��J	�(�R9ׂ�݁�����K=�)j�	UX��^�~���n���ڼmӜ8
��<��{�:��x8ӐC��%�^i�
��hs�"�o%��aT�׫
��B� ~$�ԸsG	whق��Ig�I"����Ab�R��#�	u���+G�s3��L�1]�YC��z!����:�;	v�k�-e�b��,�[��J0���;E������H} ����lX���K���G�a�&'�2��	]�2�``E���U���!;v�vh9F��!rYsH��t�/���]t�.�1N�D���j^t���:�HV���%�����b�Y��Fبl,����?e���ߢr��>�2�RL��R��р�
�dK�¨��Q�J����iY�|��
����	�}�fq���pi���a���mr����{,�m��E2o"��}�Fv���yȲp�[I��<�<�i����\�Ȣ��h�����uc/��9��骯Sy��:�T��mD3C��w��yw	^�4kk��ɣ��ٮfy]�hx�B�'��������l�Q����(r���w���
�)���/�:�6r*T���7>KBk��?Ϲb�dB���d�VKuj��x�N�ތ��x]���Y��qI&�}� -��(Z餔xy��]8�K��0�=nz��8+,����� c����p5Q1g�\��5(�綨vYӨQoT=q�<R�?oc��b�%b��bn9כ�q��4��<��L	"�����^�	8H-�v�̏F?�>�����ONo�3�}./o�C��zG2���z2u��!\��-��V�T��RQ_�x���τ@��k\�'�G�H\�B����	@:� ��Hؚ�^��)]��5��N��(���i0�;��wIֆ��F)� #���_�o_�����T7�	
z�;��Ƴ�u��Z����G�1�u�l����]�n]J�I.���Ͼ�ܛ8����\�̰V����ܭ�u�"��y�.(-	�NA�����\>+�[�O��K�x�Ѯ�����	.w;WE'ճA���]y]�씀�G��pF����@l���vʚ��L��&uk@}����j��7 E�� �2���qv�욯6��a���GXFӰ���c [(�tƤg}œ����E����xp .1�"����=_>W���C�:}�p��>4C/��v�����ȱM�!A>8i���$�c`�#-Q�DE��-���iGL0mY=���ӷ�a8��&M7��Z�rRm���n��ٗ�j�P-���immLn�_�#��n��Y���A3�+k�';���l��H��x�`�?U���;�)|sM�w_�4={ȉCfCqR^dx-����W�J��D�Zi4��c�\9l��"��r\=�����Xl��}�ֿ;� W�#*���5/�n��#en�,�QS�|�����˟�(�4z lP�ŢS�!�ɨ)�t9L��%������ pC'�<���9�@��Az�a=r�[7����p+Ё���	��GJ�5��T�RFe[vъ����g�!A�g\8/,��ܦ��_�sV�a]!���-�A����7�G��B��>���L8j�_����r(MiN�J��DG~�{ P������3��n!��hg�����Zt����J��v�� �g�{j-[�lL�S�[�	ɺt� \#Q�j�ﴚe�{��M�V����$����*�pwl�K�ۙa���u�d}+�E��/�'Zag����6�(]��z�%=����L���z;{����y����ϨZ��|�l��?]���{磾ǲQ}���.��u`N~������1���j>��S�{���o�E�ue��g��^���yP[ K{����E�L�m\���x(p�!vZ��I�*�}�?"F^ck��֚h�v�R��"�26����F8��$����T�x�6D�qD�
v���"�x��I�k�*̆n|����GQqo��	�/u*X�&�{�Ɯ]�Վ��@>��ˑ*]Np��2��6����R���V�j���B9�wh�;Y�j�W��2ᘫc��.�]ĥ����w��֫Ea�ZS�.(��X��S�l������,�exk��k�e!d!~�h	^�D#��z堩�N��c����Q.�3��e�2�{�g91�	�[#T��-���=�3M{XxvW��gw���K�Py;c]����#|�!b�"=�hs���碒���7��!�h	~�HNR耱�H����"�?��N��2���+�ߤ�Ru��$b�������gB�Ϊ��~�7ӆҢ�����P
�79?�=�̒���
��_�$ɑ���BΦ��=�� 	n��k�����/=y���o�Zy�)���"q��i�s�U��[�z�`��t�E������ܶW:ua�
�u���F�u��0�X�C�_h�����������1�]�����r���Ī�c�oҜ��"^r�>}�
��)��}��Z��8��u ��k�{ӥ�vT�̍wO�&��a�������L��?D<_�����[��ȷ�@��j��#L�IRt)%<���?�vu��E�w�ext@�9�~��ka"�X7�š��uQ
!!�'��Bm��D������c�2�$mT_������ �V���q*R�MWX���C��b��c�{'N�ܺ���4﹦� 	����$e�@-�S���'�/���֡enOn3��+�I�Uo�cO4pZ)�Do6ȣ��'��s��X*�� r����o��o�rs�;�f�$%!bn��aK+����������#q`_"ve>=�F��Փ���-K��/Ё�X�È�e�V���;�.lp���a�x@�H�̦i�ML���8*o���F�5)Mߢ��V$�!�Ŭ�Zt�$l������+�B�R�����ǈ=a�'��'�B8F�ty��F�L�p� }��#ӊ�H�M$��Jݣ(�WD)���ͮ�f�_�/�´�����@(K�Gc`�ʠ!~6L�M�tW�M��č��Qe�c�4)�h�(�RO�Ag����і�@��*fƝ;/�~"��)v��씷_��klJ��O�T�3a닇��KV:U}�e����(���@�(������I�=��$�K
)�I;*|�>���i{y��)V`.AuO�Z���P�ZWؕ����c�Ft%�1	5�|y?�V�}�7ñ�K�.�A� 3��Di2���S�^I�]�S�%F��m\Ry�@4���C2�Oz���a"�RY�HѸ�I�J�a��qh�}�k(���[G�.�:���5$��/��㑁�n�GҨ!)�����iE�0��[�u�B��V�(����Y�KT 1�N/X)'��4�p��Y?��{�Ȗ��4��Ƴ��7I_����N�-�"�����@�/��,����
!tg��Y>��f�{�ec+^XU���k�WlatMɗ��ˎ�^.s�z�� Ƿ���k�P;~o�s�ey�����f�})�ډ�{օhk�9ady��AV2��u#�a�13s�Lg-�Pؔ1�u����a�$`�N��d�� �3z"�%�{-�r�D��$��x�s����"�8�ϖ�nI���^�i���$����s���1"�2�;.�0=�0�����Y+\.���Q;/���YV�S��'��`g�a��'�[^c�Y�tK@+6K����	�I4$4�4����ɔ����Y"-��9Gx�T�ݕ���w�Y��� 	P)����!��	�exث$m����^���q��m� ��7�(VٛM�1�埻ũvΗ� Ln�G��\��֬��k1]�D��Sr�S�R�����}�F�"+N �ӿ��Ι<�/�Kح�  �N;$�nڨ�Q�߶���"�S�MF�e�]bY���v�f����z�R�:���yjuH���\U�=9g!}k��Ӱ���Ю��=��f'h����
j�fcj��r��a�;$��Ӱq�-Q�9�pH��GFD�z��Ϣ|8�g.�������Wm�&�.�ibY�,� a��b�]SJҴ(h�Ǉ�ܧ��a@�oGQ�{�G\D\�_v�J��,#�m˘�������}���	���:{�7�Xd��͚�!_�0�pK9�������ŧ`�,m�OA��%�����0*=t����#D� �I���?PzV�ཛྷ�u�8@��ᎇ������ҔCP�2=yB�g��d,�,�6�iM"UU�zI���t��h��Q�Dh�֎����q�ՠ������~,p�>A����zK����q�߹�,��y��_M.xr����� �z8���~7��k�Me�x�~���N�[/o]uD��Y ��F�u�:�b�Oo��(�G�R�m3��)�k��X���6ɍ.+��>Y��%\->}����u��K�h㠳��j�d�W�V2V���� �)[��F���.XeP�|�b<��e(�J�>{η�h�'�?yJ��h�:'�������HƪNS�S8<h쫇�}I����ؤ|�`c����[Q��R�$�"E�B���l1<��� f܃��|�my$�G��P�IH�X0�\�"���q�����8<�s4��m�7�\�F�����������?�q֟��5p�g�s�����5*J0�_���5��'�[�aզl�~/B-�v�����4��G�`"�B�d{�|�a�24$�<�����8�Y� \�g�/�јf���7���.x&0}�
!��_Vn�ͦ��ܽ�6���lM���ݙX�h�/��8+�38:�'�b�Z���<�"�f@=�Js�'A���i2(��?B����ea�?@�z))m��������OBG��) Dg��z���ss������?����\��s��(P�����*Ry:e�t��>��n�
�]�_�~Yi����3�Y�`����� ���L�S]��r^.S���M/v���W��̑����1p�)NI�&���<�4��l��X\�P����#�SԸ�3�a*҇�|�_�!�@��j�M%�P���}4rҺ3wHi�%��H� ����ֶ��&У���`���u6�h��=�}U*ҧ�v�+�I�T�Cs�q^	�d�YS�4��M�$�uM52P{� ���n!#��)x������tV�1ϫZ�H�yh�����Gtx;�����@��ag�0�Q��t��jE�/'�}���2@��oVo���LM�u�P�����O��M���������b�B�8M�r�;R�x�̋��C��%�#p�p��hz�#[��4�a:��!�N/ҫ��|d������r|!&���c���MNb`W<���%������P�^Y{��9%���p�H~��~ h܊wu��G�\#�4~�|`��:`�]D�+�FV��q�]0�m�S���l�oUP�D��5��&�ӯA�7�mŮ`\���e����Q��_f�^`�!�-�un7م�|��S4l$t�%�JYiѣ�N�1�NXbVЍ����qא��^bۆXcܜ�+Ag:��d�R|��:|�с�� #GZrD��.�p��+�qۅe.pf��+L,�\��o��f�P�t32t��G�;!->�� X���cF�@�nPE��ܮ�Rl����/e{�*�)kO����E3�vG.�e�N�~���!t2�m�$\���UǍHV��֫t(�Z��$� HDټ�b؈���b��iAG���C?�FU����@��	X�M-H_}�̑Ӈ���{ԜC|�e8j���*�,��$�ZJ*�Q��w3�~���^�s|��s}Շ_g���Ʀ��z���n��k��l�����'�.`� �A�X�ȸ�*H�5�)d��r�ۨ��s#��6ag}�fh��'^{'��D�N\@�d�����3�P��.�@��S���tV>3wy��i��F��A�i���W$�?\I������!�>�#�?3L�mدr#��(��M�d���K��^Ȯ�/ܵ��96���i�a�M����F���g��m���~��/D����%a��/3z��(l�`'�C͐,:O�M�@@�^'T�=]�F�IX���㈨r��%d�Z޷8��h�l?��Si��DQ�t'30وJ���g�%U#O����%���r��>a��rw�^~�Յ�
�Q���ȃ�\�go��LY;0c�fr<�W����.��K)�d��`��M�~J㛌�r�����b���z�'5�l>�ou)�B+"��`B�6
k�Uu�;�"mq�}�O(qUx�96�m�����d6�4��J<L3��6:�;i���6�qd��~C�	U�������]$��!�$+�,B=c���4~�Q�@�~�{ծ(/�bA*�3�!�2U�g1�Q6�F���F�~99Ɂe�����7G�m֧�KW�ń!��(���"���FѤ�ǽ�rK��|�0�׹��q/�v!�}W��%bK�2�&�=fW}zy�Ǥ�lc�Oi��pj
�7�#��:�9��8G|�s����s��E=�g���O�O%sY2�%k|B�e��X:���X��U��������Zd��ʺ���W�_9�����%�Eǜsn�/��5�@���Ώ����ߗ���vZ�l�X&A{��=-�W\�&㶵�B�t6Qt���xu���s��cn��za����t8vl���O�n�3����	���6p��w��Wa�:L�XX�
��΀�A&Wc�3��4ձ���/�=^�@ ^��#��ʚ���Td��W����5<�� \G�P���Ϫ��=]{����.�@m\��?j�:�`*A��R�{�PDeؾ��=�;��8�L*�'�L�����Et�<Ѕb�����	�
û&�I�Hy44���A)D��K(Π�J��|�1�| �]�	�YE'�K��*nÛ��rPW��s].	6�VP9����$ @v����x8��i�,���]y����WK�/�Ҟ�`g7����>&�)��zyE�؟�m,wA)�P+$w�[s���x�ܬ�2O:�a���h"|� '$���g�t���=X�N��B �(zTԞ�%�n���$ڞ9A�/��!4�Ѥ��J"g�YY|إm����:�ѥ����TY �{�q�O�9?��C��(��O�]�?�1��"����Bj� p�dn�n�� h�_qN��k1�Y� k�d�B��`b:S�E�G��lrJ��G�_������Ou�O�3v)b����9��:��e��4�Nf�Ef5�k�I����ZL�ny;�5@	kT� �~��(N-�����&�A�i�'��/�0練�)�D����)%N��ύ�̞uE�f��ڜ�^�>,nFbV�4��ݾ�x�Ԛ������r���F��;�/*K�G��&L6%c\�KZ\	k�ƾ���8��4t#З'�lS�"�Y�L�<{y�rP� ��l�a���f
�
�Z'5O%!����D�����������r�<�Λ�rR��<:���6t���Ih�M5Ϡ�4D�D:Q�,C; r��C�ݚd3�>����d[�X�D�-��Z�A�p ���8��� B!7c�h�JC�D��.sCL���Ama3��Z@r�`n��2�.�ϥ�y\��Jn�r��Ӧ�ym�e��7ӡT#�1 2M����ZMe�M���ג��4��<���P�N����Km�l���$��Z��/?��`�+yz�V��N���lK6"��</�{U��-qI�jX�Xd��,��}[|�o=�*�ϕĖ53b�ώ�鵤��p����/q)�c^�k��h�g�O8U��l$�� :QW伦cm�4\��'�9j�j�,���a1�M�X�@�X�̌�y�SZB���k{�m���#X�-o`���Ze�U���-�����p`=jGO�c��_����˗v�2���>�g�Qi16Z��%<�zX�7�/4�lq������*��D���0���$��~�]'~�S�6�H����OQ�>-���F��"F����榊��c���Z�	����8vo|�L�r}�K7�$�g[���?6~�G��s- ��8H;�khT-n�K�ƻZ��4���rE���{�M(���r�J�x��2���M��K��R�\Pm��� G�����w2?��D�ŕ�J.�9a������#tb� -k���9�8yʿ��"�|7���Y���)n�1�����fd5��wFZ5~�R3\1#��(���yA������C��W�焹 ���g�G��p�&E,�Ǻ��-&U��,>l�~�+�!���ݓ����Z��-n�N��8�O���t+��R�>"y<�E0*�����p�<D� �=p��_�����AK��hC'�3:�V����E�[�i������߻��@�z\Y����']me��ɥ!*���B�<�lj���{Ɉ\��*�0LTF&���I2,U�zd]}A˸c{�f�"�uZ��S俲t�,��_ovV�*ϴ`��S]������a���u�ڇ���g��CI$�.{�2�˒	"�%z���CB H�T�	3-�:��� ��˦�l!�a� I �?m x���'�b�^�V�]�཮a��t	಴5|MO�0�}�SÂbr���(�}E�b��������I��ߏ�ƲL�����3s5{s����R����;xn.�
6�j� ��j ��f��04qd���5��܂(ʤ���}`��r>�+M7��u��n�ܓ����&��C�u%� ���_�j�3"K}�����j
��߇6}��V�V9N��k"�U^ϞO�����[����sx��-�$�}M�D�7Ƀk��K�ҧ�y�����v���?o�pC��+'1"	�NC/����f�U�#�P[I�¨]'��ڏI�~�h�T5�r�U���Ϳq\&��&���逞�OW���{d9�5+�~�����Px�T;�eDlG'��r�#�%~\W��hZu�XA)�T�r�xZ�WuE����X's����m�Y�.>�bm��ҭԈ���{����,E���\␇r��ρ�1tгp��W&�ԝ��=S�v�}U^���a��:�[�Z�r��ƹ���Qm_u�G���1ߔ��u��R61)q9w�
�=bt"-!E�������Rdސ#-��m�
��;s���TD0j���ܝ�ˣ	 ��ԟ�X*^��T�K�[��@�vm�,���;�X>�A�I/�=��q��P�b��j�U�~�c.B~x��h�(
51��D�\��ەm�v����l�*v~}��Z�7�B�`ٓw�L�Tg2�cg%9�<�>x�6L���
�ZI;L�Z|vږ�Ɵ�q������-���(���J5 ��Ƙ���*
�s3|��~���U����P��ʠ�U�Q�z¬�ء���,�`�µ���{}�g�@�~<����0��c��^)nA�4�$#�:ꚙ��:�M;8_=)Y��-KM�Ѯߍ٘�-<R�O��h�*��]����0HEJWQ-~�~��Ǌ��ְ�R�����=V�l����܈�h�<b�nm�H�ie�o���+a٬@=���U�.��D8&�&lP�S}y�����w�2���h�<�r,��䳥7XV�z�ɷ�f+�6�F����3�ˮP�z�k}C�T�d����\}��}��DYN��1̴����R:�j/�V%���R�B�ߗt �_&*bef�(�ߟo���y7(9�j�󛛔V�k�}��+يqH��**~�_���~�~�*������>cZ����4�8��G�
k���gX�$��P��ќ2F���16Sޥ͞��ow�-,.�#z����S��A�c�\lWK�S�x��l�8�A&��g[r��[��`;2�I��=s����t!W9��\���"2�J�6�BC!�9�)��I�[>�<�-���@'Ӑ��L��K�ڈ#}[iC��J�����y҅����EȞ<$n4�m�8�yYsj/�ľ��1���_خ|��T}k�p��Ϫ!�̕i�1,�;���o�KiAu��NW*yz3F����;�FX���"�����X��@e�L��!�X��W8Yz��[�mW���{�Ŋ��X�+�N�身R�_'�-�'�[�K�k��ha��:[�xU"�j���c�}�ݝ?�s+YFPN��C��s�J���GC77���O���w�� J׾�V�9T�ay Ƀ��Y��9�
���~�-%6�=5r�E{C�.�Fq��	.��3��Z��!!z�29�-Ѳ'�Tݎ͊��̃��П�j��^�\�c���f7
E�\v��78��s�Xr2*��M�G�HO/sj	>N.>��B�C�E�	|�ʆ��S�V[���]��&�.4����ߣ&ѕeTm����4
j�鹍�!NW�G�v35��� �i_�yȿ�iܵ�:*>~�M��ť<4��r�ib���Y@�m�J����#6#��{+D���Q?��(O�I�7�:�O'�	�w�=c���c��<2���*[�Y��O"�]*�� &/�ݣK��*��%�b9�M�97� *�<AZ�t_���D�1���6�K{��,���d�&��ҺkT݁�,D�%���^�ޅ$��EH�=D�����0�1�H�����)��ձ�k��{��.�cL@e���P����G�٠�h��N�o���{��Ǿ�&����7�y"�������̅#����_��֕Ae��B��W���b�'��Ź�I�v���<��GW(��qT�zH��2(��+�=ם�3-o�}��$���W�O��7F=ǷC��i��::�K��?1{RE7�8�F�?5�>0�j���ؙq�
��FZ�ܲe����
��x7��[��W7�:�����B��60��\��B�%�S�<v����B��x�y�{�VGd��{�drcZ����Hזױ��*0&�:��f8Sł|���o�����K�$��=�u�{�YJKk��>�{I^�E�L�������O��؅N������}ZI����mr�ٞ"9g�'��3�����-��;�=�ˋ+]׆[�}�*�K"�L�K����e��m `i<�$+�"k�,���+���>fy�k��r���u�Md���'A
���[�=R
Тm���VH���b���ֈ����2��CV�����r�%��Hc�;MS^j'c���weۓ5�:��������K��FS����b�!@��*w8҉"���*I:�&��JX3����KҖ���š���pt�F������ �t��lR�^cd�,�v�c��Z�,�{������w@	+(�� }Pq^'�S54)7�����ݚ�K� ����S%��I���\^�|�lо53�w�c4sՏAk��7	G;��=>���q]��rm���.[-
����g�74�=8�A���)�~��3�s �Ir�Wϴ�=��rK4���MB�ӳ���Y��>�t�PԪ�MDJ�}�s��	'�VI�Z��[�=�D݈{;��cD�E&q���~�w��ڬc����Ok�Lm.r<r����=~�b](ڛʮ2�_\-gL�rQ�����PD����!{¦�E �m_Nr�ǕRIE�����8:�� ���j�a׻�v�w3��hY@�3����f��4@�D$�D�����۵�N�aoj4���$}������O�T}���ɔ��.�<�aͳ ��*Q���>B ka<�ډ�7K� ���[47��:d���!�v�#ћ���%�)���@�U:B���k~�T+M��E��t�+�o��L���J�ٺ��Bͼ0W���,�X�'a���(���8B�.�$�lrkv�ק0��4���3iIP�aF	.���{��n"ct4�s|@Z�o���k��+� ����EK�'��7��Q�!�G I����P���r�}������v.o��(�����r�e&�Uw�GmZ���x���@��=��-��̫��
P� iA� {ڱ�~\+�/�:$����@�B�A��[����,����r��zI��is/;��dv�ԏ����yz�u�����,Y���H(���Zo:���JW(<؜�+���Wz�vg����q����#�^}�L����F���jD0��]��4�XΙRkA��$)}z�v���t�8�i�����O)ԑhh���cZ��K���(>��aǭ� ǵ�{'W>��Eff�|0o�h��|RE�䖑�����hŸ��.[ˈh(�mQ,&�+�L�b,��v��P��!�H�0��YL��ȭt�=��J�TϬfܹ��N��`�x��}\Ԟ�դ��U�(�qaN�6�\�1�Y�*tAl�dj�����ҡ�>���å�68�ur��1.�ZR�[��Pb����p��~{sЁmm*.\�ɕ�TTz�d�L�=A����s7���s� M�"��wTyN���[6�M���R�m�7�;��TF��\$�0�3JVj��E-t��UI����a!Ե+�)��e��	ӯ�I�WAኃ�
j��eF����D�_z�ي�L����ɮ �8�����,��j�ݎ�L�߅��[c�4D�q0�w���U
fƍ�Bg_Q���>���nDK �k`�����s�d����Z��2O���q3�\�=�<��ْ��3S�� W�����`DoY����$C�n����@`B�xX��5��9N��I	��J0�u��'�_4��=��qs�~|6Le[K�Oɳǆ>�E�;!	R?��U��4�m���E�ܳץ�c�:����5�H��BXre9��G��p��w�����l[jE��Q��s���Pe�F�jUdM+�i�����Η6�w=8j�����㦢�?�D�k��jG]l.��}�l��DDhBK��}� ��rռ�[�0K؛Lek�IfI��0G7�k'1-#]|]�a2&�ݩ��E����S#�&c�����t�$� �j��º0�8s�$����[�J�;�>�kӆ�}�z�^ON��E�S���|]b97��I��
/2�[�Im�|��Aɩ%��,jw�B���vW4��~��#Y�db� �����A#�"�)%}��g��K��U}�����F�cAu�2B���eP~?�3&)�*����w#�Z�01����}�������{V_*(s�q�1;]��5���ٌ�m��۬�K��U%s���3g�Zbl������������C��t�%&�D��ig��D��t�%����>m�'a	Ղ�ysP���MT�;x�l�{�CJ3XB�P�������TI���w'SF$���iE^��g�+���!���q�@ɮ�Y�s%ȫ������9���g}�I3���u���+��it�-�3�ufh�g��P8tu⡇��zM�
���N�)UTf�/�I]!�����=��=�i���3Ɩ~�]�MZ�����q�;�<: S�2������
.X5�x =�Z�84w����b��uA+l�;��{ϑm��0���w���C>���Vk�s�e��0�砹��v���l�'nV�Z�(KY�LΦ^8����7�f�qؚQ�?7�#�v��V��A�v�uy�ԏ����Ч�lz�w����H��t#֢Z��!�8g����	��<�)�l�U�gY�m��.�FlW�83@qH���#�P�,I,:�G��%�oaMߧ`�:���(,v8��{s��u��.|�P���bfF;������{*�d�Z��:��R��8�����NG7�g����o�.ۦj����RQ��GE�p�%Y7�e���v'�:@#$�������)Z��ʎ�{Zc�uJ�/$�%��u
�Z�[�r�Q
dOx��HK{�M_�Ň�1�s�'7����Dǩ7���ش�\Z�3�,�u{�
�\�q ������� �kE�-��:��{S<v4�O����0���zs��ٽe� ��z0�� H�^(��o�?�6�q�G¥���-�$�2"�8+�Ȟ_㛘e�d�%�&k�G˹ȖVz2O�QA�b.���1!�j'�X�]�lk��}�P�/F��5p/+nM搔RHwp�f&�|$˟%�O��0����B�s(D���؈��V$��U�T;�y0��l	(U�n�XS�I�y�l�����t�^���L&v���),�o�,q9|K�]��V���ͤ輼(�<�k����B������m���/.VY�&��s�Q=R�߯�R�>"h'%3'\W-�.�1����f��)J�oY� z��I�c�V멏�nt]���Ը�
.�t��~���|wX�[���q2>� H�� ��|�n����SaDe|�im����t�N��1Ƴ����|KX���󹩶�v�����3*]���_L��{�.�O�Jh����ߔ����㈣�8Z���%����Gu���/�[T��>��,�Z�NO�k-���k\OF?�.�m�������q� %G|^>�k#�8��nD�r曊cQ��ݑ��kr����� ����[��2�"/?�� �b⼋�O����l^+��e��&�%���C1ե���f-F�ő�4���~]}��]�gIT{s�0A��^/�C��QV{P<�\��!��ʳ[|������]���N�$K��f�y|Y��'��((��w�	m�W�ոx����iVv�jQ���,�O��+�i��I��.@(:�=��w��]�-�X1��橉�r���!jJ2˴@�d��a�Y<�g��{��i��EEpU&���a.��߿��U�1o� Q�Y�$J/��)��n�!N3Y�n���7��׫�+jT�� k~��|���Qh*J{���0@�����p�w��ՖG$�K�xƕ��]���Iʀ�	�8rT�}y�R[����c�����M#�N	��+;!�NsQ�;6q����J'���{��Ak[�(�c�L���B`#��__����N"�C ynP^�p��f�s�_QВh������M``��v�P�Uz�L��U��(�O�i.�� ��'�U��Rz�7�?_<j8���}��4�[�y蓢Z�a �ϭt��l�L�f��R�(�9M*�%�g���8R�����WK�ӣ}��-*�����|����2ؿ��J�|�5Ϟ���bК��6G�b�V�ܓ�|KH���L���Lɋ��v���b��L���#M����/p�dU��V�@;8�s�;.l]���SS ��K�:�>����|;��M��i�b7� *�g�kgݿ:k�g�B�b%c(eIvq����OV�d���w@PT�kD�Y�0,
�/e�l12JI%��C��T�1�
<?󶆓����3��d���c؈)�bHKC���!�Qwf�{(�b
$�ņf[H��n����L�|�֟�d����֖d���y�.^�%�0�/F�s��O�ލ�dj&�E_�a�����(\����KhLь�8�޷��>"��H�̇��:r�޹�Ƞj�[!�yPp�1E��h��V�l