��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��s������\�Ἡl-�y�f�����f� �ѕ:�nA�kb-q��_���ѹ(4�dê*���7��N2�ɐ��+ٞ�4Y6Mx�ejǴ�y9�����=���D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�!��
��%Y l�׾�U�����w�7<@e
4D_��R�iؑQ��F�[�����G�8�h�Q�*�2�|�ejٱ�s�t�w\T_�����U���%yXAl��/�/#��Р���*�Z�d:���x�;��4��6���&u�_	d���Nj�Ւ�x��&�A#�+
q`�1[�[�$���W��r6��I���nH�Ы��O%�T�(�eܭ���L+�?��.��F�$.;�i01�p��Y۾����4jwu,���m��Iӿm|d�Y�0*�uWs�b�E���d(U0�1Gw�?w���&ӊ�2��W=�\v������q_~�s�� ��q�#K��R�S�k�WHً���+��#x��G?��f���
�^�^�߇�ś�j��}�<:�0`��K͡��#l������F
0u�7�:�3?K���4��">')�Q�G�Ec`�����շ�����L�y_ɰ� �T�,7x���_��F�r]�ΉE�9�����k6!��f{����m��	�v��|q�9�b0sz��/�P6�7�_g,�l%")}����2�������qs:�vv�mV)��X@=�&�ݨA���4x��X>�R��XO�!Dٯ1T�˦I �*r5�E"Ҙ��I�N�	%�j���V�Q=�D}^��׽i��߫�2 ���L�>����ܼ��\�v������\�xP?�h�,�Q���9c����1��,k����r`�ռei��:�4% Z)��sѠ q�F+y�\�.V��W�&�����%�7V/�*#X�%g�W���%���L��51 ٕA�fa=�n�y*�	xG"r���)b�q� �F��p�6���\7�����#A��S|W�J�E���5����	��� ��C��p@Yӭx��S8.���a�k�@ҝ9t�8��F�h���f��F�`�����������@80��.��*(�D��:�����I��oo��~_��V�����f3�5��ei��2�?P7@�j��ƞ��A��4L�on��)}��l/E��7�JJ����,tS���A��n��3�� �:��>ߖF�=�܎k;�wU�;������QS�却�Mu��0�;A�׮�.��s��u��ﯶ�TR[>��/�ͪ�ل
/�1�9��5 ��MU��V/�4QfT��8��0�pI5��
��������cR�;�Gcۂ�s]uۿ���2��;�;��ULo�z��OGp9T��>i�)�h:��.��<mP�2��5Zc�X��@�@��k���湵���g���lZg�^\�I7��F>�fT����@��w�ʋ|�4�?� Ȋۯ��[/>9*
�����s1�XzG��فV#���ܫ��W��F�8֐�1`�Q˘������@g��|J��)���C}v�y9�;��:�;�����~15�i0��;���`|����PA����~��X�~��j��$ʪ�u#�2��0�q
���b��=�O��b6��r��]7�y��×�dd��8�����U1µ�f/!��40f3���e�#b����_�a���� ��f]�e�@�M�z.��H=��s�y��	@[��Lg٠	@��C��/��a�{[nKC��ؠ�]��J���ܖ���V���e��|�������x��Ŷ��%�|:v\��A�u~;�	�#�̒�k�p�F|����l�V�lx���v���g�k�� �� �GM�p[�9Y�����i�@x�H��B:.H�$��Ɣ�VQ�<{M�\5^�j;�Q�����˪��k����|�f���d���Lb����I�:�J�¾J�4��m ̛�7Q6����N���k$�Ղ������r%�J������׊p������Q�T��i�~�[�si�0M�؜��+�'�a�2n�SM7t\ۭ3ޜ�C���y�K��ܕE�(�?����ö6��m�>�*�M����\�IGl���z�~�Dd�[k9�ql����R����*�:�Gl �dN<��g�/��./�J(i��	�To�ɯ��Fɦf�uj�ȉL�GxURZ�y6J�fy3��̓,����2�p$Y�<0y�|�0�~�V ��:L�X��k"0
�>��g�n�L��,�� R��,���!3����7o�F��n��}=��(^vH7r�sڇ�Qv�I8b����%
 �����vL��ur��o'�F-���t��^��X�[�i'8�*v4g�D%�6R�2��\b��*͜!-u��J��.?e������ }�`[ �etG���Ǯ��mĖ:�-�1K��U�jՁ��\�� ~�x�����咍�W�˔��<�D��p/tfk���#����s�.�(T��6��3	��D���v��Ň�*���ђ~�����Pnh=����cg��O��6�+�4�Rr1�_RJd�72�O �UNg���Yc�x����Χr��_��3��*vOt�n�'�����N_(��טݗ\�Hk�x~�	�[�D
������a�)���X;>J�$.�~^�eW'�r��d�zg�&Q�#���<y�rb�ֆ�IF�u#��5o�ck��������[yBKL���(�� �SC�va�NKv�r~��|ڜ�L�"�w�vҊ�����j�������oL�D�8'tb8NW�ka?vP�p�=L��Bލ͒(G`&F�@��x�fK�g-������۟�
i�GQ(6�$��l#��}���rFX���������Ιy:��֕8������}2�����3�U��&�P�������ԃ�s-@��HV�:ÅR[�̯�|��x	�Ӏ�f$N��=�ՊyZV�r���P.��;B�5��>@a`v988	w�����B�)�8v!��(Zf���k����@<��NYI%�o��F�uصKㅐ���ښ�+����gү��1y�z���,(8���ǚ��+���]�(����b��i8����Ý_g�{�nB����z��ǐz��-�"":I�t���q�أ5VV,b��T��R]�Py�F�_���U4O�Ȭ�5�X��퉦��"�$�V��t��\�xx���K(�f��58b�Us�����[;&�0�!~ �u�<[�P(���j,kL�dfԖ�V[%�)���N���։��Ts8B�4,���z�_a!rR?�;af��r�[h����մ�؃b�`j��\R٣W	��!"�a$ϒ/�B;������&����L�P�_ߏ6�*�h����}9Ψ��M�F���"���g�ԾT3�7�\����Y� ቜWL� �,z*	a
9���iʙύ����}k��ޫk�Gc��� ��+Y���~�4�m��ı�َ䌄��z�@:j�����_C˒qE�_����`��B�%� v���M�;'�2 S ��г%���e��=mk�_��9I�Ȇ٫�XB���50Q%\2����	������ƿ�h�ja�R���ܞ�M�f"�k�[g��}-)�/���H5�9GM7z�:�jˊ����\�5F�K��x�}ܰ/�~<`i���h8����linˑA��~C�/�"#Q��:���9�� =�X
7�,P�h�pL�F� i-�|�F�6��,e=f�����_xӵ3��l�͍iɸ�+��(�C"mS)Cn�Ej̟OC^L� 4�@^Y�18"��7r_�
���A��4I2�.�t�cea~�����hh�-&訐%X�K��.?�m Z���˥�V�z'/�#�g5>��ėb��i��Z���q_M���YQ����^�iQr������TM��;]wm���(�0.��ylǨ��a��8 ¯�G��B�"<2���� ��Ǯԏ�ᳩF����|&p[�m��A��	x�HN��[�mb�>�b��}�,~�Y�U'��� �ʯG���.�Gs$洪+m��L�X���u{�4��d� �{[ ��2X�'�C���`�]��}5���օ,ni�C����b>+�u	"a|����k���bZ�]��wk���	͟��"�ѧ�D�����,u�YV5�E[�m�K�3ԃĸ��H�d������mSt��� ��w�UE0� O�ʼg���)0aB���4�];T-ҷ�S�+��CS�1`�=[� ����z�8��r<{j��u��#�^(���k �Y�hm�����v��Uq{��M�݄g۝r���.��.�������3��� ����;��Ԛ��7ƪl�a�.���\��г�Z�l���0�Am���<*�eל��?Gh#G�ߒ	���n�X�G+�|�|�s ��$�85�ҥ���,�Ȣ�#<?mؓ��&p�ɟ���r��NE��8!A1����SٱQ��� S�M��j�r�xq,��~���V%0X��<����7�.j�;�E�������+SKU���=lGc\J ڰ�QhW�2Ƈ]��Fx�j=	?�ba �k���O��54�����;9?!Ro� ����]z��1DD��0���\����z��%�\�ɛl�>��'��F�Ս*�gܡ����u6�j���u�_�ǘ��u\$��	��M��=�F������|z�}܊p_~rpC,ph�����܂}c7�)ݟ&U��,z��NWG��%3a���\Ůˎ�?�/{=eĴ����a��<u��W	T½f1�U�0��{Dъ�8	}}��(`�G�d�*�G�"�|Ӓ��W8�j���?��8��ݎ�urf���D��P
�Ę�H�{��u�N~���W)W��]�o��
w�D��c�� G��ڌ[#I�@$����+�p-���e�"}(��d�N��\X5���-�� N�*7����OVޚ�RV�_T��)����W� ̂��r�Ώ&��\�W�:&#�g�nTyi��6:��w�>�"�߇<Q���@��͂�lxh���w$�9s]zR���*%�t!>���{f�&;��Y�F[�_ A�K*�$���J���V�ұ����,�����K`��u�*C$f�����&��^�hE�9W,6 DluU��q�9��9gkg��C�>y'<����4]$ͣ2dX#���g\��v�R��̳��h�[�ҡ��ȫ��~���9	n�떲K�md��N��è�Yӂ,$U�w/��F�$�\����m������:hE��=2�R�U���|�SA���m)D�K;��8(����ۓ$�a���#��4LN���%4ś�N�fIk���E8Fv����9'��E[e�Ε�A��:r���%q�o���z�n���g ~��M:^a�&x�Bx5��NۚĬ$7�ڥ~K���l6��K�+���}{�fFJsA��܌A���r�CG|��ī����Ё���2)�M��:���S��P��2f�S��)�&6�ig*��䔣�b�w� ��|�@{$^Y��bQǖ�^[�at��r�my�=�
���nIg�8�J,!3I���zm���Я�h�&O:�gP���h ;rG�P�D�-��T'�߄3Υ���G]�H�H��AL����`@�7���W�����\����R*qlX�,�<��Zf.V[�����y��v8���Iz�S�z�/,��ik�u��@/��a���^���v��\�X���*���+|�q2e<k���.�l|�Y��Q�2.r������|?�T�1�����/~��؋�&ؗ�vEI[H�3���$�_���D�6!�X�����1U?<�0]$.�}����&��r��4�ȗ���xU2a�T��>U9
�|�~b��ʋŽ>6�"d�{��0�ۜpqׇ��&8�<e���]�,�\�qE-��{U�W��UQk��L�Y�7�Rr��tid1�^�F��>���,k�2���Ed~�^C�������*��{���*��܍�u���I�/N�TM�S��J�.\*u�Uʈg����C��UUxڒ�V��p�B.��N�A7�L��g�����Ij�Q��4��T�#��6i��L39uaT�P�zQ	�Z���ji�I����0$��V8����\P��9x,�ȏ�T�?�Q,8��!6�� }B|�I� m�HbؒG�y��r�`B@�������%���~��Bu6D���✾~�`�@�� ��H2� �^~�oY���3'|� �N�oP��`�#�d���䰥5X(�^�Wξ٪�������kq�fs'I�ˉ�%Rr}^]�ELS���=;}�X������hk4@2�,��/So��R����-��=�a�t���q����H@S�0��,Y\VF/IcfyX�� �_�w6�he�S�o���
z�� s��l���U����J��2$�@����m��<�.*�c���O��ٵb+v�.Q��$ښc�x�z#^E5�R��\}%��MW����v�R��U:�P�s-E�d�����hS�=�%�T%A�PӤ�׵M�8���YA�J�Y�H���j��W^!D����\�����̝��6��Y��E��KJ;�YL6�_�-ݮo@ �?K^�zb8��;������S�\����o �7������7m�ÿ:��WG��OK���-�UB�RP��_�&�{=���y�=����pN�&
g]�Y�<��|�ڕA��A��(ok��h� �>�d���,�Gi:��7>C���P�6�K��+Ƥ:��E����(�zO�\�a4�B�'� |����X���d͏�j�ٖ�	�6��Y@�knHi���U���E��Bg� �b3ۏ��	쟌!�Bj���dVD�:f���6��C�/�K��"����r��q&��w=�~��2���p`�f��1���yw�1�64K�M
Jc�-p'���g>N/g�|wIcTKɁ�J('�!3I�`���t���'
i{>i}
���� `�OgJ]8
��{�� "���&%\�������tu������N�mV
{
��/��l����C����"h���%�8�����;�/��W hONm�׻��7���O��������L���������g]vQ'jW�I��)���L�VQ˾ʜ��V(C<��+����!Lџ|L�)�YC���}�Ŭ��Ps"!�J�U��e��̄p�0�D��Ma�M�9�
�5���q�a#R=�.�{*�^�CcG��Wi�J�8���&��)�9K�}�m\\d�W�%�������}��.�[��^����<
���idz��Yq�'���B�|��'��9L}6��Yx�t�/I�0�!t/�L��Q�-�q�������ڒ	7�`\�CR�Ξw��~@#d����s��^�6��Z��N'�g&�����K-3�������r��٪T#�	�����I�O��N,�B��4p�e-|#"��f�xR�i�O����W����m]�"���m�7�&�����y����G]�D�bl^]�0߃��	@@N�����2n��F`�Ԝ+�C��"��5�_���^Pøi���{+�VwLܞ6�Sjg�3�`*���~wN29��d0�)�%��t����	�X�*+\�����ngr�� ���$ҳ�l�jP��}��OPū�h` ,""���J>T�>K2�!4�=;������Wc��椫��sRsE>4�0.}����a콮�e��8��!,{���h��Ѷh`�����݉�/�6�r �F�u���~=�u�kP*qJ�6�ۼO����؛~��T���j��)�.���ܲ�rbDڛ�����T��jZ�=ȏ�٭@����&F�i�h�s�f#����׻��NHx/�+v�#)Wz�rJ��c��N�Ì�+>U�>(�d�� *�}]M��(���Yv�]�"�GD��#�M�3�� ������y�/eJs%�A�J3���B���J�>��<�x=���j H���&yՁ�ED2iG�����n4	W�B�%�&��m���]�Lf{݆�'�8�9S `Mi��h�&d�.�Gh�c
swZ�������h�� ���_$��ۖ0ӿg�m����:@�*�gv�~*�����P���Z�	B��4��M��*�i\=�#vd^Cs�p+�u�K�Մj#O�f��i�X��+�P8 l�74(淪]ޭ2�[�9��@�KNray����me}*���Q%����Ez�g�(<M�:c�}y؏�?LwKkE53B�y�M�u�P߈�}�����DT�9��aPPe&}�ow0�q6*R�'�
z%`V5\4|���
��L�o:x��/m��M;#�Q��?�d�;��9��^���r�p�'g�;@ص�>7�{m�N�R�9 �L���C_��|.�/���	�q��H9��E�WC
?v��;/������h$sZN��V�:s뫵\A��ܤLcU:<��Ǔ]�{k X�`Z-%�d��o"^�⥶�%�ׂ�m"{�o�qr�J�x���5�b_�J]BF���������$�|����ž��jV36n�GC�%��IŬ��X�*�V7�'tB2o(S�[�ݳ>`�l�X��o�a�)�y���D��2�q+��,N���p ��,I��{Qo��`ՆJ"qd=>4����7�����I���&DK^�86�X����j�w��0����I��Ӥ���SQ��K_G�&F׉7��9��tͅu ���5����'�JƱ��!*3x�$�_G�̓�,��|��,���2����4.u��0T�nko���}@�Gnd�᪘��rD<N�M�~KYwu%2��B���}le�����3����NZ��'uY�=�`&�?�A<��}���J�ʌ��2f��z���{�޷�)��n��oQ�80HU��_h����2[>�Gj��:���  @h�@��ʉ����<{[���)_���6CdJ�J�*�3��a�1��k�/�R�ժ�6�c�W���"�A��A�dl:�'�F�0^����Oy}��M�s����~9oJxۅ`�>3%�h/�8��WkA�ɤ��M��!S�v�P&���¨�z�)�S˹3��w��p�$(^��c�mL����d����U>P�>nׯ�����ޤ�V�����Y��^R�GLyzF�*Dˎ�L���]ن��_�L�}2�1Y42�8��S�;n����Zg:�thOk�%�|US"O�/�Vp�yx�v�G)4��H#�L�5#@7lo����V�KnO��;M]��V!�����2N-/�Sɠ���Ý��0�?/��r�3��y�p*�?���g���IPظ���zbL�	 ����U�"z�y�<��0��$�ܦ�f�&����C��_�����f޿��$���~�o�dN惟U�u� �+�I+����"V������{��S��>�;;��tRq�Z [�>b7��/0pd��Ab�Ր\�g�
�_.q���� $�g=���A�#�e�Os![mʷ���2�nyV��hsO�n2B$���v�P���`�'�z�P-���44��]���*��RcF��3�G ����%�=�\k�������~���<WTb� b
mnc���g!f�t$5�>oC���27�:���k��6���ʛ�/�VsA�Q��v��D ��%����uT���g���X4?�q$�ܺL=����<���ɝ��d �'��ozо���[f]��;t��8�?琁!Ѹ�v�2o8"���j�ߌ���_A>����<�AN��t�u�b�ڙQ�}���0�x�J�@�-=�-� �*YX�ȧ�F��:2����[��/eۙ�`���`�0x���,���n��[���w�zN�k�V�ˑ�s��[�x-Ri�XW�?ے�DK�������I����ʴ�qJ�\.�/��R�Jmj�!���H+ʀJÁ=GO1ct�o�}U���s�d!�����"�6�=�n��0��Ȝ�r�z�X�)���]L[;����tԵx~0�j%KR��CP��@�ҳ�X�Y��	%���%m���=K�\Q=�j�y�Z�$�sTc�N�$|��s��ڋP�f����l���(���x���	���j�68-�O��Sgo ��Ys��]��O����t`�3T� 	�\�&��A�f*iElW�d��/���Rv为��?L�m�A?�{K�0l\UJn=�#I�J߶��x��
�T9�RG*�s~�7K�&�
��^�M<�6�ɚXd2���M
G�ϐ~f���5�3�>���򩳸M:���~��Ϲ���U���g����x~����O_^^�7S*�����w��@�7L���#�Y�c�z���b	@��o���Y�g���ǫ���`Ʈ�c�*��z@�)���ع�5���M�^_&[�6�/��q!:ND6��rk���3*e�qfk�M�s��Un�7XW"��(�/q{�*B=q�Ca���6a�p�x�+��s{fw�t���G�7����A"��mz�	a�c6ԣ�C	!GCG�_>O��]�S����w�Ϗ�|r�ɫ<]���e^�Eg�P
�a�SxX���V�̙CB �6|�����R(��F�b����5���ۖ���z��]����6�x���8�����ϧ�:��+���ğPUcvb-�)|�cs��q��_����~1+�?ˑL���1��E��s�4�S��+���������+���*#:lՈ9/��t~�*}���԰Jk�Iڷk4#�DU�Dn$�G-R������T��qn-�$K�A~���a`�g�6�'��{�Ae�Ν��z!,��R���̾_���AWIe��l� 0�B�������[Tܦ���1l6(�Dk%{�_Ō�yc?�Z�����D�
h��7l�l�<9�8}�,�����DDh��!�/���`��2�"�;��e��D�<}t�~�a�}�Հ�և[�P���{�p��>R�ZLH������DY����5vdi�w��޴rh�+��Aĕ)o��O��[,-�4F�x�}�\立�Y�`�I�Ǔ4Z-�J��Fo�	�!��n1r��@"ç��j~d��yx�\�a�י?}'&��	��uj�ͅ��G.|֌���@(p�w]�i�f�ۚN���lo�u�������˒����v�'�\.�11�{���s<B+6ǥ	t�Gl�6(�V����X�ʴݬo��<
����?E�]r�Ͷ�92��t�b���~�;�|�6̉�٢xWae�R�&z�>�ݳ~��uƝ��N������k��}ȸCzK0d1�T��L�B�#6���y27C];��p�<��~e����#�Qh�
2��O&K�	(�a浕mJ��0�jR���Zng}�t� FI�|H�xF��<9кO7Q�W�+x���Z���w��xi��~����Vv7H�{��3���2ű�W�I+��Ϳt5'=Ͽ&���L�0`�����\�u��&�Ǖd���P�����d4�"��=B�O�OX|���4�S?�X�|i�0�~n��y��$�\��2��4ȉ��\v���i�y��xė4� gI�:���*�TC�L��Z�Gи�!�׀HC�MI~�$�}@~-�ߣ��f^u���,"1�3{���]0	�v��`',x��x�s�BФ��Bbq8{�-�k�0�]X�t�ܢl^=2/��]�l��*Z��I�������-�¬�i�1g��I�qN�|����r����e��8��&�e�JE����C%�Y~s6M�����qM�Vj�&t�h�瓱�X�'6�J#�^�#��ZI�M�D�J]�6HKׇ�[G��p�x{�$�ȝ)���-��P�������=�'���g��V�(	ɐ�s�}iMz3�j���C�.�J1����P�.�w�r��T
R��?�w�P���GP�Y�&n�>#�������U4�`�WbJbuogY�ƾ-�fȉ��{q��x�?Oi�d:�g��#{�cQ�8��1e���d�0�"\U��^ء��J@��I<2jX��K�q�a�oޱtE���}����*~����#�rd�Ƒ���T ������J�K�o9)99�B����X���Sb6�`	�
{�C-t��/lx���0��e���B8ثğ"���iYFs�|�a[���j�sՐb@����R��e������c�j��S¬|��Y!�����}'"�c|�S8�}���T�mI��`��;�	�v�L�(�';\·�a���X �.;�F�s�WK�M��9즸?1�P�ZW���|#��7 ��𓄖�-�o��;B���h)����(�s�Z!o��-o�f���~��}��"�	�.XE�όFF���Y֡���p�G�(&��N��X���]B~�\�*�E�����)g[����n���S��������>�6~��"[B�@A�)��5�V���vK��{@��ܹ4\ȹ��K�o:�w��xr>�v�"�q�:ٽ��Α�?u�x�DK�Y.������_���JpD�4ڈ�\y���5*z����4�:ۊq(��%ωm�+>�5�,!����X�sQ�ٹ!���s�ݜY�&��%]�８2�K����eO�����������n2��'�`c��l�%���am��cɱ~&������G��^��y6?�q���g�|0%c�7`�X�@$pGEm\8�x��pk]N�B�~�cߏ#��kvh����;�	����q^aY��K� ��/pH%���&5�Tl{MO�j�d`��d�֯�ݎE� ����qkC�X #�(G\&�t�����6T����_ H�MV����@�����#�
+W[�<�a$"!V�3'(�CtfdIy�H�K����K3�99Fr��q�͌�wiZ���0�?�hZWH�N�&7��m� ���َS'_*1�h' ��!?ٗ�9JC%��{{p���+/a{�X��_R<��$�����c�V��#�M�#	7۰�4�2��Y���2��=�y���n� ���;��TJ:>!�K��&����1Qv7.�}�����T��7��m��d2�y�����Z��y�XJg��Ԃzm���U��e�l��k���B�����z�A�y�.���S�H�%�S��M���iX�f�	<��R[�ϵ_M�j�e̨�q_)�.%�IR�,ݞ;]�d5��@�g$���^�(W]�`(+���������%�L��5V�!��
����נ:
�����g|�i\M������TK[��8�(rt?e1�	o�&�j�EO"zˍY�2˃N��^ݒ�M��"����<��3C�e~����K�V�R-*�e ��΄K�}���M}c����OΆ���־���{���=k�8��o"Y�i�����p�01o�ww$�H8��/�`��P\U���ԕ�cD���p��S�ղ�����ε2 ��ʞ疣r��P��6�����l]�$�>�66"?X�tԬ�j�˫���I�sN}�\B�?L�y�l���Hŭ��)��Ln��yX�^��CBp��p��&����|�t��Ü��[�u-���	x%]��H�X��)v�\��F�!�������'�Y����Zi\mB�J$@��x�Y�g��X�gi����/"�g  �x���{)�V@�j�b8m�u/�/����"(��f=lD�:
p��_����R,0q�1�t���.H�v���P6��vgH�0Ix4M$4�ʣ��_��N0?�b�(��z�<h��,*�������}yQ$b�����\46 ��hG��ȋ�Xit�ӗo���@ݚ\B����Б1�^�S�% Z(�h��jޔ}9K�O��,*c�^�6?�)� {�/��.o(�I`�1�ߣ���T�މ��B&_�����%[T3!-ϑ�%Nք���B;m���������A���=���r=5Tn��X���R��fG�g�V,�nɜm�q?R���_�+�h3�/�N�E�"8k�l���h�E�?`҃�J`Ͷ��*������G1�a�u�XQl�/��z\V���w��d��-�g��:.q���ky.5��Je,��xr�N��W��S��(�뇬��G���)�8�����< �4�[��E0��%���'�aF�᠓z̏S
�b?�!�7-*�J�)��޺�潏��(e؁~j�>�0�	��̆O:K���b@���JG���$���o�Z.(�C��&����$�G9�h8������X~5whE��<^��2���d�i�&2���� �X��F	���It��m��vh z�̴N��ow^�Yh֑�e��=�V��%W�}�W��ᇓ�;q?���Z4D0s����"���k��%�� �& �q�t�Wәv˻���-����tȤ��>����%��F
�)-T��zV���8����ј��1hB5�B����q�����Y�"ج��k+���椠�\�����Bl��aQ��TN��zT����f��xh��x`I�8\o�ܔf7���jV��]Z�w@J�œh�?���$�H��ՙk�(y�8�6͵���%9��4����j�"J���ʚ��b������qbP&�kq�����(��^ޫx�{�{Z�9�0sy;罉>�c.��FH.�k6)H�(��:�[��3Ji�h�vo~MI��"8%�&�njO�����dmŏy�?�,>�	N���b��AP�y���W�Sĭ���\�$�U{�f�R��$�&���P�p��`���J`E�	�F�sNl?-[�v'M�W25D��]�L��J���*�0c���M�2��aƎlĆ�K�ix��+�t���"�����T��o�Wĸ�437��W��m��������:�A�ϸ��A����``�)�305p�O�?L��lS��ǣ�%����7[�d��a��[=�F�T����?�Aq�u���� ���-��3�^�i�����-�s���o�p�;��=�8q���ؒ��������A�oZܭ4�"�iԊ�Z8Ź�o?JK��'����ư!+�c�
�2�j�/��DѺ�1�_q���,�Էv��`�0�	��O�ɭ
e����H_1�8��$M�8|�,�6����jc�>�em���%��7q��h��3��*,�(�K;���w���R��h�D8���x!��p!���?w($?���� Ӭ�ft�q¼����(�(�������te�V��E�
ysR����wj�j�Ӕ��G�����9��Y-}�p	�8-��YC;ΨŹ'��gyL��N�&l}�2��kǔe<!P&'��Vs;�#=|���bۦAqs��2�֢���@�.��OA�ц�|{Gе��x�~&���X�y�
2;c���.1��/Ҕ�"��±��Ȳ�_�����I�-�b�z��T�E{���u�I�a	�X΋�?���n�8ի��|�ē�v���"ac,<�n)�^���㓇J׹	�5�FAS��\�
�#��o�G��t`���:;4n���T,׷�q��'2?���#�?�̡z/�-���`E�"�/W<��c�ò��\J�:Ǳ%��Tn�ђ����Q�T�hu|�~>���ă����+�S.��,�����(=��f��@ѱ<��xu�C�d����e0?��S<�~��A��d>.���F��u]綯� �3pX�c��E��|?��w$d���ñ��n�Gs��"