��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�!��
��%Y l�׾����|R�bD�E���y"���فų��t����:�FL�H�>����F��HP�-M�^~�h�_�~I��I����aڨ(�U3�R@�%�X�ػ���
���A�|��<l;q2`�EJΌx�&&������S~W��Mtr�ʧkO��e,!z*7�GP�'�ߪF��Ep�3p�`��w+7�N��b�
R�ly|�\�A������|���,5��cR&Ў܉q�����	��L�ki):�=ӢZ�N?�����ul�ձE#���c��R|�H�-{#ֆ�$R���b��-���X��)��ɐ�tl�j����l�*�H�{ ��9�4�`�qC"�8/��-D����k�[�;�4�?i[��Y��Z{�㍸]���������ˠ|�,���vϺ�I�u�:w2�+p_�$'�1>Pm�hLlߠbǂT*��d4'Y�ᛚ�E3�m9��2�����h-��L`D��M�}r#�䆷<nmÉD�qّ�ݏ="8���>N�dN�FU�"^g�/�pЂ���H����r�B�!� Eg��JPC����DÛ�#�p�XWyZU0e�3�d��ޠ�aF��S�%�b��l�9~��V�*�9�΄k1YW�(����Mh������1��+��]vB�w�gv�|;��\�FRPB����f[�J�=��0�M	Ef�S���'��6�ol4���q�J�U�rG=u|sֵ�>��~�����?b�.^R�y%ˀL�u��,Z�qe��dpL���:`-�"�%�����J�@��'`Դ��\^$  8vt(MS�#^�����h���s���������F>����t�����=�<� +s�L��<�8��_�� ��~��3G��3�Mb"���_X���Ѹ�rY���H��MOq���<G��~C����'�0��m׺1�4�F�2�.�1���6M3�#�Q,]��pjd1��.�������K^oY�L��}�7�"��f�E�C�c��"ι�uO����@��Ԅ&ׯ��:���PTKS��Q3�j�6{��e�w3� xv$9;���&;=OA ��F�ad�*��	�k"v���@����'0ّ��R&Գ�-?�bs9=�T���%��l	�˚��v�W�{#aI���5O*�p�QD�p�a"#	�MR���֔.4<w��[��f'r�a�֥�*��h�E���`|ݐ�K�J�Uܮ�l���
dYE�>dq6���e��P�Y�S��0C1Ӥw��1��`@O}g�z���	����G/c�5Q[���B�\��_LT-�l��}TemO! D���2b�Gia��X��3�Մ|�m���/����i�Rrxh��`�A�RU/$�X^��amm}Js.O�%uV�Z�KJĶ��e��r�����	|u*F�#������*<�s��k2=�����b�N2e��s<�̞c�ƺ���K��+O�emR띦�${�)��[G�H�o�	��$�D�5p��=�"'Z�ּzz��ڟg���TB`|� K���~�s�l��?\��#��%g��?(oB8��./�PY��& HS�0���!��o�)z�	.�84����HN)YY�Dk�H���5�����GN�l��Ϫ�*@�1��6�8�uh��s{Sƅ��/[��`��0�L�\��2��q��5��W-Y_L5�uν�7'q��B�dE�K�h{L�30w�������X�/�������3�~.Gv��L�ER+3��v���T2�V� �M���4����@�o~٩:}l뼏��L46���F�V��:�l	|#G�,��5[;�@sv�Wc�^�+�de	��?8�21n�!�U�G
��//����te����5)IUW�b��fT���;���e~�P���U�z`8�}��KS<TrM�t��˛2Ц;�z����'yJD���\B�5�<^|�42���h�*x��ƾ-RnLfK�VAg>ǁ$�h�t���&�R�*��P��6��Y1+"V�����B��7�Иƹ��*W�$����b���UM[�58Q#(�P�2�"<P�vh�sg�'6L�������3({���@��*�:&�w���f�1�5	�1���VX��5�6�5s.�j����i&�����t�f��P����\�4fߺ���y�5 ��]x^�&���Bl� m�rb�Go�cC�ЋDI(��_ R���h�p�K�y>E��nx��ׂ�ab��6�#'��J��\�g��E���j��޸<����F�j���[���'v�6d�jV����9����%e�Өdl�5!��6���,k�v	�(~6u��lh�&�ޞP��]PR�ǻ��1k��2��9�e?z��p�����|�ۂ���A"KU�Vl(��.����F'�^V�1��5;yr5���� �N9�c#�����5���R��S���X�0h*9�������L�z�ۙʮ�Y�l(GP�^�Ⱒ$}58�]���ҊR"5�X�f�[�~�:6� (䧯�����2�(���v�Dd'�L$�~��6}VPd$����w�>�~��)ˈJG��v�ػ��I��V�箞y�
]�O �]7O��On���_Tx�s��:BA�&�'�g<�nގ�Gd?�; I$�pʄ5hcMĴ���nDc2�?�(#r�r���4��([L��8�**pL�#R�:�8ȸ��t��3�%��.��zt���<S=J�T���A���*u��|�&ꅩx�f��!�D-i�Ϗu��WJ�1��/�=��P���=��	�pj���?�Tϴ.$�(�uG��s#5�/OZ���h^�����'+'4YU8��)c)"#� S�gs�={9Z>i�D8[�U��/�����F�Hl�	�i������O`��y�G�
O�)p�U�U��#C�w��\�=�i���Dz��̪/�����;�	�{)�-��n�m�Fښ� �:�o��]a[׿4+>�E�译J]�@���hN�Ұ5>���s���K�G2T���br^���R��g��1���o�̢��f:�o�9��@�Қ�sg8��F�;���K5��X(���rM	�>Y�r۠��l�ȯ�ir�c��tf�09'Dc���ׅ?Y<��w�\N�������<n��٨	x��|�n@}@�L�a~ͣ����Q��%JS����ܒ�@�>-H���5���^)K7����F; ܝ�Y�uvJD��?䙚豼�Ό)^a��fw.�@T��@K��
�щȍ����pHr��2�8ɜޖH-���_Krř��Ρ��<�V������ KG�ѝ���p�Zs"S�!�\VʞC���Ss�8c�̳C��5,a�;u"�K����kIx�o���ԇ�Ĥ^����لv
��͙������,��i�����*�M�$��O�A�egFv5��������!t�h��C��&�������<jT-��5��9���$A�F,�+)�5k�5Zp�����������;�+��y�꣚���j"��V�ڝ��e!�8ڈ���!�Z��2�$�B�~�M�V�ǚԁ
;�T��A��5�Z��	�*�P�T���{%���Rc��g].PRJ-8�_&���A��3\���|-&l�):���VͿdU�e�����|�A~�3��Jb~\C;�1���8�o�1\M�`E�������̀�V[���*��\��`���,x ���X���+�������N'�CmX<�b�c�ut�Lp?�\dX��YF�^�f��w�,WP�x��^'���ڐ������U�O��vpͳɣJTQ��݆�x������d�×�SM��`��T��b ��p�E���^��X�g�gz�T�0ɏ��#q@T\W�B���;�!�p��
���.111�Γ��h(-���mj ;b�o��N�t�ݣ�I�([�rsֿ�rR!�6k`��V����7��a�ס�m�|x�zS�/������o�4�h�A�~�`���b�/Gv�W��ΕAƏ���J�a�ģy�4t�d'�n'���i�Z����e ��y�hOZ�z2WD��N|O��x+J�V��R~�ws�ڀI=n݌�ӜM����%R����`wO?Fz�f)c��x��Ѻ�� �>�w"��@��``C�Uׂ!��j�ɭy�~�Qʋׇ�_��Q���VC�ǩg�j��w��R����I�����㢄ndg!/�td��S�q�Q�G�R���G�E�ʼ<�á�;D��8��E>\S��v͸]$�}�1c$��O��C�x�m��$�i[7OIt�;z�Y���#��<�<�@+=*ev*y_sD�M�}"��V�2���_y dd��n�U�����,E��i~[�sw���:V������,���s7��1P|��`��<x��]��q" &u��3��5���Tv02 
���� �L����i�!�Ýh[P�����1ټ� u޷�H ������&��`�wAV[�tCB�4�&; ���=U"���R���$�wO��+�S�p"�":0Zʑ,�EL~�Q3���G��$�o�æq�P�p�C��,��d��B��z1��ۄ2)�h�l&���ߎ�.��7���e	��u���4�?mX��!�8�ٖ&�/�Ω�f4�,? &�X&O�?3X���sE**! ��<ǘa!�VL�7�`��;���gkU�@)��`�"�9�-A���F��������?��I]�s���wf_�d�R�u&UwA$���n��sX����f��A�ë�<i=�6�U4�nX���C���`�%vg��a�����!�[�]0C�a�L�0��A�'�۫=�L��z�ց���e8s��aP4&3��Xk��26����,.��x��tP��g*��]���G�3هG�d��=$ӼH��R�B �߯�v^\�(j#dj�!,�5gm�2�Z�S�k]����ȁ��<Ō��b�sm �o8�����NN�^��9p��-��!F�B�����t���ݖ#��4W=t��LgY�e��쉽k��~��������[���}&-�}��-�&$G���P<�?!^�	r���\t5�����m��n��<�L���:y�De?&U�j��'<v��@_��ǥ�0��-���b���&���sy((�9e"�.u�͑\j�����ܜN�Ɖ����b��d!�<k�w}�м��
`+���~Ϛ��H��S���Y5�l��FO46e4r%@�b9V�bY>8"�����F�;~�2f�����o��PQ����ˤY�L��� �|0��Y]�&@wa��y�f����)�+�W�j@�%��6c����Ho��˕��>J�u	a��~K]��°o�]��_*v�g
I�k�H%=Ve�G�����|��t	0���e�wr�K*V�1 ����٫{w$�Ti�jM��ߙ�+n��{�'��{����^�}�׫G~����T�gE�g׍��.jq'b7���b+^ Hj"5�`�L��`f�r�ӂ�	&bn^������2��6.�1�t#&��q����O�3�=�
����~Q ��q1��p$�Y�+z�>�� *��
	2ڐ�)\�}����WN^&%�n���W~��kRH337���{�.ԧ�d����;�A����}c�P?����R���������)���;�dq�3��������*G�<;��_�EĐ�6>�hT�H�3l&���z����]{�*+Nyi� f2js�ޕ��Ϗ^:�bm��OF�&z�Ů�M��ՠi����9N�kmf���Z��.ZMJ��_" <]��y���-\'����\�H���b�<EH�w$l��9y�U���I\~`��v�e^c�K1�mr ��P�s��0a>�2kA����\�F�r��c��[��ۦ�L�������/^?A�>kD�'G9��0��M���gi'�I���t�yF1|�����G�$ːe�{*	�.����ғX�86���(��_7Y�[��� <MBI �A�rX�;`�x]+��hq�\\[���9	�	�=�k6�TG](����/�.��+�@����3l�5����}�mԅR��QDԈh"�{�O�Z��[˪��eVT���
�$-� 5{C
(�+��#<�����Shw�<G~���Y���"cf-y}ޥ-��U?v���T�/=��͎7͜�P��:�3!� w����x���c��S��o��ڃ����8�w�+�}?�QQ���X�a:��:�Q�GQ����L���3��C�^!��6�uW~�R�����m����Kϧ�U�n.���!fC���W�\|F|���L������;[�3�5?����P1a�П��E�O��p��