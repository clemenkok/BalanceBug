��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�!��
��%Y l�׾���b����d�z~�4���55���h����Ƀ�ė���
��t�����x�d�:�KԈB��2���e��qcI��;(�[xkY҉zL?�v=�aj�I���y_�f`���A�$v�� �"�����o�K��@�r+��C��n�!�}x��x�__X�soR��j���dOz8w��:�3$k���R��#��QS�i�>P@��pJ�W)���wzX�"�4�g�k��e������E0A{����5o�҂����K����';��y�R����D�or�)1 Y r��.��Ț�2%��jp��x�cD�3xá���;� UoRdԤ¦��ݛ!/�>�K�
<������K�桴ڐ[�T@�g�R��+�UKq��b��j�lK�����f ��_��pe�����u�0�^���X��rk�6�z��b��K��ޙ!Y��2�R6Y�D�����yA�◘��Ϫ;⨲? w��}���0�v��eLv��a������F��È��I�@��X�6p��"��~�|��0�ǽu��f$:ҋ���~�K�'�������`�8z�%���=6��'>}|b!�!��P,n�p$�� l��e�O�A�7�Qx��}�^��YX�8��nHH���ǌ���_�F@g��D�����}�ր\��b�^s;s5p4@���%��;8�&�1��p]�RT���Q�{R�l$g���L���Ųk[&VK#�ﹶ18���|�NJ���k�g�X��!#�!s��=���:�+����bTlZʬk!���DI��p�:�O}0���F��֘��Ȱ,�$kd}��KE{�8����w�px*�������eB�4�)�f����D�,�R�M�膥,I?��84��E͊��ѳ�,
�l�ɉUlĠI>����:w��;��:��^t�<|z����jڲ6k���I<o��9��J"��8p{)yr��4mфX/T��F ���W�	�Sj���O�(��^I�_Lݯ��'�9͂�
@�̩e�����JZ�ӊrF)5I�숊R���0�32���Q��ߚ�<�Art���@���o9�Qc>��H�l�M:�"LUı/��	��N�[ͳ^2W�F�EDwR� p�D��f�Mꊎ�<��yj�>˃��b����3��`�]�_�ro��K��6��G1�f5V��X*'LM�C��	���맸��͒�0�܀~�AGJ