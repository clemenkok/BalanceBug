��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�!��
��%Y l�׾����|R�bD�E���y"�љg 	��djꎼ�Ϲ�2��w�8FV�z%V)��sz�7	�'��]Z���s����D��H D�}����\�5_ ?|����YD�7l��0sh��ڽ�c9A��(mZ������$���ٸ}�0��{+o��"9@�$�!���h,"e�a�F��	ekq=�J�>ii}|��������d�cu�[�������J���jQ���$r�Ň9������Ɠ>p>D�<?2nJ1����Qr�L�zl��q��?����$�օ�U������r��ذ�B������\��*��!-9��u���ދ�� tB���D�k��h]<A�c�ВE���������7���=�#��EY��I��s���e�K^�RVzbP�gl'v�]�¤����u����<˭a��qZ�/�Y���p�������WuDmg��)��}&Af� �T2�s�R�����F������>_�9\�Hn�x���)�K�LI�(if�
c�kJ�,�MɆ���v��#i�F�>���|d&���]��~4-�n<W��C��@����Ȭ�/f`(/F����6�EM`����jg�}�B�u����}b�,x���׆�<�7��F=�ᐗ?�9��`�~��7�h$b~{r��gR���� ����' Y�z )|�6��v,1�c~��H��< �(x0_Մ��(8�1I؇̘)���`�B�2V�c����f;���bߊ�_T�K�9m
n�ͪ)��Z�k�g��֣�E��$b��ۊӢy���.1��(�,��S	[���l��^�\u�J+%��u���"�f14hSnM=�q#C��FmG�����ڛ7�B�j��m�mv+�]<�ф����U�Ia�[�C��cȡ��̂��,�ѡ����/�<�]xWÐ0�e�&��k��e~]��Fl$%��@�q�����h�B]f�Ң���M2 ����h����X��;���k/���ֻ�Ls���ιD_{/�F2��z$�M|���ϒ��؁����9I�,q���i���8�-(Zj�����4S�R�0� �_�&�t�-���E��<}�l%J�I�6�N���v0�t��.�����hOJ+1v2au�Jԩ4L AW_*� ���.�(��%u�2$����}`�vRP���f;X�3���ٔ��f��~��r���K s�7R�0Y}2y9�Pë�X�J��}=X�uoeq���!O"����0����j�;y��h�[���b�*���#���(���UoCpHSg������5��"2�,K./��%��z1�T#[g���V_��d��Jy$e(�>�������%8twj�a2���2R��f�PNhw������՚���$�����)���r"�H����v�j�1��f�]��
/e��#�і�p6p[b�?zD%��|��J�\g��o��x�5�וU�r��0bQ��+~{��+&^)�9�@�	$q����u��x>78��.j4�.�$<�+�<�<?�HJ�vK�ʕ�q�jE�1��F��#Mٸ �nI��R{���V�4��\���%��<��3�o�����
|C�Ԩ�n>�wګ��	s�����.X��y�f��ۏ�n���K�c��U&+JZ��+��;������e����
A�L1j1�}ܧB�a��Q���.k�ta��_��iq_�r�R��&#5�[C�����o_i-�&53h�(9�.%=�S���B�\xt��+��;��J!��#� ��m��X�Ub�Z�B	�`պ���6�R$��xr��ʫ�E��G@�D�QF��^<S&�P�nޫ�|��p.�- tW��
�šy#/��M(N3x��Lb}ܺ����&�� �'��^���*j$
���C�˷�E�ITkk��cb����X{E՘P"^0�_��#���H�P%��Cx*��&LU����m���KATpa���]�O4C�x@]����Ȳ�����%<lR���c6g�bl�c���S�%��N��u���2�k���@-N[���(�x��5�2��N�%ח^կvj�@k (�$��&*�C؞
��;j�H�nϏ ؿ}�X�R��V�㢋O��79�e ���Iʟ����C��d��Ȫ�Do�c4�BB�QR9���r?:��Er���m4�)C�g�< ��H��|w���G������|#�Ҕ����G"����yI��o�Xy�GD�Ҵ	���+TME�Y�'k�3q��O�*#b\f)�q�޸!���]I��x>�Ԫ�ԙ\��.4��^@a�ȸz�E��R�T��!֞�f� �j�5��vz~_�DO>��Ƙ/�Ђ!;f�D��T��O��9��a��	�mG3�A�=��p\]tu������*2�C�aא�� 'c����CpD�b�Ϡy�G:�-e56n��@ sl�S����Uz���������1?)β)+���Od���q����(w��U�"M��}�F�/&xg ����3���_����"��Q���V1>���J�q�v��^���(��Y�<�rudu�'¿��}X�"�������u��U�dF|�[���2c�-�;MEꂊ��	����E�*�b�H7����(����/L`�a�(1�A-�ֲW�ɣ���!f���nN�����6j��Y�O�J����p��K���Sp�,NR���SL�����[k�^YA�^�i���6�g±��\�vj_I_@��57ۄ3`%�=��DZ0C`T� �:��T���ܶ�4c��~��{�7iR�����Ŝ�C�Z�X�*y�G-ԍ�b�ߴ;���p�WH.��֌�
�)��'�X�<�s�M����� =0!c6��$$��H�֟Wu~��C������pY���cm㾇�h�w��R{�̯[��,��S��Ǚ�L�\�ݷ�TA���h��!٣D1aT���|ٔ�3aW/t��r�X� ������$\�m�b�ܩ�A�X������l�����<��oKx�y�*Ǌ�o��o��/|0�I��9}>����Ӟ��v�Κ�v 0���05��}�XT��VY|�zP�+��ZiV�h��/RkX,RԎ��ɇ����r��\̏��|���ok�f�a�����v��{K��AvZE4$��x���~��r컛���Xn���Je�?��֛�_�1Q��5���RY��T�f)�ѳ��`���x��I��7��Dp�LV��0HZ+�2o)����J�ddD��B�