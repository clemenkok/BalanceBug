��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�!��
��%Y l�׾����|R�bD�E���y"�:�@L�����ӮݧBH�[
<�����ڃ��+y��e��`ݞ��G�����F,��Q!��|Y~E'�
�jM!�:�N^r��fzA�7��q���qn��#DK���4
	�9�M5��׾��O��*�$cv4H�(�$��=��n�D��)���o"����ӢE��-U@8�1D7��������(�j�BT�IRLVri<!�f�κ=V���Jё93��|��a�q �P۸�E��oJ��M���l�)W'�lB���t^��茓+ԦJ�Q�o�:p�e&���T�<��B5rP�^?NnCb�#��֡��H�*�;TVd������܌�f���MEn�$���aT�\�G�m���p�+w��C�er)+o��F�����P���|c��zi�kg�[�d�PՂ.&��G�>@����>�<��K�P���G«ɈĨս*t�t:�K�5s C�ud��D�1�噿t��R��=ijpq��i �x��~�Ƽ��-�#'�����|34�] [�"�� �{�_��9=%�c?�{��o��X�p�LD0v"Z()�|B�$q�)rO<%#)o�ݓ+�k�ם���l��`G��Y��sC��ɩ>c�[�yбC���0="R�-��RPI��� g�` (�<��n�ᆌ�^���|�,�b��ڌ��9Q&��mj�3A��ݬWEWQ���� e���{��!_ψ���U?�Y�}|� � #��N������=�դ�����9W�oX�=�}*�zqа�a�N�j���	!�fே��.���b��m=E�i8��� j��+��;^Ξ��/�va`x!���j��oi'2���\� �׀������W�x�;����F~�*�R9�?��L����_f���4��/��AVt�%*����9�u�R%:�9�0'���z��*�N䪿"8蠗#S�v����v�Ǉ���`��Y��\ߞ�!~.��>�5<֡G�c!��>�>CR�@G_胹����D�F7�9*u&^�ƣR[����{��d�JГM�FX�k$*	  Pˋ��2��؅��3Lb�x��p�/6�j�zb��|�9�TzA!RX�/�^��t283V��ܘ���ϝ� �����7���y�9w��� J
ТD9��smT��V�d}M�B*[ƾe���?�8gq�Z#� �G�Q:hz��ZeZ����������1��]�k�]�!��ؼ�b�q8ZƔ�jj��6���(l��>�x�O�0��9K4�;��=��`���P��/��>�mT{v����oXi4UJ�|����L*ܔ� Ȓ ]T%�E0D�HsT��q��/,��d�-�_Q,�ۤ5*hs��٧�$KU�b��"~fi_x"�W
���-u+�H�*�1�ez�Y��uД�$�� �!e��±����gPΡ$�~�&��l����u�,�p6o5�u�T�/��U:���%M���[�6[���%�Se'��O�rz)~o�?�:c��!�ϖ�Xv�EF�kWB[��#����@FK��
�wO� �n��=KsG �]K�����P��
����h�|z����yͤO��+��F���F�����htW�N�Cr�Zm�8��y��͆���/�j=l��z��$kܢ�����29�.PB���@�=�+A*/�Z�A�;�g��-��s��4O�$S�ͫ�	�ی~>����'�WM�ց�a���6�p�i�F�l���̭��Uf0��v�e��y�3�"k��F �& �l��o��>����?�Q좫�!�mK�(v�� �fP�t�SupGe��_Tb$���E��p�O/>��
z�T�Љ�N/����ꅯ0?���r����B����i�MH���챊y�6��S2F��ş �Ņ��#��7�N	�jwCޅ�c�$�N�^��nu֎��t�0B�ȃ��3׫3�	Ih��"G�<��8:W�[GjI�v��p�KuΒ�Qo�;|�w�>qJV�_jd��� �¼�/Ц�?��&�&Ĩ�H�'�<m���с�F.�9���t!L�#Jɔ���4|��O�f�p/�ދf�z�F?"�l�w ������u<�,�-�����/�{dYd�{�_^_Ym���J��xr�H:�DaA����<p�r!lLτtp.�O��.��܅��B�E�hc�(�`�uР�̝�ScaX'u{�]|�NQ.8�Am�]i��Zl*l;wl bs�L�Pĳ{��P��\蝜�}m��Z�Q�Z��%C<�9@�	o�=��d.�11���7$��k�f