��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�!��
��%Y l�׾����|R�bD�E���y"F�|��ݒ7�>�z�X����*�ֱ���K������eK6��k�H`�4�8N�,��7��l�E��-\(��Ib/[��wٗ�c�1.�	3�k�R|4�C!�W-B���Zħhh�1�gF��a�n6�4�D��ռ��-� �rs(�zI�*���:��5r4��Q�2��q�����X�8��u�Y�k`�ZA3.^ c�'�{�#��z\����)~?�g�����bN�����	$��S4ң��wZ/�����dD��=RI����+HZ���.#Yd�����SɈ���r�:�"U ��*D:!ٔ��B7z@���U�����k�4Ca�Yc>�H���)2�"zq]�8ª{Gg�rB�p'	>~,�Ue�^�����;K"�2�[� KμoE<ȤLB��u����K^�J~Q�6F1od�Cp^<���ۉ�Z\���C+���/y�x�|�P1>�� �6�����t3���ILP�Lu��2�!8�/)g��ь� M�L]J�d9ژ����-i8V����q��Q��� �u�xo���¼S�vKf������F�j c;�߰g�����45�3~$���Xi� o9�I(��D4��/�"�L写��u^8<�DKC�A-��(��u�?��!�C�C����K\o��C�c:��D�3Ԧ0��T��k3 ���}�Ee�W	�T��,d��}аL2{H��kU���L��mo��Aab�<+�c?��ص.�	���:���=�=Q��I]))�H�R�R:�>��D-�D����+n�@̇��+��0>�jpB�^������#��tpqIul_ݥ6����	�1�7�F�C���3�/[���R���&�Z�	hz�:������,����M��}�������m�׌˛u�p�c�uh^:4']1�F�4Hm�*��$��<̑��X��u�u��7&!��������-og��>-�<�e[ \����{}2h}y�D:�_�'�^E��y��ɘѻ�"����4.��]�i��4���
���Zi����#�� D](ieJ:��8]���@���c���?���X��Bl�:��G�ޖU�]ѱM����bS���Hqx�Gi��(5þMǅ`�b�+7v���O�y�3m_#Q�&Ug�kkh_ �e�L�Wγ�i�1�0j8�fh9�S��yI<��C!uf����������|��3$�����wc��r�^ſCFY��<���j�/���t2�b���O)>6Y������6��?��;�0W�O������zn���X2Et���U%"F����no��(�s��"���c��.�;��?|Q�y��7�A2�3�[4h�waB
�k��f�z!<��j`䅇֕�yޫ��퉘ߊ:�*xk��#�k�#U���q�u����{��i*�ղ�&�1 `��ZO�ȸ�h4 m�c�<� k�������DI�sWF�b��*��"�U�Ԙ� S���6=�15^���I�f[�~�k�-��[�Jnb�Ip8�7U>"Y�m�%��ğ��h�H"�Y�VJ��l�D��>7�}2�[I��苰N���G�I����]�j�GC���O�)��25;�b�b �x�kv�Y�8�j*�"�2m�?5fM/fwT�c��W��^�7$�q�b��N�i�\��簂�Ƒ�U��>卉�7�R 617�?YS���_�UC�2��M�_�4��[E1��7?*�L�Q��G�w��fڔ�0���{�R>��\xPM��}�7]ҐP��wX�[��bn�ks�*���bu���t��#,J�Y%���8�Q�s/�q��Z���P�-��dM��%�G�k=�N�k��W@$-'kV��2����F,5��>Kƾ�MO���=!Š��mf��}���`��3nu�|;�+t�;2�"����������x��U�zG,�"�C�;sÇ3�x�d\�z��$Z�����b�s �k펼��T��f,�?3=ī|Z*,�ݓ�=�c�d<�gzAF�:��7��dQg4Vh �~���s��ciPR�9��퐖��MJt�C����?w�\���T/�s��7���2'�7����� o��j$�Y���(�  4�x��
�uk��q�y'F�ޞ���u]�2�ߗ1ԍ��S��,���"�By�Lt�`�Z��s���5��_�]��2�Ls�
׺Јx6 �!$:H�W�-�]T�1�~l�&w�� �nc!��]Vc���@\�]��p�����;W����� j��R*ٞ��v����R��[�T�I��1�TP� �b�9Al���2��Lz�2���ж'd ��kv��u'5sP@	7s\����թ[k�Y"��C��GmMI��Kw9�D���Q�O�Y+Bs��k���᰽������3f!��0����^H
ˬ>�%-��l�\II��JoD$��M�-u0y���?됸!�z��k�W�����]��%��*[��K�vfN��������>�,i����Kp�/�h?�j��;rSz�#<L7�sFQ�I|3���3��t�W�vJ�20���^B�UZ�\[���F�Pk�Ϝ�"������;\1�}1Z2 bjN����u�� �v�Ș\
��v&�L�3����b�b�M�b+��Rfn	�ARR��hhN%O,�i�M��O�]T]�'e6��˱�Bf�?���\c�&g��YjqP�������[���D�8wm��e��\>mЫݰ��TL�1�/u8.�B,��[N�P����e�\{�yd�E�zp�+ϼ����}��M\?�n��Єr��s#���i5���ϳ=��!t������\�#���v�����y�#�#�=�%[� �V�q¯4/��^̾^{�"
S������?�9.�ɳ~�n�sQ|���g�T�2����φ��X��sSG_.�A�B��Rq�/�P��!��Aэe�m)��#"d��1���S�w_GKO�&���y�s�<N����߱,a�y�t��(�Ȧfl,�ZIn�V@�NxS=����Q&J 5c.�D2� d<j��X�S�ӼN_�gʙT,��m��KLb�A	��j�Q&��Q<�*34I//�#��)���{�:��@�XU:�����_%3~��2�ԟ�;�i��k�� R;�"�=.��:��.��z�
$)]��͑ʫ
r	5�܌fʚ�)�yи ��B打%F�P#�1�8���r�����J��^�0��q& ��R��Zkeӓ��7�`O�-D�.q����?�o`8kI�����ɺS��fF1<=	+f�P��<���	��3�K�Z���n�:Ѭ0�%l|���0���ql�I��1J]��?I��O��H�u�����W�>�û��J��i%c�|8҆V#�ɋ��3ۓ��2���]�J;0����g޳�SLf͚D }�.=\Uѳ��VP����j!aڰ|����q���ȼM�RG�% ,lll �+{P�1g}�! ���M�M���;_�$kOE� �M����vʎ�}x��%���׊3�ܫ7�C��X�6��b"6�����6o�սeuԓ��R+o$�Ӓ�j���d@�x�������c&y?�:9و9��)�5�J�������� Bp(��^�#����6��|x�^��rx� ��6rb�2;V��x�ˮ�Wқ#�D��')2���>����FD���*(�n�\=3XLW���ߕ��1kx��M�r��S��S=�'���q��|4�)�y�[3���%���?vu`���}��s��.b{Z��n{�V�bv�W�C� ��W_&s�;sٯ��B�r���T�D@��sp�(E�)Q���ul[8	S�U�7����?Qy�F�4�ɪnv6y�tZ����ٝ/�[��?���G҈��J�����Seݚ���Vq��Ig�q�v�~ĳ׵unMJ��̌���{D����K���q���l���$���v;]rIX���H:Zv�F�/�qIC�6�ݷ�O�?�a��OH�:=�N)!�����?x�Iy�VDw��4�?��^����YR{�}M�W,�y��{{�q���Aji���10fն�'j"RkO��r�©�Z�*nfǓŀ��.�Q�+_��'����~ ��s�"�U��,���z�a�]� _�e�<[������r��N�o;ú*\d��O�F���_�*:㿉�Z
Vu��ȕ8��0��v�r������Ao�s�]#��,�-{��=*��.���Z�y�c���-��Y��JE5ܚN�dj���7�v�S@&w�w²����i�_꽆5:����Z崃3�����+&,�b��XD�*��f��!"o�G��^���W�r�q�$N���o�:��X��I��Ե͢a��� �eq�P����@Ѫ��6�v��v��逬�8M3��J��i/�,�ZI˽J������)�ۚ^4�m��=��^��|�:!��Qڝ����������m V��h�g�C�yN��N�2�.@�)�B��_Q19HS�����yE�d]N��oǧL��3� 
�o�:��)SR��9s��h[��IC�vxV1��h��_��<��+Ќ�[@ʉ+��wǯ3.,%�U��\��6�I��1D�;o���y��;�>q�X�ˏ��-T�L�MY�?�'8���� �N����ȴA��F�Ӛ�P����;���5��X�(��G"|�������X��=y6�Ù���b��H�B���'���tb7��>�V�ǣ�-�Tk�TŨ}՟!�%z���&�s�S����5�i�\�M<E g��4���5���\J-�$����2�)�o�5�F���%���xWi�ƌ���g���w��l�@� >��{ݜI}�+� ��V��[yesY��ߑ�t|l�F��p+v|Ӽ�,�݀7!.���R��0�|<7��ވ��m���9cp����O���f�+�^GYCa�+8��� ���������>�l�b��T��q_iHe�}�@e���9{.N�ȥߪ�_�I�F��\���b��� �_U�dZl$��<_�|Ϡ�aRE銏��A����,�bA�Z!���������
��)�R���^�j��������z�I 5�ZG\�͞&��/�W�{X�S��ι\��AYI ���?�XK)�����>�t�e�K)@A�8��vg�M|���N�Ͽ��#nB��߈���:�>;���c�t6�e j�r�[D�����������\]�Y�ȷL�X�fn�AF�@y���k#��G~���ԃIq��#�P�rC�4,4FS�t�fz�*�����ć�3N@�#C��r8�[ �DO��ZOUg@�B�nR �G�s/V%Z<p&�Jβc*�76*{k���٬y�Zہ�K�6��}8k���Yl���c�P�}U�6���TT���T�j?q���aZ�г��0���ې�f� 9Ь����[]O��,�����s|
�n8a�
��Զ�TH����y��=��,910���A�y�$H�>��Hg����|�@�������@ä۬3®�@���D�NW���$=����'եS���8�����~��h�l~s���@��["LLh��1��
Y�٩ S����$D��&��Z�2j�b��b5�l'�I5 � ��%oL)ʯ���#���	��Pt�uAS�ʕJO�7�+"�����8@�2Z�/
�~�ޑn��<7�C�����~{ʹ�+��0;�g�J�$o8m(���wj[�=j���W�ky� �^&����c,I"�pT=+-#&�C��o��t�u5n�aT�^6�A^���{圭cT���|��XY��tL�^�H���El8_����ZM��,�0��E�x�L�X>�C�ϋ�SlYi��
Y�*�7�^p����Qݏ ?	����GU���Y�<_�\Y��[?�����`Ac�CP����&	��|5�>�z���8{YR��&�^����9<[��!�j�0��������b+;;�+���ѫ��N�,������������/*Y/�Z߄�otOu����`�)��頡�³#2�o@�^#" L��r�{J�2	�@��l�oƱ�O\0�wo%��R��u��x�X��`��<y[\���.
����p���!��|V��U\�gL�B��1��iZşAF"���:�=�J��)9x�%e76Կ�\�MOJ|˺+HH�F&����<Y�|㿏�X�#��×� W�2%��:&h�d�?����{Wj���Q����2��%�(�ݗu�D)�<2�1��V,�
#DjX�>r���x���<����<�<�9@�мz|��TVtEZҙ�M <{��b�����.�`6�.��!G��*I�wcV�H$0��o"�#����Rц�|j�|/E�v
d�[�e�TV}��w���̜(y�\�艅s6�K�I���������}
$�&�b�P�e7Wp��9;��!.��ǔm���T�cU��?�X��~�@��eN�����&�H��>��Դ��:��K���m%3�9�P��l�� ���8KB�*��R��I-)GC�A��GY�Tn5e4��B������N N�r��;��}e2(���q:=��u���=B�n嫕��*�ٙT�@�<؋��7_�4��S£˾��K�c�R�ݟ�z&W�l��"�cGb[,t^�V	�#:k%�x��_���b�4Z3��2��]����E!~��8wi^�%>���!�G���<j��$�9��to�\�����lb��#�����Ǣz���� 杢p���K��I�۱P����)����b�O����Y63s��8U�Q���o���Po�+�����e��ݐ3���	sd���	qP�(x%F �-"�%hmU���N�|+�2[f�E���9��q�����F|����hԮA@W	��5{�R��Ʃ�.�x4��W����*H�'�f<|�L�P���{_��ի�I���G�h�4۸�~�~��Pњ1�נG�� ��di��"��(��aD.ƍ��[�f�����i�sW�g�<�D�C.0�Z��P^	n����'Ao/�Fˀ{�&i�)�݂hϬ6_BY�;}��~aL��ueQ�DgsoR,�01��)/a-�#�����H5B��ܳ�7\D�'�����1�K�&,�dQ�+8E�Q#�^���֚��q������_�ѫ.4?�B�ϴ_�c�~N�)>�e"�Է?Um���$'ުR���0j�J���$'V�hպ@���w�if�mf��*A�4�ܦ�z �1�A��K��L������J�t�o��y�/�xk��JL+@�I+
(je��޺���WdW'c�7ǔ�_G)���]:>0/u$��af�4���Ϙ�G|4K9^}+it�= ��2q�΂�����o:�땅̊�.A������גƺ���ro��N�Py��e�`��cNF�ad -�:���@���mq3t���j�k`��@�
�Pj�W"J?[@�(h@MU-K�Q�c����\$�j��$�k.��/�DY1���7��\� u�U�7�ͦ�Rb�%*�Hg"�.��T��j�����k����p���i+8X��l�l�}բѻ��(k�%��y��[u�>Pݟ��2�h���)B�tD'A��g�Hb5�����p�%8i�o���}��PN2`4�do���3���0����N���"u������dڀ��VͰP	�tK���@��|��c�!/ؐ����f��}�&3������i%�e�<r��������wg�g"W����KW�e�Q����_L�x��%��-@2�!�A�ѭW��1���̏�,�-�@�Bp�TPϤdvk���HF���J�:0�1�\���Tt��I�<2e�bC��Es���O��w�?�\�s3�T�K)�
��������-c��bY��)"ԋ���)V�d��t?{�O4���Ң�j�� 0 |$��$�mr/̱/��X�{��
вޙ�=;v�ҏ�TNǩ'0#d��A�<5�/��YOZrыg@6��w�l�)]��vM��9/��P���ЈV�Z�*ˇh���ܷ����2Nqa����w�0Ne@��W�-���b�u�T��A nnv�uvЬ�N�Y
Гay��UQ3�ߒF�*����:�{�P��Ѝ(�^���3���6PLP�:sN%j���l���D�N�]���?�L�)ل>xtx�������m��Y�"Ծ���Oʔ�s����%�Fc�ū�F`�\l$/mZ��U>�x]����ծ���/oY�u�l��L�-�@��a$3o�߸��)�5�Y�(ОHu(]�����6tE��y4��e�o��L���P���lk�W�6�)�`�:A�e�+��>R�P���Aށmc2��Z�^�����,�<�Is�̦H�>\�J?)�Dc��$�48b�z�'mS�ֱ�C��<�Du��ܗ��l%�H�K0V�UD��/��H���L�N���g���L��h0ً(����!�F�(���W�z��<v��:z,�a��s=���6���2s_^�o��~�˹q�� 
n_��%���Ba�Cd�I�7fu�B��2��~$�s��Y/ O;8�O�L�y��蚢 %���o�Һ�<]:|"��Hh�d�-	_�r�]�@������R`�Yi��������e�c��t}᫟g��TW������R��Y�p����u0)��;GB��0s+}�9r�]jmȨ��84d~-�Z;a���{Ϛ�UDM�X1pT�ER��#t�Ejb'�?z\#~�G/�4��-;�eg��Q�p�U~b���� a�m8c��r�z�3,�_�Ja0�X�i"�n�2J�+Rf#��'?uy6�ԡ�r�QV�qQo,�YdS��{>z�����n�ā&��~	6o��uv���-n�`��"r���:e��t՝�0	�_c?���>�b�>,��C�(MwZXV&��v�����_\���YH�x���(�)5Lj����r�4��,F�c�J^��]��t_��g18�Lt,z�<''�6�-�`�A�x���n&'�X�C��N��>��vN,��U�,:y͜h�cs�Y3������-5�1r�2��%TZǠ�D�XI��]�P�ݥ}j8��[.�v!yf|UEg*JO`���?��Z:R��I��^Ӈ`�iP�틤\�_���<�UEq}g���O��]lÕ�$������2��.�����<{�;��W�)�>�6��K���F�8	Q�8R��\��������%< ,Wi�%��W��F.�K��'��9zZ	�?�.�fk��� �s�Q� >�!<F����hq���.�̝�3�����~P���^����2)	*�4[�ڀ[��:8�6	���{`��)km@EI[S�ɴ��x#F?C:��K�Ћ�ӂ���BF -�|oK�fd���s2��p6�����%{���YzB�+m�E�iB ��%�ѨsC1��ʊ"�*��V��9��dq(���4�t, ْ�RE	<�����$�P����"WK~��?�q= �)t�^%��\�3���#@�_Y�o����5�1���� ��<r!�u w��KE]JQX����*ե5�]�J��!Z'{���1z1�Է@�j�4B�_�B��q=��.^ۖZ��=�c@4��
�xg�sugw����F�u��_�(��(\v|�4��W�C����zj��5a�%�5��n�g�|�8��^]+D�"VOz��q��U�=�����I����~Jt顭���� \'Cʹ���}t����B"6/'�a�j����}tw){��9�i����@�B}�a�2�a){� QT��M6�����}%�Q�1\ί�`Ѧ����V�c�\�R����BQ]� ������~�I���ߤr���2����|�l_��6�l�aǆ}t�Gd��2���ȴQ��z�)ʮV��;����r7���B�m��*����W��_�8(� ��5�����Q�;�L�������F���2]ũ�uy������ȫ?��H�| 9v_��J�Cp؛h�j|��J�UŔ��)�����<��fm�[�ҡ�r��z�>,fຢH�Ao�\Qu�S���P�3͞��/���\e$��ٌ����	�T���bp��F(�?��5�?v����_NC^�;O�obX?����hq�>~�ΊL��
}��L��(���S-�����}�=L����4)�	聇e��bsO�����ll\�~��2�~C���UoJ����D� 2�"+t�zT�������h�"`���I��",�,��7��TB+q	����t��/1م�d�~v�)�� 4�R�]�,"��Yd�72&�"P}�`���^��$�m~Yԫ!S�[n"��w
��zv5��Dp��k��ز� ��6��R=ʋ9�8�N�U
��*��S� ��KxX�e����N����'�|�`Ԇ�����Sc���Ju$�Vɛ_�s4E�&uE5|�[�v~��98��,��qg|�Rp��kO~����(=��U��
 ��mx=a�߮�#�sZʳɰ25�l�Ad�?�K9����Kj�N*Q�X޿I�*�CWX6M3�Ǝ�"X����v��!�~"�ʓ;�l@�c/�ac�N�*����uhX�Q�:��T�H^�N�v������9�F����u�-������W�M�^{��N��|�x>��d-��[�wP�����?�,�]���b�ⷂ�9���.�0��17& ̰�5�Ά���(t�G ���b%��H������8�����[8/J���:
�GMF�l�ƊЧ�40�5UE&��B)����Վ�=A,]��G�U8�����G6߽�+b!����o���:�b��%�=G2{L�o����s,흔*���`��=�c���񮨘Q������4n���}����%���\���h���[����_�����]$�(�L����?�4�\~:9o`iJK�Z�Ti��B��WS�c�7�����E��n����:/�/,���~�:��S�S�%awH�JP��d��
]�P������o^ǔ�P���D�8�2��!0�\\��g���[{�yG��2��O�I�y�sC��ZR�2��f���cSkN�&�n����xi(�h�=��Z|�5`|ONcx�����/x�A�P�0u��L��)%�ۥ�{�N�i�JZ�W4S�.�b�T���?{��ƺ�ۣn� ^Uw�F� ��/|��}��ئy�Q�o����m��XO�����~�� �
���>ǥ\�����|��il-Da�+�Z���)�xx�Y2���!�W�|Yb:o�k=G���-Be��{�'��?���O�`c��^�ޭ��D��S%\��m�Q�m��5����3�aӄo´�:*c�yv ���iQ�������N�'�fP~����N?;(�PU�l����.�Yn!�E�1j��R���Se+�%(��]_�c��ehڪ?圗	�*��G��ҁ�*�����e�̐
�Y�i�qz�F= .�hV��I��Iبs��ߢ��1}�EC}��)���~DWM���)����|��@�AM���p�����Ħ�=���[Pb9@���X=���W�TG;c���c#{3Z�Ã��,4��4jq<��ϋ<��>gϥ �0��ݛ�Xl��l�� �-XvA+{��W�(=m����l],��\j���e�q-�7���l��R�D<����^�_���`�ۑW�{Kmү������NEG�]V�th`-yY}��(!�0^W6��RV� ���2��6V"!V���������σ�;�JF~D'c~���2�{^��OS����s�#l�N �?�儍�
;]P����C�jM���e�T'8��%TQX@�_���#�9{
˔Y�H���3�C�p��a#+f<T���@��?U�C!О�7K-�Y�Rh���eR�4S�wO�Y,v�?���Tq�Jg
��6�h!�����������lX�~	����W����5��������RX�<�Fv֛��ꢳϞn�((B�&�>�Ѽ�����l@ȅ魒�����T.�]k|��{�k�B��x_/-�]n\�L��\��wS�,r�"|��N����1kk4���@���yp51;��wy�
+~�Tl����H2�Zcj�/���6�vN��
�J��g�b ���"ZoĆ�Զ�態��Һ�l�~��l7!�@x��9�ɭK&��{�w> @c����A!����E7rO>���ȉ�����᫘"=�}�7uǚ���;�G��?\%3|�s�FyD��/b�`n|�W����tx�1K�	�ĺ�aTnO0� �x�4Q�鑇O�1Ӥ�'��b6C��T����
�S=�
>m�٪���: �(����`h,�m�m;�XN�k�a6W�o�g�H-�/��wK�2�h�B�B�~5��,��Kdȷ��J�}��e�T�f��D!i%-�ը8ۯ8�n�O8���4��&���&�b�HsЌ4F�>P���g�"���H]1�&���-�/�(��~:�d��K}��]����3�y=`e���S�j�����!X�P)�@|��<P�h1x��?��FN�גq���k��L�hZ�s��K��Qr�$�اr�pk
��s��3�~�`���=�y
у��E��,�����#�]����R!�e6�ɗS3NټA�5A�q���	�Ow7�**��^�,�x1���s���P�ȱh�3�����i�Zq��C͢���f}��L�������UUjg=}�k����(g�"�+�c���������|��sވ ~��u�1ɂ���E\�B]K��������Jz�ž�r���_��w��J��C����\4
;�9�䁎\�{sV1%*8\^{]�A�o�^A����J�-��v'`6�4��ߪL~���#+�]E���Q��/de)�4o�����,���ô]X˅F�s7k�k�xZ��b�vA���碱��r IB��݆�!�:]l�Է��S����T��=&�r�<�,�PՕ-��?�R�NW�s�2�g!-�U�w�M��T���j��G��ZpWV�>�ل�A�t���3�0�1|��/`>�WLf�E!%�����LX���ƫ���`��yE�u�\`�����]��4��m��z��g '���=�Q��Q?����1���P}:�a�ϻz�Wp�!Q���T"y'��D�|m3*�8ׁ]wuݥ�U�̆�7s�k]u/���
o�S�_��6�aY�#R��ᨴ[8��y0��W�XVPZ�40�
Hu#.�O�OҴUO|qu �&�0.�4[>}�Z�����9��T�ˏV������2��]�?/�D��Y�D�ͮ��"�z���l�1��h�qPJ��_%F����]�`$��C���H��]G�U�Ű���Gy��Cm
&���_(]��!�լ�	�ug�!�~��fm�h�Ԑ�Tی6�@e�;L��2Zi'�<4�7I�4�}ҿ��=��R��U�Ɗ���"�/Hx?�B��A'�R�NТFs\�H�@!Ϗ�G�<"���R�Ǡ�0#���s��ސd��씒Ο�ؕ�T ��h	Ȅ���u0�n�	�Q�<�D�OhVGY&��m7]]�b!��:���è9�
���䑕
���;D�d��*�;�?��[9%XU��W0r��b��W���Xc8 ��|2*
8���@h W�3��?"�4��X@�p���NѰ΍�K֟�(C�P�GR�ua������#:Ǩ�u@��PIOǷ觅��
�x�z0"�b�L��rkw_��&pB��'���DnUAuP�B�W�6�z���{�6�i]��üj�`�}~�@ҭ�CJZ -��9�6Ɣ�yQZ�ی����aR����\��]0~�J����$i3�)R�6�<s�;�ˈ�"�$��y�vρ}�&z]f;,%����퐫�[�Cok{�����?=�S]��f�:�����G�����$��M����h�j��^�#�V8��~��I8uu+�������la�?�E0K��P��!;Z�����Pa46�D�@S�Ġ���F҂fi"�$\�5 �ͩNjǖ�-o�������`}Łe�q����T��O�(|��}#Pa��?���+��%�|�ƽI'!���Yw);G����*�w���E&��W$�44(\��F�Z�u��������Q�K��(jx�G�<?j&&O�&g��.��H0AUg�{� 9�w�E�_�y��k1a>�I����n[?İ�#_�q�j1GnY]y)m���c���90#5�b?oW������{�j�������RK�Dߤ G��In�I���!h�Ž<cKC�"-��YA1 ��s)v�veƵ��z���M&�b�Inکac��(�m7�>� �E.�N1�s^sy�=aK�%Buf��2}"?	�S���=��{�d i��f�(�g�Wu����/���gih�誤��ly�y~;Π��E}��l�
0��:n�#�[u�v=,k�BFހ�wAܔ;\=�������$��{J]
����O�_��[S)S��j�
�H����X��Øq1'ScìQ�HO�}P�Ñ	�* <��ZP�+Л9��������&��e�n����`P�7,S�@J�!&��20e����=%V�Ks��g/J�:�Mf^Wuj�}�ʶx��ވ���R?�|��j";A䄡y��ٝ	�O�̚�W:��i*���lh���"�\���r��Eu�_�"���E��u�\��>���h%��݅�6@<|'�z�u�
q~w�V�U4�_��5I��?�iG���)��0ˆ|d���{X;��&;��ń��X�9,��S��f[o�a�z�s5{2=y�>���;�6�w�SSz�Ĕ�O~j��ƐK[����!"H �b)�9�5�g�5���^K\�}��܈)�B��xaT**-�5J����Xxmz>�s�%ɐ?}�g�,�/��kt%�;T48��:�7HU�2��j�<��Elf��U'�����g�5����l��W���%]N��>v�Sj$p��
���D��L~z�zy�&�ygI�l^#a�B"^Z�D�[a;�b�7��7�P%�M�f*��˛�P�&B��{���(�=�K���S�O%��
1�#��E��k	2ʣ ǒ�Z�f���$���1�;��-i�'�g�A�*��!�{��$�!�HR�����
M����ڈp�MP�k��1�7��O�&�,��q�^ɠ���ƚϳ$M��'hBH)2*�6c)�69;�F�`S�.)�=�H�2'9���ze)��b��f1�������(e#��AD����m�F�nM��kh�d��\Q�B��0o�P���_�C���bEQ6��#��ubl�ݩ��>�̠1��N(9�?���V�\�sL�����-�wW�/�K<�PZ��\�p���IךH����E��y�(2n\gʧ�����Ъ�e����:~�����H]e�9����=X�tZ�M�ՈX�t���:������B_�k��q8�mI��
!��w���]xDV��2c��pbQh
�@#`���_��1��㽙"ɚ�����Rupf֬bԤT�)�	Z�[�P���c��c~L���Z7:j��:o�!"\��q��!٫��X�o��A?x&^�Ǭo�=����H,�����?�ޒ����{%G!�B�vg��	W�am3�\j^�ݭ9�����j�!��3��T�#�{<D�Hx$#�GjsY����u(�P�]4U?�j��7����Gf�("�h���'7&�w1���=@�o}|�vJ��l��ؙ��y��Ɓ��
rC��l�%&�y1��w��*�	ȴ�D��1*dq|�mk���G�g���Aa�:��Ypp?k1? i�k%N忓�͘o��\�PgzW(h�G*�K�I����y}����Մ)W�
4��Р���ım�KrړynPX��mf�u=q����!�DBAٴ�j�W-9Į�!N�t��Mtf���5�c����L�h��OM0_�e���g #**O�T.��7�o��§���`�j��0��g:#TT8�Ik�o"��jfQ�ݒ�	��"����F6�7�D���vd��'�qTz���i�]�X�tI=ҽ��rԘ|
�C)c�@*��"�m7rH0�x�$�e�c�J�?�5���'�W�{�f�,���VΤ�ܕ&�7
� ��k�v)w��3D����eiv�������4�y5aH��ͦ444���opHh�c�Qk�W��}RGqF�\wX��+��ޢ{;끳���W�x��w���$��{I���0��1���a9�׫yȿ�#��,���z�P��t��N�ZI����ޕ:av��1�#��y��x�ŕ'��vT=C�	����y�~[p�s�辭�;8����	��c���y�1,�hM���`08"�Wr�1��_��|C�`"�#�e�'q\aV���F��vHҙ=�ݐ��l[^�#�`�	�z�:�#�R�P5�����=������Z<d"T-�}����lH���y�b�σ j��,�vS]Mg0%Ln9A嫟ƈW��d{�Շ"���v>��G�&0�A�G[F8K�>��}D1u��>q�)�[�X�6�؛���`Ey*�����(xþ���dV���{��9p�+_}��B[L�>�a��'�JI�;	U	�ԍ,wKد�O�y3�I��i�82>{U�|�E�{++�|O2B[���K���Þ[�±�Hp \$��[g|a���E��4��4�n�K�	B���q�
�f��0(�d��x��!��ɹ�R]��'>	�O��g��	q �O��]J&EVwvԫ�j~Y9��#����y]���G\�d�8CsI�m8��P�(:�I�ݪ�aPLS:?��I�ն�6d��K��9\��f��>,yE����v���u��#x��ܢ�a��Ar
z� �:ň�5+C�p�{��|z3ojM8ǿ�^' &{��h���Ik�P�w0�j�SNp���'��ہ[6��߻I-����T������odx���ss�N�-}UlQ8R�H�P�%N��V������p��wU�s"��i�H�� ��W
���f���vȻ[��rX���JGA72a�Ѿ0fQ�G.�$=�����<?��]��'�?8���R�R�o��4o��Ϳ��z��-L�^i/5�NW�H�*���4�` ���e�z�6TC]��e
���C-YU�A{$fwD�7l[��X� *�R7�J��T����A���d�
�WO���i��N�����Sf��'Cr*�´ٛ�,��r��(��ݯ$'�����^ɜ��Y;�K�f
�K���b���2�����DE�����T�ؖ	��ь���5��.��Wt���`��U�|�n������[F�A�kY�?�B~�.�������-ZL�<�phd�wƇ�A�2�:v�d��'L��:�2�@VyY��Ä�֌qRH\��k���ww�av;��H�g�'���χ(r��|y{��4QN�1�Rj�����R2��� �3at�	2V�?�;�4
�,*z���Dۓ��
n��H�Y�+�Pn�׉p
��W�Z�n�SY���j��:�ߺ�������BڳZ��LY�R��Ṃhˈ�E�i�̈v,�)gr����^��@+}ud9���1̐X�̕��<o�Xj9��5���Z����e��@�������'�br�/�$�A7=��dC��� �D����%ELPz1�=>�h[��du�U�s���2ikz�_���u�52�ο���F��<� qU��ʪz-p��@Hkv���jbb�ɗzN%p/�׽�2#�<g�ќޤ���̠[��0�O7F��G�#�k[q�/��ȸ�x���%�ɤݒ��(t��I�:vx�tT뛥�>Í�}�ug��o��;C��'�fm���
�LG�A�#��6�%���Y�����f�]���B��Zz?>�J�~�0|��d�N�E�:��*`��e}�H�f\8��<c�Q�@����G�<�c���І ����N~j+��.Š�~�>��K�R�U6��5��6��j C=���(D�KoI,˦ <6����r�q��V]i,�b��ȑl���<e63�A�e��� #��4�|�|��l(���2����ѻ�\�A���w����l8L��sϏN7���]%%h�����Bݗa�G��;�d�ٌ��ϟ�r��$(e�9���Gof|be��HA/��C�̠QR�S,>�����_N��m7�B����潫�CIT߸
K��h�T�m�As���/�B�����$o��j@;dJ�����Z` �4�Ȭ$-��2^���0O�6�GZЌ��p�4%�sq���c�-�}.y�|g"� }�kN7`��!L��H���}(�^������w'qjd q\��V@H����|��k�O�m⃋��o��]i���B�K�pҶ��c 12)���,O1��\K�	|q+�o�hk߀]N��aʚ3@A)��l)�Q�.=�N*{�o�x��d�zW�)=��3�\?+7朑xy�C3B�O%kn���{�
!�����e/�ZJ�����cq�R1	������y��s]0�$����m2����AnR$�E�no)�_��W��F�������d�$��fz�oZ�㒞3�tBq1 $��{ފ�}�]�κIl�`���{�x�.�J<��p���I�Y%ٱ� ��s$ϼ�~��� 3I�q{�����9�p�J@eц�ϲ'EB���"���ݔ#����*ќ�����bf{���]8>9�l��?v�S��o�����Zt ��}`W�%�BNT2x�-Mr��sFe@Ŵs�?��O$������qt#O�`�¬� t�ꝭז.	�U9Ҹ|hs�Gp�W:�`8�%�����Z7ݏ��~��E�Du# �?{�bkn�`�Z]cC��z�pL�n ��$�Y櫹{/U` 1됭�%^�q�)a�X}t{n>4�_p�7VO�fn���#�=��-���{B|wfVmv��_�j�c���(+W)(�e�9�NX�3�1hO�p��m}��d�?nj"�@苂�%.�/.٠���۾!�����"!J
�j4?�5�\����"�[�"����c`AǸ8�^�m-��ysxSԺ���y�[O�%�6�($C=���Þ�g�׾S���}�l.߮�����W��K���b��R�}�1]$o||�G����^Y�����^�#$9�BF=Y@��I�gQX7EyO����Jo}Jq����}�R&��aҖ<������9��K+r�ZNP�q�]�6&���P�}JYCxǡ��`D^��U�ב�3���͏ZV襺�&��W\�8���݀~�啝b���� *}������Q�׫�GLU�̎tKAo�i�J��6���0�OV�����Z6���m*�.�2��S�+�D�L.����8���pxQe�͆ߗכ�����*g�	+���8��gg�6K�B�\P-��������*D�gx��O[�rx�~z;ɉ[�6��9Y�VQc�}�>9>D@7���J7�?j�?�v{�(��(_�����g$+�[�JD/q�@��@���oj� �U��lH�.;e[� �_�<M���kzJJ�8��|��F�ć��]��0��C67�1���+�r��UQ���͜e��rLr���n��)����Z3�T��&x��j�l���KW�G3���j.��=�d@�~�<���!��j胈��m�̂5�c5��^L�t�4:#����n�(�@��=���5��D�r�hA�1s��:�N�Ž���5_���h�f~ !��w"[¢AƟ��fx�c�02�e9E��o(���n�����YR!̘~=���@��&J>{�����W�OQ?Χ���!灆�_i�AJR�C}�������O��������R���vܽS�s��'������&�������������&����	��u�F��H�\��x�3_*��)km��(!����4��c�=֧��I��Iı�,6HaE��LG�G�}��0�v�Ռ�#&M<�]O�%`���9:1zaf����W�Zym���K���l��ܷ�S�՜��ݛB�����#p�q�4Ѱ��^�JM�;(�"�!vѬ�Ɗ��t�g%Q����:���X���.挒� �S��`��D��sx�/d���j"f����c��ˊ�+-)����d����WE��3�����"�#��;�gg�.�0+��,{tۇ1�~�ﳠH�řM̅ F����b1'{�S�>��8͈�|$��OX����lt�X�$/^���s1ko#@غ\>��&�k��G��nLxF��v���s�[5PR!S��*
6Q�[������c�$c���{��d�[���:�Bs~Hi���B����I���ͅg\Lo�|��7V��Y���k��+/Yl�W2%���8�����^E�Xeb型U2Ϯ�L���M#��!��&6o�E�A~�e��@�d'������e0�c����e
t}Z	7��+�e��t#����oU��_��5���R�����]hݑۮ5����w4z�Loз�M�1��FCf�{�)^�&�ع=�d�<Q����.�'�ѽe^|B`.9��q����z�����O���\ǥu��jE���ĝp�%��l{�_O�QKE�b��S�Xm����QD��;�߁�A��+nlZSh��8+���}�Z��'��8���|P��Г����gY���:��'��'�g�'v�IU�m��}�:����"M�9�v���.�kc�u���o]�d�hܸ�
��z�`�aT��<��S�$�Ȅ��4p�����k]�ec�(h`Ŗ\��{r���1��i6H�������4Y)΀K��瀥���d��R�p�M<�ڛ��4�%k�ښ$W)rY�y!�r*ӓ�xb(	?0��ov|,�/3(���B�ѵ���16
�Zȳ�@��w{v�Ӌ���1G��fK������p�4)�y�����[����^�C�+
y�J7\#�%�8V�~MȻ��)�5P�~�Fb��|W]�j�����ﶝ��~%� aڻI�����p�4������d���)�>�b�/�mOt� m��{���ST��k�hÊ���/�褖 ���Î
��A�
�la+�H��5%~��N���W����ե���>���#=��F$�np��.C�wj��U\h����5���������'ko�ZTU�{�T1��"�o�F��]�`~e�Ĥ&UIiMA�sL�<�(�&��_E�'RQЇ��q�2.���ao	a�O���b�6�
8���0��o�r[K�����ڊut�z.�iI�`ξ�\�tF��F���9��A���P�@	�	�O<G&�4E�,u0.�xPt�!����'jb�@��/���,���Fb�_�I��&��4���A2X|��[~��������y�Y���Y%��ꯥ��־�5{7���q�����Dy/*ʡ��ykwy��7�Zz}<�~~�xv�)����<ӎA�~��QMn8\pm��-fI�N,ÛG�A��ZƟ���n�Z���F��JpuM��& ����Kϥ��[�e]ۧ�R]�ۥ>|dz�E9M��]��3pf!S?Ӗ��M��S�(�{�-�eq�v?B��zIx����q1hŠwu'G�����TY��y;C�]T�E
���2����Je�]�l��1��6dd����x��Ad\�ws�#)�t�$x�
�j�gW&q�#2=}�{!x$ahmc+�nY+}��
H�����(K�I1x#d} �'�=����DE�/���v�mBϡ�i,]�<���:;
,�\�!0�}`���^��`���v���p���g�uA{�
��L��9���b釞�D�')D��q`��5��׀�TP�t��H��ԇ�Be�j�|���\�H���Imޝ��j��WZ��KR��_�9Z��9������:�Ɗ���~{�hb0U���t_�0`.����|�&LZ�@�O��G����iC�L�aZ�n�7��RI��KچGs�%��n�_���{~tSkdKg��-�N�\�w��!�������Q�@c���^ n�i���'D�m @\&�
�٫	O��gt��Į���.�-F�ks��������f�[k�g�B�[.�n�;fa�;��\�KG#st~�ٲu�'ԣ���^���\W+�~,#�VR������{]/_^��X�Ť�=���Q��>V��Q���9S�a�}���C��