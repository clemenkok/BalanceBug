��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�M�>LA�����QZ�DE���	��{�i��ɮy7�K�I���9U����k��@A�'^�p�[Jr<#EϭԞvВ�w�6Q'�3�r��i�G/�����	��D/��Ob��,����U�*i��7}C@������ `�o�<�J̪įyg/+ݑ� �C���R�g�M�u��;��ѨD.�ڊ��Q�v���0/�S�Ѱc�B_�,�z�݂�� Mk�����fo@58�H�ɡ��^�[vj\�ty����%%�!��h��ء���1ӈG��-aQ/<ត/��q�_"��������d^���P���A32=�/t�V��!�$���IS�ݤT��s6ʻ"/1���L�ǥ�|��L��^s3�)����[��RYTn�;.欜�jNG~��OP�;�{e8mmxxMdc��`( �Hu��|��$�n*����ʈ�����K��3�q4��QI� Z���PߩܺD �Q�f� ���#�6x�nfзaУ�g8؃��c�p��.c�Y��B("lI1sՀ<�:9@�^y��ΐ��E�� =JVD�']��guj�����廳h���TR�p��Иv��MQ;-?ɋN��;�fE,F�!B�A�OK�;�ae��,�U��I��(	��2�N����y�脸,��!_ s�ȉ��F��D~���`-�e?�nIm�rJ�Gŵ{_�a+ h��Y��KԐ�u��1K�y�8TB)���{�F�kSm��m*��a�v3��׶Bb����4?�AZ-$P0(
l^�z���B��1G��pyo��ƽ9�ɺF=��~�b�����P�x�D>ܧ��`2�?�7��S�}"���]���O��t������v6�g�Y��oT���ђ8��*񞳷ʳ�ܿ*�<I�k��'-��P"!��#�mA����^���ZZ�K|;�����d]G;F���ĉ��O�k����V�?i �Y�xK��W�9Dv��*%{*6�	�i���o�!�^�U���[Zr�)Ø�^>+�BdA���C����"�����<��4�lwta�C�:}��a��9�'v��?�kͬ�z�u�vS]{΁�h�JW[���M?�E!�)k�݋�q��:�B��-݊���)¬��WE�.|�:�I�b���$�K\��8y��{hP8J�ׄq�-KD#ۮ��1�~�����ꐜ9J�P��Ui�D󩍽��	��\�?Oʮ�PAP���;� ��ޖ/��@�q�73�*��Pa|NX(����~��}MԲ��v���+@9�u�a��I۸�^ FidG~��T���c��~���p�+��4&��E�&%L�`Jf@q���bB�>�~�0 e��3Ag��v5��L!tz$3����y��m���f%"E�gY~ މ�a�6��lK3� ����]|7��-w�]��0��Ԁ��fX�>����$8'��"U������K�N���ع�~Sq�X�qN�)9柍UU)R�K;C�I�sТԆMؘ�{�E�Yn����!�?�^���+�㍈@�e)u,��)�!�p`�L`�D��.�%���Z��_p��3�p��S��Qjqt��+�L�`mj��-�>E�K���m\;�O0�
���l{��y�N�I�Z�Kɵ��$I��S�I�[ޤ�DM�k.�<��ɝ9t�B��)��|	�@�C�
�TL
2z���O���^�F�d�*��4ƸD
(��a~�i|,��'*�R��Kb%<|>D�t����J����2��~iD�����XS�@�w���<��q���Ao9b\A7@����NҲ�(ڰ5NM�{cQE]���&��P��/��Βg�gœw���z����Q#x��oh���:<;K��P騸�ا
ӄ�8�MZb���6ڨI�NJX�T�U"&�/�� -t��O��a�K .�ߠ���I����m:��� k�$w���<D�sS�;�w1:��x�6V���ѿ$A 
���X瞍��憟�MM�{�4o(�,[���K��x�K���z_f^�ޤ̫�9����&X���� r��%�95$�\MZ3Q�%��5��ʖDx[���1��l���$�-s[ֆ�N2^*�:\��%�T�z���iV���.XD�L��aFFn!xQt�&؁�6��Qq������ʈu�&Ь���WT���B�FTMSp���Ըr�uR�g����/)ñfD��j�a {>
AuZ@*���fM�O������];�!����%�<<<�Ndg셣��U.��;6PI�z�ף�<٩n�"���y���+W�ǭ}4�&�n0�+7�����n���L��p�=fwDƕ�|��G]L��q��<�$CY��o���d��ޛHK������$��S�$�^8�˅��#�~9oլ��_�����a�NI�r��C���w��6򹽓��G`ne������$DB�5*�Qs���8�Z2b�l�����f{\흙��?%b ��DgC|6��Vu��e��2�� z����v�@{�c{�k�\b���m�u�ȱ2}��C^*�������Y1�>�|����c"[��ǩITV���r��V@�w?���%+;<�����#E�6oh�ƍ�-�鯊nX1�(d�N構"]�T�{�M5����C���!����8��A�R侦opb��D��=����F��[{��}������j�#�������[E�CF�k�M�x�#���J��L��-[�[��˿&E�a	]W3�R�dN���;8޾C����5�};� �S'�H���.�T6#�����b	l��eB"��%����!|�dOh��i�-��z4��.sDƩ3���GC����W�4���U�Գ�"�{(3���W�ŏ��X+i�q��;�)����0k5�:�7D?�2����!��1� �wgIS�V�ZJ{
4�5�S��'�Q��ù����HB��|G̘P-bG�I�F/�ề2��E��x8�/�]�50���Z-���cHX�n� �i���� �1�!~��Tq��>�`�1H���-�G�22�K�!�N�2]�
b�>pu	M��y���6K���`��A?�C�E���fv�p`Xս �0��d6��R�ʇ1⅁s�}�8���'��Pv�(��Yտ�z�)���q��!�>wt�#0�*�\1}`i���U�u�ײ�`�-޷�����2���'���K���v:���J+��g[�V�xi�i���z�秧�H��ŀf� tNQ�4���r�`s؉Ĩ-�F��^��$�B����7�7�L�O������8*\�:E���iv�}_���OP��-�]'�	����s��ZŽ�D1>� ^������jTZ2�]>t�M~��g����̘a�/7|�ّt;Ϸ=?rs-���͉��*���Jp3���Y|���������D�U�y�uh�;��Oć^�4̼qHҲD��#�W���IŲ]X�2k�J	��^��Ǜ� {%k	W�����	A�m!�ǀ7J4>�+��$���XT�܅�K�=਀,�V�}�~3�r���^�3�y|�E ���X~�.�6��,@���xѧْ}�!�����i�$�=�3�I"q.�T����3���xh�q}�H����i����&�(���rk&�M*[x��%@�s���⏉��LX!N n)[i.iF���Ii�hk@V��r�N_]-���7J��.���l�b-/#CeO%w��*�}e�mm�-�k����PkC\����Oa�p���n?���yz�^4�����]���Y���%/�sO��W����emR]���Ab�+;F�w��]m���icF3���Q�\$�aP{pT��e��~Ջs@�s�?����ɫ�+�����}�h(�Nh�X0�[��v(��(�a���}�c�c��y|K㸰���Åq��.����>��3~�'��m8Œ5}7�Ѣ���bݪ��䞖��$���5�e��H�l�"6b5����`�}�ƦS��toNu7VЫ)����8O�Ӿfq�uR������l�|��5	N�)CO�K<5qm��A����J��JK��`�b����Y�j�|ߦ��[���ז\u�\��a�Zf^�j�x-y/��*f�|��o)(�O��h��1icT��[���&�/��/b���BvkfO�no�>��55oWC�DM��
�@0��t��T-��TRr��bWc�d�dq�T���=i��%����]
�b��;�KF��j<u����9=���v>|0��j����׽<�X��p�g�*����~��^����1�N�D�x�Qq�����Omh����uy�.����tN���^�P��z���È���pV/̔��r�:���s4#�0BM_��W��?HՉ\c'�p����=��v����$�fV���H��&K�	��KS�w0����h�|k(�5k6���V�Ǩ�=�����]�8:��&��U�m��[˼�"9c,yJKڤ�o�{����Qݺ#�dw��zf��E��aF���յ�S���|W7�\����ؐ����{��:���+���:�OԌ�aǇ���[^[�2�f�D?*)�g ۄ��g�T䷱�J]�l�j���6�����������B7���`�;��gW�����^�0A~�	��m�q5�rMo���d@Nܷ���Bt�Cv���2v�Q�I�|X�C�@����G����&�z>��>b�<�G���S��J��=�(�w�
��~���8)59mI���R�"��k@Z׬�n�3}AO���Q���Y�iЇ��V���p�jV��:zЀ�[Pc�<�h�y!�M�����Bǘ=�ͱ�:nP9K�O#�C����!�-��G�(H�(^2�w�!{��6:�FwD? �A�d0�H��& 0D!�o촷b��O��YAuj\w����O�����^ܼ�&�"I���Ȱ��Z�a���c��hu�oT�*�f�n�"�"ON��:Xa��r!��
1�L�����U6F~F\�1���gD#����#��o�Ң�����K���;�IjM�ƨ}�{m	�y\�����c���R���q&	�G3�g54g$��ϱ�?��p9g6����샹�����J�4�Ά�����5kOB�^1��DWla[3a `�xC	U�j�� �:$C<���L��p�Q��կl��cc�����~C~��l�gW�4��q�O8�(p�$�Q] D����4u�jA��K����簬��4���C <uD⇟�@Y"Ds��5�Xh<ɐ�w����!��eZ&d0�S?^�U�=�)��%�:+;�,��p3��������;�!��_Lk�y��-��ǿ3��AY����%��W��@�;|,�v�iXi�u�sϑX�QNw]�х��#���N��H�k��r@�Y!��AE*`�j�!�еe��p/�W�
���n3� �����`7�YYEx��t�VW��~Y�������(X�-��4���U�q��{�'�Z�=�i����M.Z��r��2	����H���MS����Ǳ"w�W�(�4���.�:�_���ڊ������A�'�+G��� ��_N��9��,~���~���,�?����ݞ���yZ���΁`�{䌟�'�W�*,�G�|�	�g4'�b�uy��R�Lz��?��<s[�q
̰�0� �@�CJl���:���� �<B��lN���2P������2�	����&�"�juE�[bIZ+.���H��.˨[v�������>enҚ���$"��Ui}��3��������������SÇ���,E��D{�m}�g5��`J#5�`�􇴴db`���S=R���2o��C(����Y
7Z�i��H��̹�6��n$kMB;R{�!�G�6� ���j������L�_)�&x�<�sֻD���'�e��ή:*�:;VɎ���B�ѐf.w��7!ؑf��6��w��u�/�c�����>ʿ�r⪷E�٢ר�^�K�-��g<SJ����ٻ��Ո���na�ϳ��~���o��Rx�R�5��' �a�*��]�9z��~�It�c}�'�Hv@��R����{i�A�P���POG�4Fq}�%T	��<��D�!V���J۸��j�"��|�^����Ս�Tq�:�����RbD��Ŋ�A{k��&O�2$����tė���7-�ۓ�<@h� m�;V�0���!���y�@�j���FP�
�lm��=7��2{���j�@��mo%�E ���従�Qy�7�^�
}B7�Wv��|O���k��zK3s�y���w��v�W�����*��s�(�?
�ϾE"�_F>uaYq5[�Q�`U^fhE�[Ɖ_�D��:d.c�Gb���O[����8��1��*�b��Kiw�k�Q��<�����k�p����� x=,[�VJ�y֒�D��ָF��?�Mo��Bu��b�w���� ʽG�}c��=����-`<p��4�d��yMnY��0�	o܃��ja�(�H�+��������3����IP=\~�v��Z�'n^O���ac`�㭢�퀤�+\L�2a����J��W�r�9�`�$-�4���ye\ʚ��p���qI�������Yyҧ����`Ĝ�S�U3y^B,0�ۗ�o��8�@�L��l��g���	�bb�9/h�j]T�Q�V�
��[����!k�X׋��YO��7�d|"�H]<���.H����U��ҰD�����!�*�~�
WG�lK�#,�x(�Dܽ�  �D:��3���%�H��!a��P���'�|�i�;�%6u��� ��
�jrfb+�9�[PM������V�-�V�r�h�V��K��P��"?.��D��岓I�J�2�^?�l�s\%g*x�<��wA���ha��#R7�(>�	��"�6"@��U���p%ſT'^�zb�p\�.hw;����G�>�mn�_5���1%���(V�Y�a�{��)�au�nB
�����������Q��U�B@i ��;K�>:!��K�kt��B!G(�V����K��Њ���'��>?S��ł����gmUO� ����v�N�O���!X	V��T��������vR>��'r����3��;���*�ِ5���W�l��� �m*Am�N
��@�9�]]*,;Q���Mɜ`����3	<Z���8Α\}�Ԏ��<�jdϭf(����숎�e�=d�mP��
��gy�P{��(�)�l�l�m])Rl�G#���V��7W�\�a�ou�<�x�V�IH3��<�w����I�M�!;E7�1�� �Vz�΃m�x�uvV��}7빨Y�yП��u���If�!�@�풡� Mz��Ab!�t-��YHg�ˤ6��%�ʬw�I�%��.��|�@kB�X�*�&�r�$�2�(=�乺	?�@ z�P�����H#Q��D�z՜p�uma �G�U��;��?������`�x����T��(	��xz��"�h�=GQ���N��� ��Ǧ}���3s�N@�V|p�Y�~�'-���p�n�B��ˮ�R]OԒ%O�C���M-�N���8������s>��u̧r�O�����C1b��F��
.���Ė1�N����i���VW}�c�+�b����{�9*Z��9��N��2�@��^b��eQx��2z�d]���G��zpÒ�G�(��}^�N��ϝ}��Wӵ�+ɒU#4���᫐�t�;�9!��^�%9G!����_�z��⨻�h��.�����<Ǽ�6����|��Շ>�cfw�d�~��յh���D���6E�GW����=��R�����0��\�"Ws5-dQ�K��m��{I����Զ��!!�#M:�i�E^�ӹ���$��<����i�.X�Ӵ�ޒ����Qo��J�~���ڌ�?���6n��}�C)�!��rnI[5�� Q��8�r�k�:! �$Ob,tb��}	W��UB����Bw�x�v�X��j(�mL>��Q�ZM�^��'�0�8��\�T�
'�>[2�	Q\S�[E3s��{z��Jd8F"�ެ}gZD��`JAJ��v�=�|	��B����P�&��Wi�V�N�5����	�����G�+Bw��4�TlE ܓ�]����a7���t�PfȄM��A8���O��nz�d�	��b�;X('�a�/b��܋���ٻ��Ϣ�HkD��Q_"ܻ�Qd�#:O�\a��S�#��me}���`�rȏ��s�YX|�
���x�{L���j����t��IF_�����7��l0���Z�@3 6�W��X	�3�:vo�b�� �vˤ�w��P�x38�g�>�jδ9���sQ&`yxǬ����3^r$�+�ǌ�X�R ���G�h��~��q��z�$�7K��_(�}f�&WVVy�-�U�i��It�݄�`.���6�'gϾXՊx׵L��&���}�8�0h�;'�B���d�ݲ�Fh�Z�@��V޴'��n�Y
!RM�����O�"�oKh�觌�hA�5XeT"�xc�8����_.�oe5�:�l�
bzund��S��ʊ�t`���h�0UA��.W�Y<H�M�0���v���Yɵ��&-X��eM��K���݆I~j1 p�'���m��7����@���Ӭ���3����H;���f+�8����kD�2�}2�J��q��Z�*Y��r���p�^hVǽ&���Pumst(v�+�B)?�LEVU�g<�o�J�{������",t<kEr3�0nŊ��=��&��9��Ce�X^O{SjɃ�C��Y���)Gih�y��M(䏍���j�lmJE��)��K9�~��;ַlk�!��Ii�x�Ͻ��B��.{�|�q��Yh��2�E�tz
By���q�y*\\f���{GNM'^H1H��
l'��C����ߚQ���S�:_�j�"xP��,���@&G�ӓsW��n��E�n�܃�im@7���b� �#>/�������\�#�u<Hȹ-b�Ξ��e�HV7B����3�]F+>���
����0=՜��\��psZ����^��Wm_�B�8p�]þ��/�O�I���1����	E�#anM>e��6�<#܊�ѥ�nz�+�VE�@D�N����[-R+���N�R��KyK4dWĻ�N��O�{���.�ɓ��	״-�x�1*��
39~a�}��YX�g�>-��(D�*Ĉ�YQr��L�
����ޞ� 3��Ǻ_0;x4�����b� �W��]�-њ�Y�c����$b�JC����p(Ż	� ��-��7gU�'��]�BQ�Da���������&�R�,�s]�1��7Q|0���i���/Y	���RN	�M���ړ.HP͛�����ޒ2�bXT�h��C"�s�Sɗ���BQB ���|�DwQ �S?)����/rZ͞K��gE��P��P�g�AGG�,׫f�J�%�?��m�ox1�����vL��X�J>�]�8HP�ls����gY���  �54�ѕ^�����Uyv\��!K�Q0�>j��E���؛���׊���D���S×P�9B��e��͵���*l�Gf�N����'��6-^N���ۥɢ��V��DbC�����h��Ǜ�LDP�Fm4��5��}=���QR�&c	J2?S���J���S�w�����Y@^�S�Ԏ�����S|�^���jZ��w� q��
=���s`��V�6t 3�~BH�vH70a���m�'�H)Ac"��\v$$�������"D�'uU�+��Y��+ ���7�J�=4�:>�����N�73�1��4f�	��<a׼6j��$�?�h�s�x����A Cslλ29��ȼ���6T���s����T��żW��k:���_��W���G7jM��M<dx��*��A�;-Ӽ-��:���:s�<T���/�T8�s��l�Wac�2^_�a1�oߴz#��^q�.�)����^�|c���4u�^!�~�-�@�����l+���`W��7I=�&QMӽϵ(�E/��Ȋ���.ā��f.����P����q}��w�O���u	�=��m(���w(J)��Vi��5-�%���8~P3M�1����$�Q~���W:g-T���q�D���r��H�6� �.-������lJ	F�-C��ZZ�ŉ��T�M�$���J��&��o^��E�����aQ*�{`�!�C�T�,ԓ��{ˊw>��JɹA��,�Ps���Y ��QF�`��}�˘U^h?���B��X7�CE���$^�4��#���J��%��[{3y��F��5�E����a?B
�6YR���U��&�R�~ύ�G������ f�.�� �~jY7=�$��]�t*dQ-/�����џ,y�H��#u��(n�_���a�c�'�qjPU5�I�h�����7���LМ���,��-������G��Z�I�w���/7�*�Ǧ��C1��%�)zv�m+Gb����X�#4ڻ�VB�2Z�&}i斈��a��Y����t���i���i;.LT\EJY�q��G���Pƃl:2�5��:Lm�J���g�n�'M�dZΐ���{b��ٕ應^M�����},'����A�<샔ۂj��(����ƫ��>��@����+�s.�Ds�Җ�2��0/���w��cI0DB�c�%�pn�@6�&�c6EA ����vP?�������WC��>$,��1�o��Y���������
錳DI:���;�:v�N4�X ����	,�P!�A������NP��4zvB~�� �E�.�s��iCRN�eY1~U9
:��9�+f^CjJt�im�<����f���#f��C_`��?G��u����>��;�rs�V@�LS13���]�=�x�B�.M�<P�<�&�E�;�=�:�7se�[!��������(�qt��J� ���U�q������3���膞,�.k���u���!EvV5R�h��ǇM��	 �s�TƘ���t�,,�Fٓ}���GJ	fR��4�}'!S�!���k��C�G��W�.]�_'|��O����/&)��,OvR��s�k~���k� uë�`��/��Z+��v.R��&���=S0JAn��i+õ�T�;@�bK�cD����9B�p�׋���������B�w<���V�r���i��jW���×JX¸b�f*A���R@�
�_��r��A@LcQ�t#������ReW�c��'���%�tAK�h�؄�6��>ə�a�r>���g�R�l���<��rJe߳$�"���e|d ��CLj���<&Դ����w��T�T��ZF�d�!Xf�#$/V�%f�c3J0��.`��.)cn����sXI4���ToE��+v��:3k�yr?0���!��o`WN��_'���� d�PeL��%��;���{�=��-�t��d�!W�d���������M�U�`e#����
S�l%K�Vt�{l�����O)����ᦌe#���OvEg$+r;PZ���e�����]��%��r�=`$�~q�� ��i��3�Ͽ���
�bV��e�ffŕ��OX �S[ <��QQ�r�j��9�^��~f�%yAHn�y� �~�W���!`�Ӱ{E~��/"����WΕ� �&n�o���Ae$�r���mI�K��}F`m͑M��"µΝN�	h������U�������������6��g�l�s=[�/�Վ���W$ 1Q6��]�>#��Pp�O���T�EE���kǝ}���HL�ѩ�T���(zC����*�M�2%UnYs�ҟ7Pp��gE�YCZ����T7ý�]f�E�4���Lb���`6�✧�Wϭ&�}�qfS���r�5ڠ9#�}Z�<���*˄\MŔۊ	�L�9�~!0��p�	Z@���Q��m�Ϋ}vȶaV�)�>Vz��e�^����%7T����K��a���J]Ǘ�,	����ܜt�,HH���:L��8RT��~�A,e�))�H؞�www�RE4��i���+tg���$m��$
	��q�>D�^�2R}?��yD+��A��fZ�3���U��r���)q�������w5�k�y���*�V4�
f��M{���,Y`����<m�D@�H;I��A`,8l��\7���XP��,�޴��_�t�&�6a�f&�1���7��zp�-�}1K����t$�]�
@����4=Ď*X�%��Ņ,�iyۥ����A�x�0�������7�B��Ʃ	'-_̵�Kp��z#�!�L��!�|��:qn�HK2���e����jS &����v`�PV�a{��/�������5O=p<Hܨ�&��=G|��@)��,�z&��w حG�E����/4L����|t \:@��;�tǃ��QU��nUI��ڜAl�D)���;g��w�.�i����� �ij����n��J-MZb
���GQ{�3Em�{rɚ���� ���s$ν���.{Oչ�툐2FY��m���`j��
��@銼�L�!��Ǩ~ �&fHL�+�� �풮�ޜJI��D�u�|��G7���aRT��X�i2��BwQE����K
i:��Dt��ǧ��oB7-���3��R)(�Ю�b���䷾`$�����7$����x�)0H�~6&���!6�d@�.���܊�:}������j`�m��XX�����^qm���5��	�^���sI}�Μ�d��ڳNGעЗ�4S\��������$�+�9��Si�pG�@�ST:d�g��'�����T"�Mˣr�ޜ>d�����#ӳ�PC&拾0�[�"Z�Q	����/o�d���g��Y�<+l�#׮����S�dm�%�}\��`'�'5�vX5I����G�&@��e u�7�;�U����1��Tp��+y6=��,ek���#3�!���V����G��b�ɩ�U�x�x"2)Q�"_����`�Fm�����x	U�9��4l��VH0��
�M5� ��
%��Κ��p�=�����\��=U4��4��|轹��6�&��;�͟j'd��<h���B_���^z��1~��aV����yu/�v@�9֮񟎕�A��B�{hs�����Bl����=-v��}av�_"R�_Us�tTDz8r��^�(w�F_�Z��s��^S�-2�e�'^NE�#E�tz�{v:���~PЋ*i�?0,�x�Djf�cߌ�.}������re!
i7M�f�}����0 +���=6�@���E��S�I��]��]�<���h�xt((A�̳�a}P�g�95��bx�r����>�$�P����a�78���=��gN��#�%{S�p�q�/�B
�� yK	F����:gb/旪�U��M�|W
Ov�>��jۓ' �[ˍ�,.;��>w����*��{71���qo���ьD�B�7ı��>��X��(ڽ�M%�q$l�y��2G� ?��1�LiR�q��&�f`Pz����c��b.��{�g����rJ+�����������Y]b��A `2%�?)�%"�)D����DfLM�3�Ogy'���܎is����Z���FR$�ZQm˦>|���ܚ���?z��ڛ�+�Pm0���O]��ù��rqH[���?��<��? ���>@(Y'Qhc�r�0@�t��@d:͔Z��I+��!�[춖�,hk�|�r1�vg�U|{Ky���:���Z��pM���l����s�@-K��."��dbM�6�O���m/�5����q���ѩS�jF�����W�e��knԂ?�8/��hM�D&���g���7湲��_�ySa�·����|x$������/�v&�25Ĕ��=mY
x�i�2�L����8������a�N�,�4�E"´=.������Y�\�2u��%ڋZ��~�Ms�h��n 6gE�1T3��gK��k�5qϞ����8�����\k���"ѯa����_a+�r��1k2�T@O��^���/� (��4�;
��m&��BA��ă>l��qNTm�N�Ո�'����͇1(����I;j�5�"
C4��!ς-��|�_�b��L�2���f@�
�\qI�������k�5�Z�$�|҈�
��s�:�q[N�ǰX	A�"~�c��2�����
�0
\�v���G�i<U3�L6s4���6=4���;��U[���Xa�2�tY��|T��,�_��%��{GQ^k���VU���zk��x�!�193���a���D�`�M���%��Ѡ�=��+��Ց�М��K��!�z�{�����4� �qn�[c�w�H*>��f��$�7�,�uu��f�Jٗ5��(�)��c�g�=�=��],>`�>����Ȕ���+��E5�3g���{¿�Ȫ�
t�K5
�<�ɥC�L����\��nx����@P���䱊ճzTIݰ+G���I�� ��`����0�J�es�d���^���{"��߼o�*Kmr�1��ɓ�Va!���3������N��!����i_~U.���Sc�~�;<��"!<�?��Z�s�BS30��Y�� �>����t}!�'qu%���d���P>9I;�(jW��'kۊ�n�o��7D�G�,�K�7k��a@�7�o�nvg����̖��0�Q+E�+@u/T{Q*{Ƴ� ���Nr���Ks0�!:	�1n3�=
�S�4f�cȲ���E�a( "�%� X]Ѱ¼��	l&b!XT��'	ʩ7��dzCl����(['�9n�W��0;l� ��G�2b47*�(�,����n8G�vK�� ��{m����[g�f&|�ٰ�`�ڏ�.m,�����J>	�p�T�^yɕ�*C�&y�8���ZD����O��,��g��?��t%��HwZ��cԴ��߅�-I�~��K*LX؉	�Mf2e?�~1�疒�@JekyU����1X =��כԥ��'�����.f	�w�U�=(Sl�Q�L�rNy��V؇a�L�)�a�0��f��MUg�m��Sؖ�q�OzH�����~RrsV��M�����'U9�K���=v�w�E�\���X��Sbw,SpL27��u����y\�3ٲ�	�j0R�m<�/��G�@��g��i<j��	�i�2�hP�d�G�K%K���l�����h�I��������� �!P`��C����G��'�ϐ1����V�(��{B-+�^�#]?��m����/qV�{�0�Ѫ?�ibw��P]�l㓮��4��Q_q�g�����$�#'��~ω�����]���hKF�ϔx��d�N��/q�����b�\5�} ���;,�i4ǊF_�d�����Iɟ���P$�.��+�=׽��\����
�o����tk�h�	��0HRrh�u��乹��������B�	�eAH&h�iN1��M_��	�Fh�\e�x�ր�
�Igl{���:�H��й������As��Җ7�)w@(G��� RW�<�L7���m���!��w`N����ݟl3���K~��" �0#�)?��Gt��ێ��&Ǧ2$G"7Xԍ "]Jɕ�� P)���.â(��N�2t4z���~=F���@�D譂�Y#���"ÐSj�'h�ZV3|�ؒlm.��e�qLϿ��mNn����}4�`���>!��q�����arQl�V!��P͞WGD�;& �B�Hơ��j
����j���J5ү�=��*\�Vfv�D��V���׉{����N�/��7�k�Ϟ����Ǘi)a�(ʕ�Q�f���W�"���2��g�&�)$_�G�t�X��ǾC�k\��8���|���g�g�3�ڝ�V�(�������/dP/k�?ǬѴZWzҭ>�-3%����b{���蹺�7��`�V��q�������7�ƿ�y�����l�a
!�z���B0k[�7�8���_0��c+Jqע ���x�/X���)�>z]���{��)��>f�
�<<i�a�f��K�2�%L�I\��d@Sy]�1��b:���IN�:��@M4�=��±�����G9y�wi���4}���e0�Q�۵s;��I��3��%�֑�u���ol%�0�Y�-�Eg�%})�!xf��+��[%��u��8l��k|��~n����,s�:���j���@�f˝��(�'�f�Bn�I�]{�fj��EY��zK֖��-"e�bS�����߈1q{� ��)R`������A�Տ��z���Mk��H�<fƔiO��Я��Fd������j����ǘ3��~�$"�R ���s��ڪK��8�c1|�@.EB�E5��ٯ��$�[��K��'��TRa��couc�e�Y']�9)n�gSk�XL���JF:�ԁ�uǯ�.
�Z���9K)�L�PЕ7���5ZI<�r)\P)��A{�qv�<������§`*s�#�T �E�ZD[�dE�/�m��#�����Q��1|�C+��Q���ߍ�acP�޼y&���FA�
ޒ���B����Q�o�i��3��6��vxYWE󏗙�2�@P��q��D��i�B�%���2��D��lJ/g�Mh��fR2k�����Szq��	��R���f�h�1��y�(��e��1A
bY����Yp/�[���1c�)*1�(�u���Y�'�]�u�>./�l-�az���B(7�6M����6��C}-��o�D�zT�=]�ҒZm SY�Q |��v� O����浝��L�KI�����Č�� �R�^H:tX�`.�/�ό����[���2<��)��(���d��c�V��u,�����R ��S�:��$Q@Ŭ�Ԯ��A�ۤ�������u��U��J��/���c=��[m?m|M�n�΋�e?�{���74?g2]g���������G�w�}��*�27�AN^�s�X(1�j���u�X�=�:͘ь�%I5��6̈ϭ?��+���`*�nU�<o�Rez�\�T�3�(��q������=/��2��Ǐ�g�{(O=���=q�����+��y-����2ϳ��큡�����}oO���\d�Ԕ���n/����:�w�;���(M�`�Q�4�C�y�=$�K6+�3)lD9�z0g^ oY�HLG�G���~/����j�X�S��Bt#�x��cα��[���3���nأ�F�����nSp]��r�4v;�z�2���~�f�:� 0��@�۾瞼=R�F��!j�����+���b�g�w��v�8u\�ɍ�E�wk����W7)�s�^7� ~X	����2���T	�~��zPҎWS�\$��aŢ���#���4�ǘ��ku(+�Fn�G��Z~�z��C����m~� T NdG[�O�W���ݜ�Z7����H�V�}F�෣�!�b��MҺ�\�L���iu>ܰ�2�+T:_� �f�RS�[����$t�c��U�Hd<����%�{\��y׊�����!��JV�Q T��s���,�|�Z���FJ��4O\��nv�+Ôo�-�[�x�Vl���l��f]��hh������J�Z!0��~|lc=:�"�A�g���3��J:�����mJ�Qb�c|�:���@$-l�jŢ+V���^g;��!�g�#���L���hK����/��&\f.���1?èB�xW��!�� l�|�����:��i���eV�z�����	C3����;_���^t�[c��6���ț�����
N�DY�mNo�Jraa7��B�Rv'�+E���.R��V�^�a�3�J� ����u������sa���ίדQ]��Fm��JA�Si��@���a
���8@����FƬI����\�l8�:��gI�����r���������vh����\�GL�P���c�v�R���R5�D��%�b���Xڻa4�ۧZ��j���	����4��&~�F��O�[�(���$�M4%Q�2�v��78���뽎lNA����s��Yݟ[�:'eA��	��7�@�1V�S�y�ҭn��������fyᄤz��4��I���$1RҴ����p�|��:`�d\g��� "_<���R�Yʴ�H��\�eF��I�~���4�f~3��+g�A6�9��̒Y��2Df�5�3��}r�z�L�jCqg�0��I��?bV�]p��S���G���ڐ)^�]>*�����|�8���)t�Ű�q#_�kHh�-ۏC3�t0�j����=��h��YJ��+~�R��Y�85}�s�nL���c��=����M����4c�߃Ěc	qCM�.�נ���R�V��Yr�*(Uhv�n�hbI�˕��z���R%�!���^{���[-Ui3]��(��oiꀴ&�S������M0f�^8�0C�da~�Dٳ����9�Gֹ[NC48�B�`���k�c,8� ��WR�ʵ4�?N�ޝ}������}�QW�P�j��x�[�e��b��G4]�?�؇�%)�rBf��c� 3�W��PWl�O���#Q���������O���v �<'��:������Ҳ��kB��M$"RF��Æ]	06+b��]|z5 �C���%T�H���=�BE7S�%0G*�7p�Y����z8�)�TI(��\%+ɬc�(u��T&3eSK��r_��0k�|I)3v4�l<" ��W`��?�?+�H�X>�kwϔ���������1�X�D9.�I+i<�"0� �a}���E`e����c�@��&ϟ�U�`ޠ������k��A�йf��Q�j)Q����e�a�����7���it4zէ$��_Q��O*V^ǦC��جŀXX�	�Ћ]= 
"������n.�>����N;�� �6!�h_���A��]�c�4�4�3�bٳ^i@���G�v;�Gx��h�S�܊])@�r픁��W��z�v�H���bnGx�q���wI�@��݋�Ĩ0�,�9�ĘĀ����D=��[�Yh���!����V��=-f�_E��:Kg��#�B�d2�^��4����:��&B�}3�
|ޥ*���K ʨ��s���$�a�.�I���	��$$\-�����4B�4���^�Qo�#F��x��I�
݂,���v���bq&~~�ct�%ѯ�P �֖�gk�~���+�T�;OE	��쐔��tA���	x^,�K������V��S�wB%�j�a�һ|X�GA�0�g�bsO �c{�p�N�UCU��T+=@ݚ�,{�kH�l�9k�զ�iNH{�Gz��ir�W���Z@����ה����ͣ�I����%������H�-"�*8gVV؛>�a�$��%��`4�a���d]풌~Q\5�C+'g��G �������G���*[���*�h�5=���݅z
��D��><��O�u��4a�� F�D2?�ͷ�M�U�z��ٶ�E%���<������e�F\^��61��s��+�x�p�\me�>C�4B�(��l_�8���9�g���d�7�q��E�����a}��69 �qO[ 8ԛ���3�����D��M�5���`��$B㧓�:Jb�)x
�,l�V-�xw�J+�W���PFʹ$5����ɮ�R��#m��I�A�o�x'P�����ٲ������/���chbO3@��"�w����uy���J�BA�rcEY����Q;[m!����qc�����0�]�ۢlH�wjs�<}�p5�θ�촿�F�%�t�URY{�)�^��cRC�w�R���A!�v&�-oȆ]��om�� �s�!=�&�B�C�+� ~�sGuסXd]�%h�eY����I-1���6 +�I=)M���vS���"�Rt��;I�ђ�w�G�a՗ޱ�h1�6�s[��I�ެ��`A�R��L7$_�|5J#j�\�#/�ྫྷ�%oι���X�^�rY�r3������8	�����2���p[�iL�B�Yhe����&5�9�����d�L< ���HO���']��:z6>KhK�n=U�9���<zZD�"O�;����^�Jj����?�l	"pk�*� ,}�8৒Q��7�_֧kP�eaC~�&���Ǻ>��"`)=����P��^*x�ߕI,{�,'�-��_?�@|�Zk)����KD�Z��]:���&�r`�K)-��ys�2_nO���u� ���z��9��+����* �Q� ���^b|c�Q�J���x�)�}7�Խ�1�p#,BF���yء�W;�j�ޢV*�9�ƋP�cLW�����:n�� iіJ�wů���r$6#½<�o�8M�$���XrJ�q �,�$c���SX��V��6����i#�A�œ�@�i��ʦ�3�,5;�X��>+��P�U�4f��wBX����~�O�gM`�Z�G��#3�:8��w��������%��
�5�*Ia����l�*���Dc�.�~����� ���7�6�s��*��12���R2U�PkeЌ�S��t���ʀ�M�uaC��:2��`��M���ۼ2YX6KB�}�5��B�B��?��%�*���֎^��9���Mݚ&���fOǤY��y��H����~1�k=�_��x>���Pй�9d�N�k�P�����*.�k�� �F,F����ၺ� ��@ȖV�[s��)-�6��eܩ�SH����P��b�OpH��t�V���.�~�7�r\ �$c�Y�Z���sS��@rT�ʅ�@?�ߧ'�7��GR���,�m��#��� "��&�L=��2f���U81+�Ճ�!�iƇ�x~�B�v+��LW%?�p��� �!���\�2�7Ծ2�$��]�E�>;��<�����4s!��X&E�miiQF�~�	�yX��E���G�����t����5�|Mƞ��p�;��$�0�,Y*_gl�N���ϙ�$o�)�%�,�K�l3u���^�5��_���O%������D2�_S�cr���'�w'L����=�r0?�q����Oc���y	��`�3\M�DqA�H�yT��=�H��4j�x�,�Y���F�S��0�����S�;W�MD�![o��G���[�A��Al|;�� ��R�='��\��x�o���dW���1��Z�^�:�:M��,������'jC|xp$:��i��&*��}�������&`n��d���U�S�yS�w�1��|�]����L؊�O]��Z6��d�A��	h��Ja�Ȱ�Z�O��'�/���z��"���*wgx��$��!�2������c���6)��G>vF���R�>|Ѭ�0+�=;��OSM?�(,B���	�������[�Cg�m9��@�5,^�J?yh�a����K1��B(���M�����;�m�����XF�<!�3b�q/�D?q�Ϻ�bh!9�KU,���f�mHQH�D�j����/e�����5�,��"���)��Z�^m����M2�K�e�56�㍄-�ј�3�;Lk����kF:��{O6=	R-y7�K�0�Bi��l��ˣ�Ф2?�qsa�Q^�%��6�-X�*���A�p��y5;c���kԪ���r}9���o+��=�����P3I��>]+��ܕk-]�do�.\5��1��Ӿ5�{���0@������� ���MA�1
���Wխƶ�#����{,h��.J���M�����5���>�GyȻ;�yG/�~������MA@!|��
V��h[�פֿ�_U/�M� �:��Q��%��Ʈ��%�I� �� �E��b4���NBs�b�����E�w����*�Hpm����]?�!e�]>"����a�'4��Az�R�g��������
��}�G�kE"?)[����(�U}#�6q:�J>p74�b<���?�.rh�hjÿ$��dFN�V�����*�H2 J[�3t��;h�g.9~O��O�5�F���A�f��z�6/�2k�jiw"��e?�)�L�����_�	q�l�,��y{�w�UC�m@641��W����ɴ�Q���*E�NtA郅�x�P��:����ⳓ$��J�q6����5�,��_-������R��fS�dU��j�:��Q�א�1�"0$�������1�#�jǺ�췢т�`�2�Lc�*�
�үL��������x�B>iE��s�d!Ko��`�>xʂ�*k��J�}~N�Q�	%��K��Thm� ݷ{j0���>xn<䘟�U[�ǯ���Cʽa!޳T��*���U���.x�����>̯U�N��Sȩ�.��
��S��h���V��}b=��%��L��W�%,?(����4;tUU:n	���ԟ0���u�A"Y���+�`eV �:љ	;Kao6���$��,Ŀ
�Ke4���&{j�k�8�	�����r{9�7�:��ӂ���o�rNۀ̼�*��ho|�#�^����}��>�^����,M�[(�[i�"	p7��¿�%`Ɉ2�×�<&�I�<nU��[�?�S����F3o�I�(�DT)��`o&��#L}D6�d�N:�v���Zx������?8�*�������C�ks9چ�H��{fHjF��l����i4����� z?�����ǖz����l$\�@�I��?���=n��W'�/-�Q��`��S��{SV$���/�S?�B׈yW�=x)����0I�OF����ujǗL(���}B^�@y#��8B�5VR��1�h������ܰ+�t���~��<L0\��q�N�o3�J�A �����	Y�ר-	�һ*\/W�s?�q!�c����MzF�p�֎�;	��%߸䣔���4Z3r�g|Z<��VW��-�s��y��D�d�?�y�G#��@~��k�k�����"|�wx�g�)[�z�����ҵ��;5b��
>��ZB��v$��
G�ԛ[K������Jy�O(<�dSK>ox��E��uYڪ����4���U�7k>��i���-�
oE>�K������S�wK�'�����6�!<�x�2)�3���;���ާ��;�{�����V���,�\-(��A�����,~z~��:��P�l�;��H�1'�T�P�M�҈`v/ �s�(Ǔ���fT��|��,���X&�жyr���l�%G=:��WI��5�ϥ:�b,1\J��M%�DP���yĳ�#��.Yw�h\�d�si���]�n�UGt���)R�u���J#*���E�չ\�kCň�uPqN�/z'[-��E�&��`���
��E����4���(9�9�1A�h>>Ba����3�Ț���}o ��#�
S��y܃۾rQS������.��}6/u����+3l��K�w��1*�n���Al�*ؤ�J�����rX��ҼG��\�a�߶{=�E^S���ؽ������g�t%��d��!��(z��$뭺�=�?��Ե��I.(�9�]���P9�f["d���!&(..b!����0*Ij;��!}p9���L��E�Ѕ�:04<�`������}R����Y��}Ȏ�1�@��Ot�>Ҏ^����b�l��S����4����)��+�Ext��Up�[�k[O�;�y��jN�����ƻlE�����)��h��(;a�Zw�A���d��7�K��CO@�C;��i�R�b���bN���e��Cx�([��{ޓ��G7I��v3��.}� U�I�4������l�"l@��.���0!��(I������<A��eZ�� Zb<�����x��L
����^ˡ�\�`�MϬ/J���TG����>m�7�Y.EM�ݠ�*��_���#���s��u�xƋ_f�`'d��{�4�15_����J����)��Z5wXg#$K�0�΃��{wQyn� �q�	R�dO�%�H4���o7���+���@P�|��;�t��6�`'=e�ea{[C�3�-9R��~��j!� {����VrkZ�T7K>o �y�M�gWH�V��Nz�̡ؔ�Ze��*;f��B]�bL�.��k0�W���l8�&|�R(�?�&���0��A�gv�4%,M�G���˲]k��;����ݺ?�a*'�G�ɛiv{n�bf4��#ZM5�S�$��7VJ�Z�TMǥ�e���
��WVµ���q朝Ū�'l����1s]�%��6ʆ�r��&1��o�&�)�O�ᮚ�)�F���_�o��6(��|�rX�Q��p�o2�,>��W �'�ϖ��n�\8�H�x5_=T��F'H8?��ɘɃ��r�ҕ4 ���ݜ�Z����/�e6@��H��JS��l���\^r�TS����h�O(«Č%B �S>��M��Cȅb�R}P.���.A�	����F�ad!kD�M�ݮ��b�G���o�XJl��x#֢���7LS�5xYH�<���Z�W��8�l�jq:�����|5&��TS��'���=�K�p7S��ck����f1����U�놜1H9���&�H���\�Xe�i�Q����,:�@ ��^������#/8-�#c�@�3�� g����7����1w��(A�'��SP�8|�cL~(��Jt:r@����c���I%kyT�ג,zʎ�S\��bt�n����d���4OpY]�@����f���b(�,��p�?�׬E������c(h�OX�6����BЅ�8�yw�>���L0R�&����T٩�>Y���2�1��y�����E��mO��9�/��x��8�v�i��_�`BC�(�L�H̺�7пL��ۛ^Z�d*|�����:��>_b�|�Mw��b|'�
���K#����/��E\*�?1&��t|�qf`�ߨqN�����J�^s�Oܬ�ό���� �ˀ�&��U��f���1�B����n���B��:�qXm3y��M)+|	��:	?2{�٠���˄��׺溢ڳ�a��b���"dX��Ų$����ص��w��q颬o0�
(%ꨪ�C��T݄���m�#�8�ِ ��;6]X�-$TY����X���V�0�s)wzv5��>m6z�j�3ɣߓ�L�0�0Q���g<���@��� �Z���gE�tKA�`���$u{�y �P�A�\3)�����E�%Q��YB��q�g�>�򴰓�5l�_*P!#���[%��Z��
����JiW��bU���X�^d%�ؕ1����� �b$ȟ�]a�"Մ����sQ�p�]E���§)W���D�Z�7���;�����{ĮӖT��Ŏ���^(Ҳ��������@Ό�F�$q��-L~�*�F�jF]��^XDU����5��-�������z,����y�c�O}���FJ+��m��Y�:nʹ6lbZ��]J�.:�W���òW����$K�$v�T�Y������
E���h�+@#����q��Mɽ�˱����!#I\㼽���ǻG�y�n�����`��`x�$�J�ç<r=[�k�bKh�4��8�Q��OlP8l�e�p��+~]Iq� +�f������X��-��ŭ�U;�tGi��H���cB��M�cBs�/�`����-�2Rw	�c!�-Δ���C�ۢ��e-�!�\���-2�vc)ǻ�{��q2�Y�jD:�|-O��<:O�tכe+��C*��������������Tx~���?sʧ���z����W���ȱWK�(7��t�["2  �Շ���{�E���Wc�l����J,5��,�Ԗ�6���Vh#�`�㘎t�8r���'��d'��wOl��������$uxY�,�ڬZ��v��;|ૂ���W���9�Jy���/c�Bx�<"E�E,�jEG��;=� �Jz+HZ@���L��	�-V�<S�ٌ���%��^o�T�O��A�{�^2y�Nf�g���9�owW�����!�׵�x��D5�����.�xL3�L	4{��gV"����^����ß+5��1�t� �ݗE�Wee����`�C�n^3��2�`���1U����I���6�H}�P���@/�*Z�4{�y�L��VK�l�+�F���,� )A�)>Fc�O�XQ"�J�]OF�.#KR���p�i4o �HyDQI`�d��1����} ��D��Y
���c��״��XH@�u^����@s�?��)�XT0��^���ÕM.�?�׎��;���+����eʯ�QBRԁB��c��#�%`��o�yit�)�hX�����[+I	@��>������"��H���>�HN�.�c!�P���a��2��!�В��K'8z��A��]��6ʮu��M/`2�@Չ^�'���sqt�X�,���*�p�+�m��S�/���:���O��8�6��'�{D����{�r�w�0�-`wm������c��"�x5IK�q� ���r�o��sOB�rXU���AugJ��e�g�<�@�/�w�]���r&T袐��#��fe� h����g1wj@��:�_�Y)m�\�-=E��R��L��]��<s���K���#�o 5�ԭ���f���Y0�u���L�۩�`c��:-�@�k�z�����E)�ñs���C�-�p�0���Ɂ�����DU^A�M#�s�0�3^~e3x8�����k�m]ۭ��?Ϫ������L7O�>�>Se�+���*krȼm&|�Bܵ�@�Sĥ��uV�+�9$}@��,�]4�N2o��&���~�eR���]�{ay��]hR�1%g�X���g8��#��ĳe��MH���,4��!t�W�L���[1����,w[Ce�U�V��� �{��sR3���8�T��~#�0<CFh{��9�F+��-o�:(��|�حT������K�'�{I�rby������v��`��h4)ޢ��A��V�Ъ��Cٔ�@�h���W�^�Hb�`V]2|4��sbWh����l�2�������̮"�(���G�����O���yu���'��
��4rLP &2�J��5�L:P��n_�]�cp!k� W�5��~*���I�n��p�SMG՚�Ο��:,:��n�8��U�j�]F�,���	�JN�nT�V]2Y�v�7ۑ��[���w��,6��oټ�ֲ�}�Fc�u�b��xx��/�;}�߬t�}8͢$�$��^�i�I�!���ɠ0�����3hm��Yyݢ�8��0�M��oW'��7�h3~Z�X�O�/_Z��DK��;���Ǹ�.���!rO�+�X��"G�ȫ�Qu�Sp�𺆤���P�����.�P���~�F�|���6~s�:�{H�..��n}5M�MmXM�2�Q�v��ע~�m8�v́�TЏ��=[a����Ӈ����wvA�,bKYqGh�(�1�";����?G��*��1GЕ��F���ikj�_iۥ��v��ߵ�=:U�4���eW���w�鸃"W���n�h���j����&����$�� @�R�!�L� �x�X<�/u����-t���C��P����ƕ�!�ؑ�`�
2"{,�L*�\%/ �hR��&+N_%���N�}��}�J}~;Ҳ��D��D��Z� #��je���G�I%��t�d��K]׮��;��1g�f�L�Hf���7�jZ�h����0n�
�q ������4ɞ�'��80v7���/\&��G7s�fR��c"\c"�׶������4��Z���ޢ��w�e�Ef�b�;V5({�C��A��,1�sV�v���u����Q�sp	�:���i/A��vhm��%~�j@�'W�@���	�Pōa���§1��s����Π� ����!c���3QY�20�7�+b�k[c���,e7Y�?xsj���� 8P'������9?� ^U���y��#�#�>L��O�ζ���kyU`S�������1��A��p���W¤}!�7�Gq��&��b<j�V���D_3ev^���W*�y�r����!�f���Ғ��0�n�ǫ�w�2��ւ=$kl���6����4��L�kt�剧A07r�ӫK!�E:|����Ÿ@\��rǛ��noi0w'���2��(����^�����oa�	�À�� Gf�L�;��[�M@?�xl�,�v�ٸ|�ȿ 1�VJF=�C\�U�&�����;]�E	V![5��5��q�Q7*� �����@O6=@�0�Y4ʀ&�����Oj�ñ1#6��i{zNZ���3JH��4ջ$n5BW��}'E"�cُ�?�8=,0�$̦U�����f3���$��qPFllL�9����,�WC��^G������A�>M�V�Qί>uℌ%��#05���;K�E��;.6/��&�:-�e�U�IF��{rW�}%v:S�ڀ#���o�~�
�O�oqgS�c�-!&�G��*:f�ߴ��poC�g����,�\t	��z)ѻ�] �/?+h��_��"� �w���g1��� ��=.�� �A�꧆!RG��_���
r,�?�5>�-Va4a��>�ZX��$_���^-͢���(0�!6�1&9�+�LO:�qS���	'�zw��|�'i�����NiѶ���e�57�� �6\�:��kP6�Q�~�9;��v�l,'��[��YܲR�(ȳ�\&���Bm�8�	��L�ZП<�k��!��"o�4�jL'�l/�6�3*+����Е���]uel��HI�{�Tè)�V�*�NM���NY�:�/�r@��,^y���AW������6��&��P����߿���9��v�h���MKSˊ��̜���k��P��jޗl0ܢ��j�*��7�H����ΫY��$Q��>2�H�BA�#x�X�r֖H�w���v?j���6�B�jW��@�uY*}���muA�~FM+r>� �����-��ѷ�Om���_qD�{�39I��/���1,�H�Ƭҙ�?;s���Ug�@H�+s����@F��o���j�=֏M)C7	���c�xYs�ρ�r������Y���7'%��D.���o������R���?ǸeQ��|�Ü�k�!�8��ː��M�M
_�\fAKń�c���I�n��^��#F(
�����-#P��$��;!%��.�`��|�<6���"�R���[�-�q�,p��[��SO��B>M�����`ݟV3KpP�6��Ȱ�D��m8{ߢ8�[*z��V��J�ۧ�z�苆�n����/<����ʴ}����R�����</l"n�S�є߉�=2h)|c�P����P�X�*�?G��b�b���9�����A(�8�0A��C��<Lu��-zV+�/�ȃ�l��B��`��O�IdB�ǆ��)�[�~��-��������8�Z�9�e�� pT5>/`��ub����6���_��MhX{~�xr�j,���a����o0w�ܚ�4�݊��W-��r\Y���P�'q&i�/%T
QTS&z��ߪԛ87��>*��rJ�`;h!�Tm�A	���Dkه�@|�$��{��ߦb@!����TM�B�jv�'���d�\h���ѣT� =�'?�/L�o�1���� 킽Ϋ�d�t�ً�G��L�C7"���Z���<�^T��a
��if:#��e?��ܸ��N�������jQ��쑢�k��g,�"�+�*�������4M`�1#1�S6�II�^����'�>�XW{[fX��';&Mfu�O���mSIp_7���Y����c�"�Y?W ecr����po���'	�/Tΰ�K@`��Z�T,�H�T�Q�Azs�F�A3^J1���8�����i�ԷS.���7�q�=�gG}����+�){������y�q}K�!��M6��y=�g�]2P�MPzW�2�t�n�&�3j�ʹ�=������"F����b���>}�=#,���<��"ͦ��9a0P�yx�n�U��	�9�W
J�u�D�sޣK�[���P��]�OV<�BP>'O�ɏ�$
g`�5�0ʼS���5���bs���Q|W�O��T����|[�/l ���l�w/��0b�j �F���9�d�t�rt^�Y f$�a��q��b� l�Ĭw>2�8Y=y'�r�[�՝y�� ���I�N��U����Rң�&�l�;�/�u"�05I=��,kZ�1ڣ�{��1��d\MN��e�(2(�2��z�=����$	�.��z�g�.�60�X�����Y؜w��5�7ӆq�^j��i����Ry��U(��Xg��d!�5N���"v���7FZJ��g꠼��b
"�{�x���G>���뗫!�N����f5ż��n�2O�֮���j�u=�����P%)d f��n�(��8�-5������k	 f�Cf��%P^��:�v����$[
��#0:��TSS�{�(4�*�K�D紖G�{�`�s���wZ"K��;��d�r��~YW��>V��wV&9��,]��*$/�1dѶ�Q���? >y����;�1��L�¼N����Ot�Hp+�V��2$��zГ�q[,I/N,[�K0���uQ���_Zx�;������t�Jy3����Ӱ&{�T�R����"��o����[�ef6�}M��Y{UM&܎C	�*�u�S���t��$Іi�yi�!$�y�*-�	`���<VK4' ���~S��?գ�X\"d��C�w3� $(vl�D���#��EئD\��Ȕ�Um�����YO��/���Q�����Yc��Y�kƠ-��x�s,�� }y� <�A�'sG����@�F,�MQL9N:��̎JHR�DU����@�vȘ��=���_�d�dO�G�R xR՞���P!<^�e��H�\���۞��6JHǳp�Y���0y�����~�m�����2`�4@m��.o�0+�u���(��
�d�� O8i=�7��S�QF�q뙒E�Տ�1G��X������a����zp�L0;�բ�W��	bd;p)��ϩ��/���K��hm��1�*f�rzQ��B&��ۉZ/�x}�~1¿��+120<�W��K�H�	ݔl�C�l�}Zl��o��k�gGW=���ci�`1R�]����BIظ(����x�|�Rx>ds��f[y��&H�����&0�s&urƕ�7Y�dqa�ds�~����P4�B������(Yp��^Է,�9uNE뮟q��ݦơ~�Jv�54��a����p�l!�!MA�UE���՞���=�6��#r�1�[�/���`>K`2Tc�~�S�.��T�������G4 �^ ���̸@'e���J��!�>֒-��v�q�Q�e�ˈ{��ypq�P>�~����f�� W\���M���dp\�%�q�m��TQ��\`v�\mܕ��������'��ܹv��i]%�񰜵J{���4`��=�'�ӔM�0��4��~�n�5�/�
��+�� h�%X���$�~gy�|f�D�E�K�k.>�x𭼧��Ի��|�2DF�7��g�R�ߛ&��n�v�L����O�F�sG��&��kH�����l�j�S����I9z[9��G���I ��8�]_q�2���	>Ji6�����"���&��j4/���d-h� �6���h�Hi�<=�Y>J"���@c���	�	�f.=��'WX��o9��������&�u��S1�~�)��r��q�%��(��kp�z��2�A2Y/�й�E�Z���g�i�#�]�C%�Cy�K'�z��kK��̞խs��ɾ��`�̎RC�0���9O��4ܥ䞔}L��R��`�[
�LM9�	�OS�9$���J�D0��+�՚����7���^!@��4��ஜo�b�F�4 �pN޿?�������Ĝ��V�i�h��Hŉ�A�ތ2&	�ȉY���[� �J?�Y�V�H��Llcwl���L,y�}� ]|�����g>������ֿތ�8̘b2�d� U�Z�cúcQ���39;T�TUV���}@�9ї�{���Wl�9�t9]��M;"-�6i$4Ao'��=���^*e�����~e-G������>�"�s�U9�o�G/��W��Z�A3@qw�w�߉���O�x�$ZO����ő.I��ۙ��ʝ�:�� �`�������*�t\tc�1ѯK o~(�蹤u�Çt1�)>�iKLv�����s����ù0����D!>�T0��v�ޱڮ��� U|t/�AI����ُ���¥�:<j9�Dy��q�Tl�r��!s���@n��w��*����nV�.v���U|h+avLē����R� ��}_���͘K�"���+�~\����H�7�R~�P
�*��Xg^B��i	�AO��6t�#��|���f��#vU>�D�Q�γ7=T7��&�	?�6e=C8�MoV0v��=�e���L�4s�map:���g/�e��[��ތ�
�����ya��0���ha0
N���bz�������-څ.�a^!�q���D�kO�_�طʉn������g�қ�Mʎ��"�	�{r���&|�M�v̾� 2���;�8��Ƿ �`�ALp��?:�|5R��P'�#��~�%��n�U��S�qX�⌨;&r�^x��>��y
yg��~3"f��;�Bփ�40�
Cn�O��$�z���/��i�NmP��W�����?X��)��
%ߔP�o �����+�[��:+�	(�*h_�� �:�qDT�Bˉ6�DO�a&�ݫ���k(�-��N��$<�K'Rq���3J�M�Ug
;�c��1�����Ց@In�B��x�mI�;��}OL��Z�R�EΛ�'g��; 7�*���X�e�מ�O��w������, `��⋏�k�����]�=.�i盀�2�z�K�/��~�Q����B�����v����kB�^�@i����L��Ё<�<pc>u�Pt!nL��{;F�Q�����.�"������Ͽ��1@H�Elx������6KK�x!�u���{��h���ŕ�WKH�f���"�!>b\d����8naJ��u:�m�N��ϱ_�/ȉ�Sz݁�9�C����RO�]�!��&4��ɪ��6��Q'՜�r�+��X���ӻ��Sjz2��U��.H=�܈J�G�wF�tpQ��ϯWO�ULf�`m��@z"��9AE�8M�潪�r�ޝU�?��w}��}�pHVs�h~�����X���:G^(T���6��V�v��>�c�����`͈"����R,�=��a������	�g3U�i[��#�hfb0�B�.F�
��X�ht�
ǈ#T���f2OD�fN�wv�y|e�^Z�4I�SH�3���F�m���3A�-@QZ��������@GW�Ф�!��ݚ���G/�6�k1�H����^[�.�Ӧ��O�������i�N,*Y:+�؜d1��Ĕ_e�$�,�̻
�Mƴ����I`���&j�����ld7�B�>������Ue�q*�#�����~�CM�AHU
�\-�+x�$'R�B�F���,� �̻�,7��۠�Me�q�Ő�$���<�(�
�8�ݛ�!���;�V��KSDf�l��L���@�f�^�5kZ<�i��3�͕Wr�qvr:�3��XF�9�B�%���_��ݗI�:w9�`�����dL�|b�I�Zc0���gm_R{dq�D���An%�a��@�pŒ�l�J�p�G(�X�6xX/ue���.3Jx��y;�T����ތ�ߧk��\�����;X�A'C	�ꌤ�X�
���������tv�U'�Nkdqi�>��Uh3 �۲K��������"�^�^���$_4� 8Mg&N�kMO|����ì�� ���Zΰd�_Z���o?�
����p�����^��l�1S|�(�1���r����9�Ҳg���:㲈�_�1�l"u�w1Jڳ��Ĺ�T���c�q��O������
�1�����?e]��>@^WG?@Yn\���6=A������l(�1a!��2��a���*�'�����9F���mx�6k�4t%�������	3z~����u@Ҟ|{���a�Hx���ʅ�-D�y����f�|ϩ�$��]�!����q(eIC�82��ql�L���e����Vq�l��y���?��%w)ˬa�v�Ft��i��|��x����rM�E��5m���}j��:��>CTUKa4xz�z��W��U�b��.U.dX2�4�'���S֥]g����=�^F����x"�)_q�?����{}�	�Fh $g�3�����U	)�0`��\.�0�aN�v��.�x���i����DB.���
�n�J�k�yvZ���)�ю\ �~hUIQ<���%*��G녕W����D�㽟�;�l��g�$']�o��X��	�x(z����?@���4Q�I����$�����)�|�j��{G�������T�Ed-�K!%`��U	�y1DiFAH����C���n6��6�;j��^�+S˖��Dz���- ����ƪ�	x�5)WB���h~?Ha�������Ə�Hһ9�~��\�rǆ���K����(���!&�ٓ�Ӆ��(�:��%�"��rXH�|U�@-p~���ҔE�F�F��EB0EIEh�{��)��`��l���M�ew�,�����[7��'��&2\L=<|�+/ֿAW@i�HB��{�_AU�=��y�%�oB��{i��p��}������� S��'������cB���S��T��m�p��2g�����U�f�yTS�Sw
��w��	+)��C��uI��-���3b,��.�%�~z@�aޒu�0�T��z�<�lm5
U�vK�6��P£�i"�3�<<dp
f���R�z/3XV��8�ݚPZ�j =�P�v��و)`9���+0lFS-:�D�*��9�$�w��;�'v��2�k�r"�A���6�'��H�
AP�Jߡ3\N���+U{9����P���1D��Z?v0G�L�p�)���
�ޘ_�SNG�`���F4h��n�L��*Q����q\������jRC�癳!Ou�5�\=�)�����ͪ�P�{/���.��y	��g��)~��fI�&��}0�b��R�v#��,�d	���:+m(�w@�6�G1��d[S�&~�M�P����C���M��Ʊ�٫�S�>hA��E���"��O�D�c������xx�ͭLf©�PyD�lZNjH���#��	�]a öo�Ev�O��*.�s/˹�b�4���cJ��$��D+��[sP-`�c{O�x,����/$<�)�X����z�E����89#�"�
R�(RW�Q#
�u�����9l	�2ۄ.87�p���C���WW�=G5�-/�x�g����p���C8@ݒ�Zm�D�ޖJK�����%r��^��ϋ!+ocw��gIK�5����s�N�M�Uw����I)qwߺ����.���x�-!Y���,�!��2{R ���@Xɥ��G��-ۛ����E�����V13�vw�`�Y߿�0������6�"i�-=ҥ�hS頋!Y���>���y&����>�#nm�����	m\��y˲iG!E�:�{�Ɲ��@TE��}��cf��c���E j`�*�7(S�����3�T�M[!fp�@�.��h��Z�!r�4
�rG^������a���h1��3CקxS�'�c�D�?.`�P
Cz�:5f��wYJ&�a�@-��&=1�,y�	��������p�1��ݫM��P�A;�Tu��\�C���L'��j�j:b��s1&�T�U�\�O\��La��w0F�z@N�	]�t��[!U�Dۆ�)�u\�# d��	D�{��X�G2�^S�T��Ɋ�F���C�*G<˂h�E���Wȟ���U�DI}���	�Q�A����|&|lUE.S���~'H��3��^�o �L�R�s��jq�=pv�繪X˲�@��ed3�L`�@:�e�C���_z
ia��Z�)�|6� ͕w�����/� �\׼�5��K:G��f��+Z����I���k ZAz8�X���A�gC{
��~�(���;��'f<C�7�J!-U�`15�2�i�W�r$ё)��XZ��!�l��)�� �O��}�R�j=�w6F��̝�c��e�~��qs���ܞ����vŹGk'I���b
l[��Ԋ�KA���b\ڷ�6B[�LH�A��Æ�!&���*ߋR� j\zO�6�NOHl�Ss��_ǸRh-�}��P���wL�v�`��f�2PĴPD����7�K���e�c����=�%r�*^A���m�l~�ַ�"z�%/�KO���-�BM)�ģC�+���o(�dw:o<�꼄7���+z�٭&ZL�38�U�3#L���,�*|i�BP+{=+qjm���<TOKe���Ϗ��W-�l�N�k�3��l��(�[!��ݛ��>eg,�o8n�O�	�'\��B&v������%e�����C�+���o�E��X���V�V���\3��ei���J~�P�nz�j�o��#�4n5��o����L���	��ݘ~�8�ܴ{�:���.}y/)AA��b�(����(�L�֦���T����v,�L���*-��ܕi��/�D�	X=O����6N�<�WLz���G;�����۹�p��L�gJ�cC�v��:X�w۠O�ۡ�I�
I��|�
��=��G"��-�m���h+fWZ��o,�0����:pO��;�D���w���@t\����r��*)�o�0:e�k�jgJm�e�<�c+��Ij�c�X���C����C�� Z���:m��!���ϲ�p��b�vΰ��������״�`CO|,4h6�Y&�l��-��0^�ܝ���i�}�Â|�6� ���joUS}s7NLJ=i4�F+)���~����s��֞�V�C��*r5�r�k�"�_Tm{��@�u�R���y�}u���u�)�d�29�.�7�dH'r�n��� ���=�i�Gz����`��;a�ot�����97�۷L%A�8@�:�z��y8�d��ӓ�.�<�n�;�n~�:�%��L�5M�H���NQ�D2M�b!��&u�	�S��/�wt6���/���ڿ۴-~����B�&t����X�㇞&�_�'WM��^�j��F����B�p����|�š��[��i����b~�o��K�����#�`1�`周�H��8�-	֧����Ҽ��������&c�kQ�Q��`��XJ��D�tQ�K���������qá���f�CL��Z�@�3!�?��6��ylS�Z.[��}��ß�*~������f��S�
��7��wf�x��nJ�i�U_���W6�����*+��n�?�T��&>}H�q���k(D8FE0�~�"?�/�Mz�����7Дƽ@��w!,h�� ���V���S�T��}�<�L�6�ڧ�� x�H����h�ɘ�(!M���*�@������q�-���^����)��LP�ϐ3����.�^��HjΈt����5[?Ό��	�)`�_{�M�D|�Cx��4{Y�.�&I�lӷwr�C"�d4It�E���'�,O�ܛ�퐍`�=��\��}_(ء~�F�b툣*q1X~�ڟR���%�U�T(Ӊm���wS�{�	��M�*�}�HDa�HU-��0*���-N �f��s5�
��(v�\Y�v���*lf�p�v���r^�x���̈���r�.V����ܢ"|h��M	8�՘7T�3*,IT�k�$/�`c���Cnq��_��)� ΂�r�[U:��h@��"� 	EK�N~�eA��@N$�k�R�U���ފ�h}\rkb/!=��d�Z� ��bE�5 �WL�QOd�i^��3K3�s��O�_�#�`��TT�A�Yߋ�u
ݟ�E�vm[F�zT��MS%�<��Wrj���͖��g#Zޟ�
�Qk��ӏP"�}+0�=��+�>5R
dT+���[�R@`ǺD�����2�P�ELD^6�pt��1�'gY�'+m�TW\��ʗ9�>�+�EI^6h��ۛI���z�M&Ö��6,��� #Ҙۄ�V���1O��ľuu0c����-�����u��n��!�=�	�v5"�A�ҍ�֞�?�c6y2��Q�����T^WՏ��@"��r`g&���qr�SCpj��N�yoq��[A�f���~�FC輿X>RZ_Ǭ�fS��H�o��޼\�3��݅9�b�wnn'�Xhy	�7Z-:�_!PŻ.Z������g"8��lke�`�IX<aǨ�tZ:E���~��	����L�R��1i�(��ڿ��S�5�t�)��<ڧI���r����(d]�A/���W�p�J�?��/j���U��w0��p�/'�;�s����DM�¯��͇i�(^��g� ㊍
6�5`��r��q��dB�B�8���]r�H��
�ҝh=D��ۜR(@K�</I-D'�o���e�l5�������M.j����렡����R�5��4��i�/-���>���<k񓊗�&�9$(�d��,$si��	m>�hLL��x�
�шK�ȅ/e5���pAr��3$��9Ԟ��.t���ݖ`�5#��������[7>�� ���/=�JvzM���.N�<&=p	�ٰ���\w/�'�v.�܅G1P<MY;2�9�Iˊ��𢕪`mt���D��Dú4C�Y�e����{禬�t����ՊH��3���*n|��IZզi}���-���|c�������xj�PKM�C3��HU��^B�q��|g:�N�X/0�1��2��/�jr�4E���(7I�2IVS,�ͧw�8ȵ�����{civ���c�������Hal=9gf����{�#x>�qi� ^O��M�ٰ���/���Kϙ�ā�$Dy����f���Qcv![�II�?�J=M
"�P�R1g���u�樍���s��o��H���?�ds�$�.��' ����wMc��.�#�q��n?Lk��֯�r�I0�1��âl�Y�c�ș]Ҳ�/�����t&|�LC�3�`Y{;((&�����w�-8�[��'��S�/0�#9�GZ��%^G�F�@�!���9����D�@\fm���\]5�m
^��b�I2�ѽ�z恬hJd���/����	�2t���q{{��=��+G�EV�_:���ǃ�>�K$9����`�w��{�O���,�% ��R�s��B뿛��2��S�WpK��YO�Yv��U���I���)aS����fj<�������F���p{ۅ`%(��ǃ��*?!�j/b)t�Igj�*�?��Z,�:�^K� ۅm)�;l�w:��ˆX�t�Y���m
»��nx辩n63��U^ky��t�n����=����#���HpD3:��&Gz��'ei��Ҷ^��s��̽i�1���El��X�$��c�
��Qnv+����H�RUv0�6�*o������ɿ�w{���� �C�k�B�;��]VP�z�I���?V�s�r�Ҁ%�)ptd[��E��6} ~Ef�̹��E��ҝ�)	�m>]��-!W�*�1��9:���꼮
k�0� ̒��@d�h��@R��VX-pl#��#F��YJ���1A��$�Τ0��e2�3���H���Ե �+$�ϦM*�wgW��K�����W�A�Q�-���ً�Du�\�V*6�X��c �'.�܄i�.V�s��`�
h,�NL=W��,�r�s�E�;�:4�E��L����O�A�g,o��,�p�~����ܪzU,�P��.ĻH����){�L��_j�t�*�:���H�LMᓽ�)ۙfz���p�qt'�� �"h9v�7|���WY���E����We�+��ͪY�xU�����]���Ҋ�q���WN����q�DJ�ď!3��� ��O?R�"m�Mf��xvF�7�Gf�_z�s���j*�5�,*�H��mgzl��֐���b�j4��I���r��x�k��`��*n�8/�&�15�x�,J����:&�3��;��y�)P�U�r��!��� (��(�o�Г����ā�B7fM�#��n6�_,��}ﶬ�Ok�cb���`"�4m0�t��
a?��^PdD�O0��ٚ$���ĭ�kT����`P����1d�0](s�X��p͏�F��|j�*]����3}*�<�J+L��무��6Ʊ:s�"ֵyT	��@���[�}[�:*�%?��Nj����hAN�x!�_czo�o���蔬��P
'g���n0Di3^�ufYUa ۧ ���0>� �Z�*��3`��iN<��>�J�9y��ŀ�ȿ�)����.�Y(ok����K4�Q2�`��%��(X�x�����akx|r���j�͐ Pߖֵ�giCʡ��U�.��B����|�N�d�� ��dЖU��!��������H�Ɖ�u�b��g���.�ɥ��:��1�M�
UOE�˄j�K_����^"�</��C
=!<"���=�ܙ��[�R��1�-\�m�nU{_+�r����� -����������LSu�tΤ쪙��7�(��5�1q�{'}���ד��3B��SU��E�P���J���,.��ؒ�׳�I�
�CK��5��y�- �T[q]�?�ɡ�Ax�y
=�[Oa���:y��&o��D!�y�*�3�+�o?4� :��P����O��#`��@k>A�֙���p�Èt{��7�Q�dJޖ<'��22�rسL�t����"7#[�*�n�OS���F��Һl�Pf��'|) �NKc�ڲ�`��f'��r����Ұ�u�^ꇤ���m�1�@�&�����zAt��]���V��Sǖ6�۳r��p�(�n)Aŵچ`~��Tƶ���S����\�R8�:G�w���k�c����R��$��nE�]�cO�A'ko��@�u`c�4m['�{���Ρ8Y�	��G��v�_��"�8c�x��qJ��{��Sq�#�txR�GYF�YM�NC	�+����Y{$�/�7(�~fDx@Qǹ�� ��i�g��%m�M�����D �?�6�G�'V�_C��.�q�'�#�҇f4��Ci2��+V�����j��b�;�3����K�� ��T�<���0˝�aH��@��º��G�-�
~��+�(v{j��b*#kG �&y��·?���Ţd�8-��������B)&�v���y�9ǯi�>{%�/�-�D�%��:=�E3C���`�d�%����E"Q����9c#P5�t���k�d�j�R�j�Q6:�Q(��fz&g�+FwoG�k+v�SG��Є�/����ҙߵ��R:��ά�,F�������<~�H�.�A�8����!78�LM��x���
�@�O�?]2��M*���U��W��,���Q���A�>)�HU OG���_��������`�9Q� ��N/V���,��O��)� ��]j���P�'Et�9�������o�cFP�  "n�S��NI���uc\��R�%�ޫ��"��G^t�Z���+Vq�_9@'�A0K�YuT�哥.�wP�H��/�ճꨧ��jN����- D��A�ѣH�y��vT�Tz'dy��k��V���?A��H���h�� �eK
3���-�=���70K4Ж5GIg-;�^��f���+�E���I�C�L�j��<ߛsy�4=�S1 kLM6 ��<G�k_�|5�O��ܼ��<��~����"!��AK���	eu��nf��Hϝ}W]FT(AQɩ���V�5�l?�'���k�E�5.�1نo�2���&�����c�Q���>�5�I~6-_3�W��61��싰��J��%YUh�|ȋG�+Jۉw�]O�^KF�T[~V(���АH�:��"5<~��lJ�$��[[p��RV���C3I�#���zñ��x���N�i\�]W1��
��;]�p�|�6�`)э�fx Ĕ+r�v�s�(����q)����/bC���{0A��7���M���3�O���U�����Yg�Z_��h��,�v����5���&Y�Ҽ����)]�Ai��y�����}zϱ���|�%W��c�yw���rnN��bM0]�E��L5�V�%DW8�F�9��<%+�t�T㱂�\y���9�L�yπ\�vFt�	Y^��Za�L6
Ƚ!]��a)K��ޢ�ȳ�wtE���u�wܞ(`�H����_�\�Z�5O���;�Y�]�2lb��lW��T�\�
�e�L"X[R���U��>��6Qk=�U-����X�^�t���.|����d�����l#�L�\P$=Q\�Z���3R�"H�e/HXӪW��N��mn~婉]tvl �P��ÿ�k>Ȫ����Ǜkv	֐kOB;�a!B�v�l�;~#.òL��C�{iZ���S�WUe�W2�f�9*�E�볪߬$^�3~���Qȏ"�y�e�!Ӭ���-P���gui��]��Gk���z�U@��A�jF��h�։4Id��`�8֋:
⳾����n�hd����s�&��7��-���~sL& ���>x~�ڕ���F�5���Y�~�j8ܥFW�{���P�²�Q=�EWGue	&��(�V��ءiG[���@��W�Vs��Q0�d���ٵ��[�m��]����� ���>�) r ��A\�� c������<�O��|
����2)B�Y;M'���m�5	P�^�ّ�Uk��J���k������YuP!����;�65�ﳡ��#
��_˙�Q��w�SR���v�9��,�#A�Cg7ȭ_J_l�k�?��(�ҥ.&A�%]�\!\���,z��YEa�	7&�Gܔ[�d��d���K��p x��[�A3f�]�m���>G�,�2�M05���O�t�И�:�� ؂O���OHe�A���Xܙ��9S>`Ư���'�J��t�Hסa��=ό�[T��%6�5.�����R��d_��\���x��A����u�w�Y�2�.�_8���f���f\�j6L, N�2`���h��4�l5��� �q�l�Le��H-*��],�3_Q ��j�t��@0�W���q����p��)8LO�ZfoU C2�e���On�>2"^�Xj=W��tj���g��UE���:�p��8l�A!@��(���a�TaW�;�*���80��[��`��l)p��w�'��Ǧ��x�!v�[�%��%L��HHyX��q'Ț�N�hG���=X�קb�����Ե���� �=�V���>ؽӁ-v�Y4J{|��"jY�S�"}M>�G1W�wng�"	�7���6����ln��~rς�J:Z�n}���rIUJ�k��W��[�W6=�y�'�wqЦA���&��6�[g��/%���E���p�XN5r,V
e�x�'+F�s`�	=��L ���#h����x c�PL��P�az�=	���A��T�2�>��^�����L�{6a��>���-�Y��k�/�������&�o[]����G�{��6�J�s�wx����A&/p�+D�5ǅ��X0�"%%6Pbk�3�������	J\P��i�k��$����%��ޛ���>lR��Z�49�WQ�����lVy44Ѣ�]��z�3S�X�#����n{������ƥh�VNk*C�dV�HK|���CJ�N1�?�п�؇�R����/�	D3G�	����ph`s5��������AB�f��&�6�d���Ǩ?u��B�v���̥ݐ��kʓa確�D��5���q5)|/`�d��p�(�:�[d�g
�����&̞��xƤ���*U��>�=��V~;���,d}�/W��<w/ 0 k!qt+y��}�p#su�m�j�]�Î͞.�u�[�*W-�RB(��;�����{�@���8>PQ4]�5m����.�?���X�N�k^�]r���y5Bf_����{]�_$�Y��]��͚������FK�ʝ��W�%��weҷ���x�$�\t ��:j5���hR
�ݬ�^+-Hz��� �H�H�DGM��%�v*��1KǁZ�:!LMIf:iW ���R�m��	XU֓|D%8f��ᨐ+��\y*#4 d]�~/��h���Ju�˔_e!B��i�#��%�W�̽9u����f��s�)�~�Q�XP���Z����#��Ɓց�R��yg��0?�; h�C����>�7 ޖ֠�A=�E�]Zs<#uw�
��P��X��1������������(�BP$�6$(A�5�痳z�����h�!�'���1��L8�2 �Iǡ���rW:�I�˦����R���Oգ#ӳBk�(�.����x�9�Ա��ţ-R�IvgQ�������/��t]��	h�g+��t� \cbtwsÐ<�?s�9}�S�qK�Ub��+Ќ��ps� ���lq�|4�!>#�F��sXv}�	:���G��& �&U�Ck��wV8��Fkn�ӋE/�o���P�Z'��z�(�/�"�����ׯ7`��[��Fv��W,!����&��=e{`�F]3�ӧe2πE���ܚ��S��M�t	�.���<�6�nDm�r2���f�Y��ϯv5Q��wF룗�� ��痍?��M�\6��q���X�
Ld�_b^y[�{��*�ruG�w�����<�/7��qt�^�+�)�6ҬJ�O���.�f<aeR����MԛF��?�/�x�f�}J��o��&|�����T�b�=��_S�6��N\
��}��Ž���g
�R�+6�_oy�~�!5�7�=��o�_U��m�e�{�,���n;w����0$���;���lD.O
~��.�z��_r�����4wÍ�<z��BF���_0�Z�L�5{ѻ�t�ì~��P�0V��_Ju���B4 ���X�*Jm���v����|�LP�
��0��l� p�g8����LQ��A4�ڶ�k^/�I���8�WՈ���>�p(,��^R9#�P���,������%�}����6��$�hoL ¸�܉���;C���%!�!�t_r�����}�mo�v0�>��D^�Z����r=zL'�*H�f�: ��\HLSF�@����"���ϧt($�.���4u�����9wF��WS���nMn����ܣ8��$-[�y�:�k��OY;�xM-.y����.�S���Ȇ��L�%a�3ۡ���i�m�@̊��,�dƝ��z����蕵V��#���&+	M��VL鿑��R�g�Ꞩ�h��g1�&�B��+l?_�g D*Ns��*L�&�r@E����4I���-������.{/1M����"�G�DHZ���AI:�g�}l��*q�
���b)t�����,a;��?������Z,�uMX��ǽE|�#��yG������,Ā���XЀ1I<�8���C�^#��*�)�[a��'$��r dVC��0"򰴟g�4�䶆[pɞ,�A�;|���ub$�_�܉>sXAt��hS�����,�a����_�/z�߉�)9śy:�B����B�E��d#ں�h-CX�ӹ�`X�T��H8L�����Bӗ`�?x�a4��G���$������A���e�#yz�S�I�S6L�X7��v�jYb��Pup
��<�yk��ޙK�itpt�h1�xtS�C�U��,���;�m��Vy܅Wu��0c����	������H�S8�&���"NC�',����~���j|��QFa;-c���z	��җe/��_AYanp����P��fq���)6�z����y�ިv��������K%�G���ג�Bb0I���.*c
s�X;����޻��!X`�G��=�ʁ�Ɔ+
��8���_�J�_��,�(=����א; �|J"�n��L3ԪIa�g��R�3"6����T���:e�j�Ŵ*�4�*�&�N�Eg��C>C�S�q<��B��c��l��^������LӇj�4p��F@�g P3-G�E��d��� �Ҏ��We,�]���SճY��:D �;kh�"����@b" �b%eϕ���7�`V}��,����d��+�DI����	�<~��_/\)�:j/o�x�RH���m��b�[�kW��ϟ����r����UK�h,��~L3�F��U#.k�u�"��#vi#���a�o)��*D���#�<Q����Sq��Ux9|�-k�����Z:vK�b��`VO��W@a��(��������<��&���l��\�Qd�hX��w��	�IX���1ȃ���T��#�+���N��\�f��r֤��ʒU�Z��ކ����M�w���и�oZ�;ntS����Z�՟	�nr�0r�=���4��lU���:�	ba3�*>חSE��	�o&���3G����Tx�`=O�_%)H���ſ��:_�ю���F/�>�tk�m�vEE���<=�P� @>K�-���
��	� �4D���E#Ao�P
���Z`IXȖHm��fk`y`��K�ⓗ��S�^}a=�}/���~�v}qu����I��̃������)���j���E���Y�U}2��U��q�|�t0ր�����~ͧn=hV�;�M����S�
V�r攛w�^(r���G�(�}V)�_�V87�M�=�L���7f�2���HѻCQ���b�Ѱ���T�+��w��^
�ӭ�)Z�pi��n%HG��D B�CG<�\��դf��}���Q|�ͽW���f-h������3qL���=���I�N�������B���s��eOs�b��@tB{����dW(�4��K4�n�S]1�$��PD�6`�t7F�0�~V��*��§,�^�~�_�+W�![��2VC����1�.ٱ��>o�xɠ=� ���"�����^eX\d?���f<W*����m5��w�;e��3qt��|=T����@[d�w<+�D�KoT�� 7��R�˹�Aj�������Tx@���7���v�M��5�m�-�vau��A�,�gt{	ޡ~�}����cf������:�>�&����f����~`�Kje�IZ-�����?j2����W|$�ө>`:�l�Ix3J�"X<GR���WzmW�{�<�-l�V��o "ĢO��&Ë��`<|ٮ�5x��Dj��V��ST���[�j��\țw�
�$�D�kk1�Ak��ᐿ��N��ֈ��I�'��KK�(�@��3��cܷ�]w������g���T	�#�<jZc:y5*�i����A���y��&�u�0F��όe*��&��H�^�d�s�J�z����T�&9�	Wq6��P��A�?�I2R!��n��"0/[z���X}O¹|y͈��pS������+��q�2�u�u����xX���e��8�׳�0h��Y�%I���?-��:���g;uy��L�&[���|�/ ]�j�w{�L4e���{�U$I�JD#��<o�-Z����(�t1�l}Q{�<X����r�Ǌ��K���y�4%cQ*p��x4z �����w���)����F���+��V9x�2��,_fԕ}Qq�ܵ�M����1��� 	?D�!��f��vN�U��X�	��~c�ɜw�i�g�S��M�#̷�z�w�Q�#�����H,4��&R�4ή>-�9���QF=Y	������P��H!Li��}��S��}��pZ#Y�y�;gfK?>������I��V�\��C/��n��p���0Iz�5�7R�R�*E�KtX
�:�2d	�C�
	��Q͘*թ����S�T�?s5����81�!�g���H��Su���n�ݿr�+�q���債q!�ڶ�
��46੅>'�h��5�$��k�����qc�	���ɨi�
�/*e���m*l�[bR�N�=e�{�6~�U���Ԯ��	�����0x���d�!�(�J�(��k4�ܤ�r
��������g
�y�5��C�>#�Fg��>�&�w��ΎM���|	���e�d�PX����$������G(���S��n Kpzo���{^\gv}�k���"����t �ӯ���P��"tg��4iڪ/KZԫF����Dֵ�u�,�%����/hr�8���l� abE�#�&���î�Xs�`T�� dE-Hgw3��1�#�V*��_���6��m�`��k���W����� d����i��b�N&a�
�T�4�a�"@(a��ӟv�w"Y!��/�� NJkw�3�ʇ��
��+�냺*=�jAm_��������E_O���XT���d����cY��B����"(c���	mH3�Tӫ����T�j�lڈ�acͻt�����A��	�
��۔I�x�#��4L�	��i��4�I'$mK����r�Ҍޥ��/OD���H;�ӏ�c?�p�fs�z�ט�$P �_יdh�r��^<M��7E��Rv���9��F���׵6��d����pj�{ޚ˭�f'��1�K�S:�VF�5��z������f=C�wC7�|d��E[,��q��'�u��đ�E�`-����%z�6����e�?�H�Py�<Ί�1��c����x�4~�q��ؔ���e���?�E�L�mvF��c^�ӛ>�s�)���>9���u�3\��I�����~k�w�n�Am����� �٫ݫ�S��̊����dy�ҭ�x�����S�%Uˉ(����l����m���{Z��9A���I��؇Pq�c+�w#>�A�fe���M�q���6�UDXr
Ǫ�T��S.t�N*}�<7�~��;��O�:�K`^�� h-"b��4����Buښ#g���]5u �.��#Q�_a�=+.� ��	ZN}ˣ�T�i�F�8u��=��3�3-G��R�#������$d��_JOF�7������I�F���ξ^G��p!��,ܷ�v��<�`���Z����۶y��m�Q�����Azs8��9�n�e�m���K=��/dݬFF��w(��2����4�<1ܥ]	-u�O�8nL��^%���i��ɱ��#�£[͍F$Jp@����vʉ����v�)e��(A���Exj}�iUS�AC+�H��[�NE���+=y��RRY|쵽̃�+�ɲ�y�Y����`$B&�|��IbĽ�B�V8�p!h���6�8�Q͔�x�H���W%���R0g��B�-F���h
jꠍ$ϛ��{�w^c]rҲ�� �qq��+OX�3D��F�j�u^����n�:9��*�����>�jHf�6��b�^լ%1�PO3����Sw�b=�� �ۢ�e	���a����zw�g��9�y���?���gs[,�8��Q���S*�ؤ�Z�G���yuZ�j~�"�����q�8Rf�$�\��]�����b}d��k����1ƈW9�1܃��Xv8 ��<M9����`�gU���X{������
M�m��(Z"p��yCG�.��ZE��a�U�8䱢���2����m�����.��p;�!��-4u�6,[���;򏒴b	u����n��QF�����iH
ن�-
�Ӫ���["<XC�KD�X�
���Op!1Bf���W��:b�N����p@ݹ�_f=9rR3:Y���e�d��Ս$��'1�)��6{���jphM{�:eLE̤ή9�1��L�LJ�i��4%���9�+��2�[nh��8�-2店\��&9�KS��� do�������WBp04}�5կ΄X�@�e`ہ��6!Q��x!~����4;�dP�苁k��ի���Sb�#nc�TdIsl����ҘmKl#�MH�r��~�bS'�Q�(�t�f�L5�J2KO�,�B�lr�@p��0�1�N�8U-�� w
�l�=`;��Vͳ+�C�>��y,� ��.�xy��ϔ%��菲�6������:xQ)Ռ�ȼ��8nQI��k�kb�%����6��p;�ٿ# D���5��{f�:h{�u���Df�/� �G�ٷ�����At��<�٦��Sg,A���K��W����j�j�\R�R���42=z���S;[�6eݛN��!UpL������G� ���b"�m�u�(��G�X��i ��y��0:�8��d����Zۊ����y��R��۸ �������ãl���;P�ؓ����{���E��Ļ��Zz�*�%B�(F[%/���)jD���Z+8M6�w��O�"� �FM'��PS�[�ڳ�[��d�Xd��a �g�#��a�<�������4LE�/h��h��r�Aw���`�WB1V�R?��-�i~��U�Z�����zN�9�&�+ީ�(��Y�4��`��Q�����F�����6�\�YD�%0�8m b�m���2^�RyU�bm���i�� Zh=�%z3�?��9��	�ŷ���Ѩހ�@-���Y���sQ���-ɹ���E�5��[VS�^p�+���6|w�}D��~ ��~�@:(۾����#�g�@維ad5<��hN5/��p ��W�ґR,=����j�HK����4���Z
G�gK��g!��'�_�R\L� X|Evs�D�9&K�sf�g�&u��ց����D�'μ
v��n����"8SL��Y��������0G��L#3l"��ɛtd+*X���";�Wy#�^z���Д�~o(�#�����^'�e�Ry�@@�?.*5��oK{�W�D�'�kk:&�����䂃���R�V�9-��$����CO�ʾo��K�$�aZ����G�q� ��T�c{+���mS1�7'�0&���=�2�@���JPJ�_7O��W�_D�$�%�0����:@���mk�^D�?$*�g6�y+r
����6�n�@cC���t6���� <Ye�q4�81J�U�pI��6�ݛ��C�W�Of���ho�{=�"�ܩ.
�-I^4�诿����;���yXb��tf��sM$���Ē�u2X��%���ʌ�E�FxW�QE�D�(�'2H�E{�� �A!����=T\�}|j.jRm�M�Z�?�Wc8��)$�X�B�4�Tv�]B��i��3o�ws-��vcZ��8G��'>���s5�e%+DdD`y�%���r�L{��s�T~)����Sq��9�ߕw�gֻ�H�N��&��Qj�6��$�v��BL4d�%k�������<� ;�����.��A��XpzCK���2�p��5^��!Ý�{�B��=��Jw,U��8�ǐ����7��}c�g�Z�O�Ђw���6r�|^��\}���b�p.��u�����I�5�ѩ7ѻ�3�Y�O^��{VL��=whb�k0�am`@V�L���ek�b����ALU|�M3�v���]^�Xw�n��\G�3}�AOﯸ��.'����,Z6�����C��;f�d�uǭ~2E��Ӑ��6�FQ��R�8%%0�^.�n�l���^`��e��a?z��&���O#.	$�Y���F�:�y�av��9�[��֮�qE������1��@�L�Cr��T�Ss��������˜RfZY��j"jL]����5�<�\|�C�m��dк������g&��ahb���u�(9��KQ'��Y
�S[�W�87o�
��'���,��Gk��ͳM)�OU�$����
A���x���K(g���)?p~�,]k6�>��Ҽ��#��@�����Ws0��MZBPU�,��2��D싇�iu�q�baފ鹦�	�R!�j�duF</�r�8�ލ���:`߅=�u�΍q�R=5�>��|G��d�t�3�Cp���+=� xpɹ��pk�n���x3�>_Cy�G|��]�/T�徏�s��EJr�;T����{�k��9��N�4V��}<�!m�Q�f�ܭ7�Ƹ��4��z4�q{W/�]m(>d�Z���\m��bc�-;4�=��br�t�-oTdy��V���x6�������95�뽨�
+̓d�o`��,Y�Nޜ�	�m�*��k�==j.�2�6A��{�Q���Ŏ��F�W#�l�8ڄZ����<r�Al��l;͠"��_~m�7k5�,*����!�ox󫓯c/j��T�a3/9�,\W�S�L�ޤt�r�p�}�D��1�M⽜~_	/��*�����ߗ}h��k昀��"vggq�iA�ij&��Y�Ga0w�?~(.E��۾�38�U����p�D2	��g�VSc��{��
51��D���)�M�����x���:�̷�s�'*�*��ڲ`Zx5;%S;�JC�JxȢ;��tʱ\ݠ�%�|���P:	3'՟����p�J菈��w�s�'��cn�FR�X�Ev���VU���9�Z��8\����;�
sߙ`�t���U�Q��މ4P���+�C>K��$GM	�d��)US�x���D��́�b�C�4{^4�	���O~t?gF>/%��W7,g���/�Sz��g+�na�`���Nu�:���9�)�
�'R�,��[�rZz�����:��9�
��p�x��ÿY��_�SN����O���^���2���K�5���?�
<�7i@p��OǷ���gX��p?�֙���� ?q�`�:y �g����606vܬ�0C���/�������M#�F���y9�9	Lh��ߟ+Vڐ_w�p�
���>!�}�:�6�s��"��e>�4����]�ǽ�����Uae,.^�\�����N��f��In��NK@6ӕU3�o���dO�fu���u)�R<�	�a+�2Xa��_���jL�}ٲ�K��"ݗq��=�����㿣���^�2�b�H�!$�!Lr!�=��3�� F).�_<ZC�_�C(/�j��í���޲����مS�	?LS� wL�8+�=��������gdy+l��-
^��( (�t��������������I3�V�'�ZiY5�`ڢ�h���,Gw�W����g;�~,���6Z�ٻ.E�ր�V{��f4����B۫�ט��<s�;8��B���2qꐛvOR���l���N���|3�����L�B�%��"�����.-�V�1��E�F�9W�*^��`p_�D�A|��׾�b�D�ʍ&�iAȚ¯%�g@��7�Z�%�����m|๥i�1�\)���7g ��k�n:#K�vr6l	~��,Ϲ`�|3�W�YI^0߁
�h�3"x6���9a�߿�;*��z_\�Q����k��nL��ЩY�:Q�&���!��k��\�5����I�Ȓr�f��;�n��������
��̟�lʛ���fk�B
^��#"g�DB����Ieu,�2Hly��܈��+ ��Iqn�}4-5�����8oiO��/�k���NN�V�W����2	ƨ;��N�e͞e�"�&�y�S]�j��K(�������KD�-��~�H�Ï`ҧP�p��FZ�`��A���u#����� ,h�N�v�8Ox�6'��)��-�,̰)p�݃�bC���ڤ�TY�Ib��Q�ۀf����Oew��� C�w$���F�<*���^!�G���KX�4�8���O��V�9��l�!tpY�K�[��;���fÎ ՜�����)�p��I\���t<���أ"a�#��Ի���yNi+dI@��5>gn�0>��*-5���=Q����(��3���;���4������"S��ڲޥ�P��U��|�x�d8�ȝ��'9ĵ	�e�i�:w�'M�W`3`�8Q���R��I~��[T�8f�j�5�ŵV,��O���ϟҚ\����G�R��,8���ܹ�;�<P����S!��hK�~ߏT(��U�p�,��v\p\�f���a�����kCa��UxvtR�|"�LK|ݙ:.I\hgzQk�e(�"�?ZPa�|L�������������'�hr�/Hr�.�r�:X�)��o�FZ�H��azc�Y< P��q>�˱8�������YŌ�,ePټ�����v�d(H�x�Lj�&j�F�riה$�0�;�v���u�{�6݇څB��si{Irz�{3���������O~�Oh�@!sr�w�P�w���w��#�߻��w�DI�<c��v��Q���㠉5&C���t�nգ:�_s���D���25�GCV�U��}y��C "����y!X�ä���g��ࢹC�����{��Z3>��(�dL-�@�����3b���r�a�ߩQC�����4�m�1��^��x&���+��y
Vl[ג�j(�I9_��B�����%Q46��?XA�~�D3����΁��	��"����]�%���A"`S��2!V���G�v>{�a�8{�I����`���uڕ���'�ʞ#GȩAc(�K�)amY��X��	ҚL�`�c�X9�h��� �F�+�ƈ)�V �{U��0���t\t�:�(��R�9�w)�����z�6�;�cƿ�$o��Լ�w�8�'�C��ǖ�^��T��ܖ2�υ�p�¿�U������C!�Vpc������4�$�*�9�tK9ˬp���D`�А�����턧5��C�3�Y��OQQ� ���<��(�6Z�>��7g8283�6M̉_�tK�V6?����*�M'�o@޽9[9�~1�so���5�y�ޟ�*��_y�F/*WX�)-�-*1�G"�zq��}p�Y�	�L�#�>r��(�M敒�+�4�xӍ��G��D�l�ѽ�|[i��tN�vG,e����E\s#3�=�b7��f ���4�d���h0��#�4F{|�h�y6'��H*�� �������/��zUM?	��du����N^�.H�2�=�z)�`��0U�h`@�-��z�J�Α�Jʋ����U��c�.r*TEi`(wͤpݑ�pM�Ym(5U3匧��!F��nQ���	��؆��o���y��l��^(��@�����mA��Ϻc����E>����{�^E&Ɖ�:���w���FG�H��
��W����X"����u7ڔe����d��z��:ac:�J��m���Q���w�{Cj�{�N��v�G������wt�mԧ��[HY_��}�����-���k�G3oQ\+2��q������Na���t)��& @����E��uFN����������rB����u��|���W����z������|��^$+��w�m{ѷnIj�A#����~8i2������zÓ.��-���5��Z�9�T_����oB&��#�[{���߈s��9�&�(���w�����ҕS��=0��z	������l~��@�6���FM�����]�l�j4��׾U[����a.=K�`*��$D?��1Y�NK���_A���|���TVM8�D�����&��G^��&P[�1�%d�P�K���7 ��|�`���ؼ[(,�^˷>�����G_�d}�e�p���q:�W��<Unf��g@���w��6�C~�f67�.�
�g��wC�?2���L65�]. �v�'B���y����cͼ����M��U��R/��5Vղ�]¨���O�k_�+	��b?��Ó��������s?L�V�#���5������c��˖9���R��ڒ�6Jdo'w��e����
AW��O��yτ��ݼ��L��H�gF���z�.&m߯��^V��ۄ�I++3�'(J�WT)|��5��3�xBeq�\��n�>�i)���zZ�O��T]�C���!r����E��I�'�v:�	^n�Af_���m��ՆHx���D�c�Vޢ�d7+'�Ċ�?a��F�AQ�)��ћx�8ZM�QG�V-!�d�5��4I)���[߉?��"�(����ݖA'��!k��8��Mu��,x!�ǤK�~���:�����-�W����M���e�5���Jo�$�C_l�8!�d��;)*x�>u��'��Kf��\��ґ?�e����k��4q��X����99�ME+��?����.�؀��1����z�	X��fs~t��Qj��$~�,���.�ϥ��xף{u�9]~d�����K�]���`�g5�1�/��n��Md<J<i�ophU����S:���n����n/�+�D
�eM����롸9|��7�_r��#���L��H�RG���D���<�ydG�A�G�Q";�bc
[`�u,�uT?żf���M����6��m O�ph1��CǨqE�{h�0{)�:vw�/��$�ѻ�Jx��8gQ/B0
��.��lh�Q(T�S�&��B݈��oD�zvRj�Nl�Z��s�fJ�o���v��7SE���O>E���2�i+B�4��SlB(8`�Z�s�֚!�j��_�n��B|��H$�)c��Z�Y� �p�ۇ8���]�U�n��S��!�2��-,B*��h��)�ܙ�-��9�\>C�ۅ�?�����!ә3�TBS�E�P�g`PE��񗍋���&�{�O6Mw��x�F�
�j��`��Ɂâ�pt\�싃��]�'�ỿ���朸�U,{����<�*� ����R���w�C�DvhF����u�uP�I3Bm>�CF����q�z.�EҶ�S{�wβ�q�U�͘ 2^�ҕ�������M�	Pڡ(�x��������Cp�^l����瑇G���i�vp5�K�4A��F52��>P�_2p�����^���V�����^��ZsH��T�z����k�����+0D"���C�y��(��<�>�N��J T@�U�}����1��`��O�H������N\`x���ډ�XaN�#�Xc	���<�3M�ۍ�+D�x��DSFL�tCr>�T<�́^=˛��
q>�u����[O_���i���*AYL?��_\4� �oɁ�0��_�ui����K*^��������"F����+�`W��-=� R�v�/ӽ<m�������|8\pa��+/���\��0���(�$���w��cR�,A�:N�c:
@�r٩��)�x���S����<ke�!�wV���D�:H�3��|U�)��pu9�HT?0j�@qL"�]�y螑j�*c��nH!�ϊǦ'�]MW�Z�)��\���>�1|�p��ԫ1�{yڐ rZ@�^��t�_h];}:��<J%*�a`�9;"=���Z�4�:���P��Xe����ƈJ�m��N�Zn<WX�����V9�ʰW3��б�� u~�`�S�o��*
�tB�`�ȤQ�����>L�B"��w��I�1�
	=f����%�#�ۻ˂�b9W�H1�}���?ӌ�-�};T@o���~�C�8�1��ܕ�z���_}H�G�Y}Z�YEҭ�a�\	���ξ��JZg�ن�J���u��m�����p��B�m�j�B�#���0�+�+aɫ�
���	�'��i�f�1��q���_��E'����k��v
k0��r��h��*�����C�%�%�����������,���U0#ٳ�T'�줔�0u"���v#Zyqku/�I��՝���l��ykbz�Q䞮}J�p��X<���i�/8Fj�93�PO�/ȭ�̫��$&���2�����$��FeT�p[P$WL��S"Mx�`T;B���r{�B�2ԫ��l���o�2b�x�A �`N��J�ݢb��(�|�����Y1�$��Z�s)d%�g9>|7 �ކ��8ދ/�5�ii$f���7GPc�*��u�Z�������%�	���WFd��U�H�\:5,�+t�{�lv�����L[+�U�^Y�
�c��R��YLQ��f|�ȻJ���MRȗ���B���	?Ql�r� �3B��%��r�ZH']���Ae|�P'�;jjOǜ�E3�����/��A׀�G
�8F� 2��M��֨
�,�D���g�؏#��u�Y�U9&�i.n�A�!���'�:(k%�[^+��-�(�̝�#�~�_�\)el�����^_�T�
��+A�m������ި������T�p0b��b�pl�܆�:K�WA�`��j��cCA|LR�O��s��s��oMZ-�ݵj��FF-�)[�\�Z�@��_6����䲇�8h{�[�*�m%����&��<�9}���m���%�
���W�%��> ���.�!��P���ks�K`}sM&ra���R����ص�Hq�Ą�gȅ����x.���3pY�ϐ�lm��7γ%��=���ulA�QJ���k��|Oǆ��2����9t=�f����jb~h����W�޶���$�+�]��
��BgJ����j�&z��������t���W3<�����o)nV�M��SE�h�Q9�ݔ��jyj�	�-k���T��r*u>gW��s��m:y�{<ʹ�⪃�}���S���mF��Ԏ�,�f#;9�@�r���}��i��V��'�M��P�w�u��QBx�=�&�I��1[�aȶ?��5����#)����};�)��r87�X/�8\�:�|��F�Ǘ���Fl�ȢV��T��զ@��z6T���Ҫ�������O�$LmeQ���ۜ�Y�������VZnB9��j�w�R0	V�O��tR�4��.؆Ȉ.Gj���ck���F�qPA�.�����X,6,F��Z�r$~�Ŕ���Gyy&�Y����d� &���!�S����a�L֠*umLaT�:%�(�R E���z�t��C�6w�˞��W�E=Es%ض!y�L�(h)�߯�T�I{�0��Dx����i�+J}l��o�a
+���b��)]�|z�$)%_E����i%O��M��M��㡪��<E���,�i�P��A�XqƬ��� ��:�����X�� a]���������wO�k�]�.��h<���$ ! �.�b/�� XO­:��]|��(��ޚ=�c��r�I���f�Ԗ2F�3���	{�y}��Ʋ&���i1G�M���IeI��TnQ�a�0`�R�Qt�I�w��X�\� ��V�F�T<��h`N.5$$5�^�ؓ\Z8ŗ&	8�j�#�W|�!����to�R�+N�`�L�O\K�jp��ΙFDu�F#ǘ0<"�ꦬ!K(C�0	�ۄ����B�Z=����I��ˡGVZ�����ڼ�$�3~��gj�[w����L�uB�d�뒺NEksdyͶB�Ov�}g������C:���&�oh�B��BV���i]q݌]�� �U��;}{J��R�Y^6��Ǜ��tu��XrL�0	D�v��2L�J�ZD�V.Pk�b�&0O��vZ7��lr��Y��ֈ	%+����`G���&���ꁪ���Q�7R�F^b��7��&�ڶ����n�܅6��_�w�v�BmW1�`8r ����Fm���;���,���0³�\�v5�z��0��u2���P����c�k�;iH~�_���Hۏo��a���[k�2��
����]��궚����HG���eZic�N%Zp����~A�32�&�u�7�QBl?Z���q�"{Z������1��<�8����������ԓǱ������X��Bad�V�ɥ0ߦsf���L=ʉvb�����M����}'z��K�=N��z�E����q)�jmi�-���X.5�*��' {:`����nB�1~�P����&�O�KdԖ��,��0F�5�
O���8�A�c0*H�~OUS��	՚τQK�$`w�i���s�(=���,��vB#�I�xQĽD�}�}��Q�y�I�`[o�^���c^rS�O:�{������`�V���w�C��$rH���X�t�uI/�«�ē:�,�G��5����}��v�Ϝ�9�#Q�Z�W����応n���߻�d��0F5���A�h��\,�)?A���<#w�7}�df���t�����{q�0\��pɁ��K�~��x���(�_����ڱ�"�/���J[dM�&<|:��7eQ\��Q�����v�����Su���^ޟ��%P,XR)��}*Z�a�o�_�fk��[Tt�&s����7%���/z`m?����j�5�)ʬ��F_L?}G˟hK����0�zp����9>�*��Mas��쑜�|�|����Ӝ���U�o'��Ζ�<5\��E�(v�11��\�=���|4E�4�Asm��I +f��U����kT ��iX�j(������5���y=Ã�T��ǉ�f�x�5����-�mnϗ<��c;_/�X��D������ݜ\
��[�I�ǡWw�0�V-�,��d��c@�PǼ���	e%�"	����Ts��3�D�wP�T���
�Ǆ^ń�~���kΆwV���*�R{~������\�)�3�2�] ctӍi!�ro����Z�Eju\*��}WK��3��q@ią�+����GQ��T�2�56:r��m�,i��w,|�	����(�5j#g���ܟ��t|q��'č�(X?����E��G����F�lJs�^KU$�f.]�H�6lEBD�碛�	�U�d3��p�#���	��e����M���X���h׫l�jI�Y��+���R���e�1Dǃ���~���kAC���߶:������W)�e����#�X�8mgQ�XY�/~�t�]wa�Ѹ�)i ����i�D�
	���/�����`�Q��v�f�d��ZZa�~���C2��`*���f�����/X�H���z�=/bhʡq��{�]��P��9�����^�f�!��\��������I�8�3�߄|֙mͰ��HXYL������1��:}P�Tjo�X�F�D��M��4X��E��� ���S�9�������m`�VC)]�^� �����B��֞�+�`��k(�I�P�/�i���t��_?�{�����攏�I��~���ǒ֫uQҧ��^P4�z��恁��������\�1
���5�D3�Q�V��a���łLuw["�X��{���������L������:((|�J�}�w$�K�r@�@A9Q����o[�W���W� ��ĵ]ܧ��3������r�'8�yL_�p*d �����Q��.R�bَU��>�8q^}G�**��{k~a�F�a:�����H�9t���wش�J�rZ+[S-xr�VO�{�V���a���L�O�$�F6�F�����YT��~E�t�Y)H�J{�1��,���'��J�{�6�5=z�`����}�=�w��ީ�S)'��dt���~稕Y�o�Rq�jGO�ܶr��?3��^�r��ູ}&��� S\��X��۪��?��P���ț��&�	���q���H�:ؤ�ͫ��
�MM�k�ݞ�K�L��d����`��ำV�F����7ܖ��z0�ɳ%l���B�����|����6[U��`��m�x��>`ˤ^m
�>���S�|࢙�����tC�$Um��.jp!Ο�*���C\�SVJ����g':�C�+V�?WX�0�0��� 7W�[���2�YA�
v��vZN�`��,c�0f�q0`������	iG��{x<�B�	�ӧ�~m>�#�Ǒ�ɕœx'/����iy�59�9���?��#����V<cseB5��a��w�I�F��H��MGA�4gy�lO,�Y�2��<<��6#%.����f����;��7����CRŅ����|>��5k^8����qP<���`���KoH�����Rg��E(=�C��-�4E� �侖j�|a�2��ݦ��տʏ��kĘd��
<�ad}ɓ�cJ8X��*_��\��}n�L~�v֍��~�P�O��B��U�'�0�z*��)�Ql�zĽ�cF���<W����������WS\��)?��+[
�+�T�Q���'�G �(��g��ᖡ[1�\�WY�����>0�wW�7����B)%���#�1&��y� G:��7�P.}h*��U���|��c)�,���]��iU!�#T�ƞb��:m���������ބ�e����k���d9�KG(.�N����\>p�k%�G�O��Ќ���(2]=�b��*��t���hW����+)��P\<s��u�\�%���drܴ.P��^�����1�� �kJ���R�L�r����LJVX�s�H Tfٝ/һ��S9�D�yOT,M3�p��,�e�[��1m�Cq����B�IZ�� ���e���a���|�7@���m���a���6K�G��3{���:b�2�`���C.i��ʾ@�4�C��`=L�|)�[U[�]f���Llþ�P�x�]Ioހ��Ձ�`bC�ֿ�qnx�{��=��0n�@	Eb�`5��h`����#@���x�VA�.��G�~E1��$2f�5KWl���ʏȉu��Ct�p��Gz�u]��k�HB�<-��Q"�[�b�
9S���C��v�KQs�	�gȌ�T���@P.x�!ތ��h��yB&�Etp[�Y���5v'޿����=�p���!7��"HJ�C#�'�C�R�� I��Ne�W@K��V���R'�A\�R�dS6F2͋n�
�S�� �Q)��R`���]���U�{�u������P�TQ�\o,C��_c���-��:Wo�X����t>��$vE'�
���B;�N�}/��Nd�
�F|��`�G����o���C��%�F�ᥝR��K�O���^�Őn�ZOt]�ΘS,n�L�Q�XM	�b� �R^D�x�/��dH�H�o� ���:w̠�I�i=0�:$_�N�Gkr��DijFā]�=�9��u���DA��B`��>@���Ǿf��TU�����_<��RҔ���lDZ�0$6J�ĳ��7�	����e���a����:5�
��j���Q�� �hl�?٥�	p��fÜ`�|U2g/'��Vr��&�?�a<9�C��DPѨ&!�������F#�h,�yq��g�?1��ժ�l|I�tP�4��/1���L������67����bsI�� �7{ၣR���	�1�B����m�[�H��uC���Eg����&5��_o��Dڸm���3�H�>���C�.�>�ae���� ��iO���<��Aܣ5��?�����c����@�	��^Ր��p���ϻ�X�U����`\��=�`��m����c"�k~�\T&ɂ��ώ��� ��b����*��m�$Xk�Dɡk*^_n�b�mJ�2z$-)Π�{ji[��Qih���������8�̽��:���5c�c�= ���B���Hʃ�I�IǜlOHE��b��)���ۦ>��h$١Bo!�K��!�bl*-~{e��ݚ8�屄��tr!��2\Ń��f5E�/�1j�d���02E��Hܵ�^9f0��Ӄ''Z�E9�!�����ԡ�l��/����3>Ggz`����*Q���c�9�݋tl��{%���o��znX��uo�S�v��+�Y)�*�V��bӶ���d �~�X�(S,�y��N��JN�0f������i}7�?c7�iao���n���������1�S�̀� ��^EK�%m�Nl�}�wB�cפʿ˄Q)%6z��B�V;%��=!\�0�'�~��xmG�T�=��Ƨ���u�&�-R� �5c���~O4c����i]{% l59
a{>MaG����2b��.M�`��Y_��؈�nV@�����p���X���qԤ?
�l�&��o�"	�f>*���u�u���NB��8�����L%�}E�N�J�Ҝҝ̞'���ZYn�8k�r���OH���`��RE�$����]�Kp�!�KN�O�\d|�O?S�NE;��#~;a���{_�4Fl./�+�V��О��;�wqHY&��ڂ�A:K��U���|�rf�F��KI��fq�z������x�q�O���=�.d�F^X;A�J���������o��)\�f�m7������_�D���&���<�z�7�����.��Q{��-ʏ<����D͖_��h�B�9�{�6�L�^p���
��}�tq=cy٤�'~���;�XV�Y��ۨ' ̌."�?_v�|$QH�'qt��x	��2������ڰӿ�J��Hf���OD�p��;�˳�*��v�E���2ƈ����Q�ޚ�4��]���:���R�y0����G�D�&֓��L=��6~\�'̹x���˩���0�2���'ό�wð�č�1�YE��0� \E�����a����Z_�>Օ�4Y�6t�����bl����u��4���M4�u�%��Jo�q���{�ES0`�Mn��̔�-p�!�dϔ�,��1m��Ba���+m�ʤƂ�A���uF`�����+�ch�� C�lel���(O���R��\�c޲>mT{����2խҷ΋VS��4�gb^�#���r�O��(�G�-�z�J�m!yb��uX�T�fG�_!��DWP�j��.p%�qsP����1a�k$�U])µ�嚋ܡ�r�Fx��~fFv��q^MK�6|����h$�d�-�-���@��>8)7y�&~�[u�#!� �E��?js��Be�&�B+b6)Me�n
bWNqo�$Ț?Iep�>��Pj{/9.��a/@��V�����s^���=��ctX��`ޡ�#���xO鏙̔F�"���ca�B g����)�}�)��i.�P��a�	�$�Z���������R%(�B�5���{���PH��́�g�}j?]�[���*����b`A��W3��1"L�$�Z�q,�����l(8����q�n~�E�k�-��V���tVs��v�����҂�����`�]NP
C>�(&g��t74�S�ApBiXN9�qF�l\��1��ȊD\�{�ژX��Lc�V{#	ˡF�N�1�T�����x�Js�G���v�ˏ��
7���f���x �����֑í�!˾��l��7�����k�;�M�d���.��2�I���� \��b�MX�>-ڹ|V_��VFHEh���PY�ӽ;������3��,$�^ܚ����0<�ȽTI��a�a�ԙ������i�9��~8�]��.�R�YxX�rC�J�ę�YEj=$��!g`�"̫D˪��U��}�V��q꣼l� PKۧ�SD-�4ٴ�8���EN-�y��~�t�ğ�,D�%A_��&�Nȇ78��EGOĂx]�Z�\��J�����:G��u�(G;6=X��GWjk���=a�j�P�*;(6��ͩ���`mf��):H*�Q\����jk$�����KQh>k�th�X��\דw�� �4�	L��(Ø�tfN�VZ��Ue��j��t��c'��R�C����W
�I1N�yib@�����sŎ�=KG���B0�R�����WU�a��7�˹��̢8^0���5��y;#GQ�[��n�"��~R�̵�Ʀ��:<�'==�d���~;�ީc3ی��C��"����}}���n>�_.z7�|�?��I��vn��wD_�4����N�WA>B���{�� ��1ʠk���q�7�$�$u������2+��}���o�#,�I#��/����F�j
���n�OzS�lG�Z�l����
���=�&{� Y��r�.�k�e�E���ʔ�&q����4�,�]�P�.TO��8-��Q���#�G�R2��b[\�߬�@�B}�q�ż��SQ^�B&^f5�{K����|���k?��}oɎDF3�|��B�876r*�x��(-�T�/'������=��WI?�~���/H���'��V��r�!W����ͥ� �fRr�r���ǔf|]-:*F�3CX���qab�V��bԠ+QG����q�)̜�:�{�ؐ�8s�l��ߵL�N
�~�m���d1���Ag�C���8��͔Ľ���H�N�$aAq U�o��1H�����}�l�b2}S����,x�?ͱ_�T��ܓ�O�,��:YQ��;q+)fW��X*�H�t�1��:��ۯ	[S�<j�e�
=�ZOa���r������.�����^Nţ����0�U�a�3 ��|�{����:QX�Q>wd[k��);�����,&fy\�� �{���S,�8Р�q^��!~����]
�:l�V�`J��J}���	P2��ek�s��v)&�>zО܃| `�_�9�A{4�Pz�����YU;���7�*R���?.9�1ǔ��bQ��ـ���	���}����g��8�)L�������T����u�<5R曁�����!�,R48�EL5�(�H/�(�k�{�Khյ��f��X��~N�=��b�&��\�5�'1��a
nfp� ��;-xgRa�#�&
�DD,�[��@*U��
�+u~J��3\��zx]1=+ܳ7t
OW�{����%����Ɔ [ٴeB#��g�޻#�;>R�����;�I��O���`d��ڛ(B,c'��E[��,ġ��#Cf)0 ���kR�/QAE��j�i.��"=޹oB$1�*�K�#��Q�p?*�T�C�ӳ:�M(}�(�:-���3:�4@���#-�I�ӛ���i��.�Q�v��[�"7v��c����!��J>v��4�SDM��+hV�:��7M���D�:.��͗\P���ck�`��W�������1��o$;�yN*s�`|����P�kw�����zU���t��	���؎9{q�����Mx�R��$�f��񮙕�GFI��s��'/���H>e��Tx
��Tٱ���is�|�v��e�t���+�VX���}��Q:i$�i���E��9�(fb�a�}��>�=@��U'u2��N� ��P��H��cZk~$t9���<�]�	Gݬ$s��b/�}��Ѥ!Ʊ���ڲ��m���~���U�A�0;r�Vr��300o�����*Z��s燜���vW0�ԉ��崯�6<�As�'!|�ᑞ�PF�9�5]𺹋:c�B��>[����/��@u� ����'�?ql]q�M֋y?Jb��Dph�,T�_���0f�7�,��{��m�?��醪����v�&�8�����c���~T����3G��6�j���MR�b���r@�1�\=�C������\|
���܊=�J\DN��]���?����	$��%]��{z���}��c���R>�]�,���>��T��	�P�8�>;^f�� 1���r��f�o�=�)=�;��� U�+h�����	�b�QqFj!�S~��\���}E�Ȗ2��7�`n�e�E�#�l��i���P����9���/�|b%Y�4{s2�	���7�>��h�H��:�l�j3,�A���-mn4r��TM��M©��?<��[�E����Jϵ�V� 5Eq=�t������@}d�1���&ȅ���'��G����3�(�l+9�AMfC��=���>�"��(TR�ZoE�6p:��1_�萌|�O`@ԭz��X�ߋ�>Z��9{� z�Cߧ�%��ՠpR������Z|�)���W^Y-kr��Y���-4���Z��ED�=�ތ
��1{��o(ɱ�;<��&��$��R]��5fY��8�7�KS�1�*�$}e_�!:�A��x�'kQ�j�m>��[���.$����^���ϧ��l�|3J/�:�r�3x\3;Ґ�\ڽ�JZ7YpQ��f@M�x[�!��9��װ��"8PV��=�ׇ`��@V3&�5㊤���' �с8��R's���:6��9��My2X�d���ֺ�q$�|/ ��L���� '�+��e4���9K�� ��jO��5Hs�<���r"�� ����U?S�<R�<u�]��ռ��0]Vy�н��`�a2'6���en�B�Y�����r��d(�"�~�:��J%Z* �f�*�+'�)ߦ��^�]�hYr�� �R�5�5��$����g���}�>;r����w�}�H~	����z'������p{{�L���\Ξ�O�cr�OďT��'���"�����Z��v��OϺ��-��lЃ��C�{<�i���R
���i<��KIdQ��f�@$�˴Hj���Yྯ�B����\�^� #?'�uݍv��^����&��L<W����N�^��癱�k�8�NPn<��ۣeN����<�W��t�N7�഍R%T���5�n/�3뢀x�~�c�O�B�vڱn!&�=�ٰl&��i[�5A=��$���^`��F�|>�o�gm��ue�"uELJ	�M�">���YEϘ]�����$A�����x�瞛�ٗՠ�h
�Ph�<��ؿ�YbG�Y(�`���bKW.�e'���̫x�L�]��>q\Gl�����|T��:�T�O�Vo��������ϭ�&��|X!2�O�l�ny��2�p� �c�`��+�r�UL�B�?I�Ԋm��j�u�����1�5���u�cAPEpfհj�D0�\��� �x�܊L{�SB�޽��A�����h��|��y�D�pݯ��PI���Ja��x/�J#7J6+�!ރa|�n��S��HYhϖ=E:3�k�N����E�>���.Z9~�5�W���_uk3��"�� �*!���L���2�[���hd��{I�UD�q��aUG��p{�=�.���?�0|3"R<=OS�O��u�IL �nt�S��H�����nl#�5E��p����&߾0��I�1�����@O���@���Ti��mV�7c[b�8R^hN�?5�ͻ�x]���}n(�~s{�*�s(xԜ���R65jQa�D�9]g��d� U7%|�0����=� ��'h|�n����F;��I���w��2�=���,Qs�!+t���C�q�i�yab�e*����%�`�/�$N��.�6y��b@1����'lT�s�N���z�xkJo�{��_=ٲ�Y?��O�,�qy��ܑ�2��ǔ��k����3��|\�M!x� )H�.w��|�`�X��"N��!���+���q��*�)����v�?�iO���N��B�a�q���&�)ԇ)���z�P�+��ȶ̖���:�ّ�t����BP��v��T�$%6�{��O�����6�
�/H��";�(!ʐΈS*v����|���&O�=2G���L`���Kڗ=����ک�*�f2��#��6�ZðE�i��Y���|���%�ֱ���:ӭ��mV}�v�@v��p	u�U7���
*F��L�ek_��P���.r6�5IП0
�K�7!����J�aQU�&�V���l��3 yct��+��i��`:O��e|�;b~�0��f��tJp�Re�Yޑ�n���ߜ��i��'%#��Y�?��N;s+�'1��ewKĭ��Cܟm,L|d�l�g��R�W�Gi�r0����Nа}݁�J�����Ywk:y�k�^� �����n�:�*�K��<�^N��}5�%�7�A\7��R�OT�0#{��ø� �&:i	?�ce['.�'��[��q���������5WM�2��FW�u�k�ʖ/���.I�����3��? �]�[����U��O6D�i�� �{�Pk��/���_����dv��
���q�?oSB��ѣWdp�߆�]���e�=(J�NZ������X��XlC���ߙqs� �?�v*�����������4x�S	jQi�P�ǜL�4��66S�9h��p`aG��%	��.#��]xO0�O�D���
��Y�9�{��R�ʝ)���!	��ʬ���'J�'‪��j���\
��S��ԫ_�F��W�2��#u�f��,�Սs��Vid��.@8�>�u@�ȸ�u\�8Vq-}��fT�}����Κ������Kz� N�9B�l�-����> �$�&�q4n���S���q��NO�E�&���K?��ڒ������o,��������A&��N���U�F&�����2��[��Q[Q�\�0Ɵf_;�@QBB���)��c���F�"¿ݫ�`,� g�d6T#�.7�RĶXI����8q!�0b�ɂ��;�ql�AUr?���6|&9l�@�	�=�cPFo�ֱXE2�]W�`�S���B;FS+���	|ܒb�2`�W�o�M�b�{���/b�QWǵP��P���:׋�V�&"wW�[��"�(0�X}>=UHF�"xh�`�M�m��9��ضxR'Ia����'_-B�ؖJ/by�mI0��u���C/��]
?͆S2�䶭O�$f	b�b���1RY��Q��e
�M�ʔ/`����7��(d�Se��E�燰G\;}� �ȟ&q�:5��]�N)2�z?�E�ڞ�C�&ee�KFf}���j�fc��*�Yky1m�a�������`������Z��G�r|�w#��B�������5<�O���s�Bt����5�ݸ���
,w�m[l��oV��LHfq�N5�;�<ty22�@ό]	}�_�Q�gTb����w�Ϫ�M� o�!�ݗAi�t����NP����ۺ�19�9��UPy���@��'�}�X8��S��m��_�;�^�g?"��k��=�J\����[�����a)q;ƴׄ�5�5��Co�Q�$E�'[�X�
�j_�ll�1^�b``e�	̉G�>�g��&ܣ�wD��*�X'���v[k���,�v2Bp�va��@e:� ��X�/�X%�? ��vSK6��<'Ӕ��Uw�O��%8t���{�p���)!�FIo6�w����nO?��i�ޤ���Ԝ� ����qR���b�����bO���m�t�
����Ѵ_��,��-A�>$ ��]���i$F�b�@k�\�=?�-S�� Ҡ�w��e���:��[��U��f�.5p/.�O��ӗ�kh����A��U�д��>�q�m)<�Ȃ*��
��܋��q�2V��L;��U��o�f�����qm����	�nq�\�eX0��y�x����_����Q�6��>�.��u=���jF�4��i�͑fn�T9d��H!��&ޖ�1M���a�ٯ��z��*�A�z9v=[+�W��"R�;�7��	�UX	�S%Ve�p�Ċ�Y��S$�a7��f<EWX�*^���oB���z�e$�<e; ��FH��.c�������(Y�P����[P���s��XI��{�g}�����v�'��!=ز2���)"��ꨲ��O.���i�e)�{*ۉ�$'�{~����P�:�����G�?I�U0�
J�flV���@$���V2����'��ʑ�Y��$�
�"\���tA��bc��YKv�X�l�3Js�4�\�����z	ܜ�!�G:�~��pH�`���+	"ދTCI����U��$>�-�E���F�~�11��{(���;�����:q�q�E!��� �	�i6��X!��S��Z"V,�t&����$���ʤ�"w��a�C���Y`�E����[��_lFs�TĿ����v�_���i�NP����w�N���sѝI�ۂpaHe�봗��W�%���(AL��@�s���q@H'�*Xά����M��dL�sM醹��x@���(��{�:+�L�4 u��k���S�����W�!��>�$ z��˹�ei�ۧ���^�9�F��%>���9����]�������!T�t5�1* ƞ�҅`y�.�޳ZI:Il�+�yj��n��I�%��X�D�Q�a��R&B�GL�)��m=`�-�����/�)U�ŝZ�<�U���:�Ro�ֈ�F`�B�խ�oP�o��H���hN $�C'��[3�~00��Q]hJ��Pn��2�T�}iе{cu���ȝ�z�I��Q*2݉[3�h�<1XIoݡ��4�B��z�¿Yd�x�qY`��tR����j�=�;�5>-���@Deb�z����d�h�R2[�z�'.� $�u#YC�c��H�?� a�h{PRӉ�b��%4���Ί����dN_VQ5{�s�4?��()�Ms������D��&�����s|��t�5`�G7J��ۇ� |��jH]�?�$U��,D}��GL�X��&�[�Wv�#d4?���F4��(��z0���4��q"r����@ǔ�V�|Uְ�j<.�s���hUG-�@�������>��bq-<���%�*�(j'|m�p�T��M���LW�`� �$�ٌ< �>�sW,;�80?�1w|]ȗ����ɧ,$��R�|����=D���f�9�����n�u��-��H����Ƚr�#ۯ�
RP���tD,%��K��2/��ug�)�l%�&ݳ�_Ki;�AL�)�*]��h\�F�O��fIM�*cB��Mu��B���v�* U�Ѭ�����)�1�Z�����oc���k���PpWZ���Yv�����ڤ�/f���=0R*U;���m̍}U�/�#8���"}VO1����1��%�6� ��75��tr7)u����َHb��<z�|�h���ɘ$o�h�����`n:�y n㷙C�X����F�!�u���{�u��Nb��9�LgɍXv�M"k��1��	/����w5�iY�z����5�o����%�E�`��G�a�m�~
�������I�𽻊0�:�� �+�YT�Z֎+B�%"GG"tv�����c4N�>�%Ϝ8�ӎh3��g�ː+�i�K�{L1�ff%��w��(�Q�	g�n7x�)v��@B���7V�H����;�U���^D��b\C*����:?P^r�㌰'��j�ZA�؀�2K��,��F���b+'��}�V,���7�\gv�����o�����i�R�͇�'���d�V�h�ry�g�@�s���Ѡ_s��xf*���9ׁG'����&4��D�"�ħo�"!���jb��(5��{Uo[����^d�X�?Ǳ��#���hUr���TM�c|�G���1���/N؟�xT�#��Q�ٓ�C�ኚo�q؋5EIb>�c|�|�K�gxd�OD�~f�A��Tm�tw�/��6������%�����[P�S�{��H�/m55���C��,���g����I|������\����x��w���x�7��a��	f�%Y�6r�?0�H�V����y��.�����Փ�C'7�R�2�'�(R��O�����n!K�K#ʅ^[��=�L�<RP�)�}):�!`�H���b�ֽ���R��5�e6�� �6wԉ��W*�R�-�I��]U�ѩ��G������ea�O����y�.�s���3^�9m_���
C\�zە�cڻ�M��Al��?���!{��U\Z��<��D+U�#;�臍��xV �c_�� �S��ѯ!�I5�����fz�W�D�#1�O��73�'�㫮����K	PUe8�r��K/�Ms������#7[~���/5����+��e{h��o.��u�J���D�ض$0O^��<K��b	�G��݁*	p[�?���(�2y����+�*��D.Me�cc�QXŞ/��uq`������tX��o����'������/�k�����42�YN)}�r/��G�>>}P'�tnK�bZ�$H�G	�zp���Qzi��W��2cg�?~ā�t�Ujc��s�$C�� �+��_�G(����U�����~�ji^ν�d���l��fc� ��P��T!��aW�-����P��~t�d���cV/�횡c�
�O�4?���}�Km{������p�=�P��k��K�`{4�I5��|�*��L�>���\/���o%�Ԁ�6ȁ�餞T��z����~��ΐ�F\[�/�I��f�� yKTL���?3XoQK��3��@Ks�O��(>Dڝ1��!��M|��S�Dͫc=�4�g��1Q3�n?�·��l#�w�5�=�}�|l>Q)a�k#��/�˵|w���XD���J�si��s(�q�1����j��|��T�֓m��ծzl(y)�V�&���聘v��zWB+_��n;���N;H߃A/�����*�	@��ꠊ&���p��F,�`Pt�$K��d�b�2o��`^C�+%�\ت�5��5r�93���X<)ϐ����I?��/�z�jU������-����:S�>W�M�@�nl_�m��A���m�q.m��R���I>�+�h>�?��"��#<�m@�n����։y�[�2�r�^�ĆW�̏'!kM?��-y�.��8�ݞɩx v�J(	.1���e�dU�ǡ\���&��Ĝr�$,�����Q�
����1��:�mR;��"�E��2�,���Q�� ����0W��+$����U7����gr��Y\*�r�	�@Q3�)��M��0/J�[��=��|��|KM����׬g�5x����F�vO����r�7 �^1�>�,�5H�{�k��e�e^���^���QS?�g�����z#{\.�D��Q��u�k�7�����ۥ֯M��,S�������_���'$.:P�������^1�Ce�/Z�i���u�)9�#u [f�yi���C�̥���§�����p���G��i���HR)��wmRb�Ӂ�.�c�k���.XF�ke���Wt�g���Z�gB[*�Ӄ��r���F�� ��N� $g� U
-') .�?������E�y.��9+([�t{���2�"���fC���\���~e641������y��$��J����W����# ��RN=6�'m:���DN��	P����Y��-����ds��_�A-�JR��7C�9���:b�h�P�G/���� Gp �x�}ܞމF^��zJ��}�޹��'���S��:՞e�a��o_���/>ē@*�����V��0�(b���)z�j�h�����Ю� wfo�KV�b�g��M����)���|a��g|?��eM�fޥ���iPn��C�_l����cUu�9kӳ�F.�Q�;ܾ_b!^d�V�mC�cU^�H�#�����e��0ǣ9��k�n���
��HC)�%��Q�|�k����O~p3��Zd�FrY}��X�HG6��Xܽ�{`�먿M���(��TR�|Xu 㧳[i����Q�#ּn5-U2��D�i{����[|�|�S�<ܝ�,���ύ����;�-��Qx �x�y`/����Un�\���}0o��%���`�p�&4����E�J�[-�����+̓�����N�2�9˺R6��4��h�(�f�	���]��0.q�z������aPt~�Y�"�@�8���N��?�a�3¤�Lʜ5Wڻ�`���j��ۼ�����)�I@S� �ℤ�P��Pݧz=&��qb�Sޯ\���)������>�W!�.��W&���`��b�jXu��r��j�&Hjx�4�|r��F5s�My?#���$0'��$0�b�F�㶟]�	����)K�G�0-�üY�T/M9�܈�6gM�Dcs�����0���*O��T6�訷ntiO ������Ǳ��?�毨����fC�
�������R��B3tɤ�=h��sb�֗�2p��U�d�-��:˓y#�J���tD�z^��w�Ԑ��Rh�Gd��	�7��������]��g��MPx|Ps�VX��+[iM���Ʒ�pV��� J�|n����^-]�B���L�d��qmΖ��	خ��C�^��|��^)1z�G�3/�*�.��i���X���������m9���֨���~�~���NI	L�6�������+]�]���
�1Y]����b�?�>=���)`�;83bԀh���	6j�W���4fZ�m޻���\��ka�+|p�7ƥ���n6�'4�QDw���-p�~Ǻ�c�#��ƚ�A��oXM��8~=Re�Jd�"C~��h]q�j�r݄�y�]�$�E���K�̭⪫��&�E�(�/�1"�B���
Lm�u'��e\�1:�m/���in��e�$�4�Y�(o�ʾ�q��e3�p�A�]�X���f��E�*!�ț�?[�̿��(�PekD3��p�d�4-$��)?�En;�X��#ҭ����`L�*�џ�f��S G
�y�h�p�kK7xh)�A���ӧH�]������S�*/`�J vd4`D�M�C� 밼�Fu�Ͷ;D������ 5\�@���T)(�"��y��_,[�x#ư@�Z��p�,ޮ3'|��`6��O���9(�C���BQ��'�َ� �SVXx	3r�-��QgU8Zص�y�l��8,��XIX�+�{q#z`�n+�%���ƥxڂ�C��P��S���(Bt.�,y��+���+n/�L���p͊��u�@��l8ږQ�����͙�1-�۬
HEP�-� ~΄���>W�:Ֆ�=[(�����@���dM�gѣqDoԽh�i�~b)�f��O^VZ5L��6���J�o킽��g�~��e������k����C+ϕ;9-k��[��J�0��q"����m��� �r��B�`n����h	��R�@��c�� ��A�K6�>��̪�$�W)zI��K>���:�_|�s��;=#lq�%s�@ez=0�;��F	�)/:Va"������>D�*����} ����Ϟj��7D܏W0�R9�rI�`:��?xv� �����l��
١?�FL���O�u�vƷ}����'��4V�@��+����u�W�Y���1�/��{1*�|��e^1���Gt�\[���Af��)bs�����^W��s����3@OK����Ɨ޲7��p@��s{�|�a%�]�����
��`�
5>w��/��f�<r�0��p}�)���߁|��K4���������םVG��KV����o�i_��U����Q���N�C
��0"8J���V��M#oJ���vȝ�@��X�g:���R�B�j�+����1�n+�M�nn� ��'�����V{���#R�U�ϟH��`��}��lS��$���)w��F��\ؓ�2xu�ۭB�O�9�u}i�_�m���/�y
�4�g��"��s|��%��Y$r�b�m�gV��%M�J�'�ap���>�H(7�� S��`@y-�Q �ڰ1��:�BR�9E�[�v��h����[콃�I������nZ���z�n��i��f��ӓ6m��)B���؛�E0�$���C�Io%Dԯ����B'����|���TL+�d&����J���E���D����+sB":t�*�r����+�z�_�j$q`N,�=���7�@n�Ѐ�C~�6���H&�2����Nk������ä�z�||XE}��*�>A҆����:lj��*8�;� �K����j����!c�A��E��!�h �u�;>� aU�v���N������)��ZCj4�El�?�Ɋ�PT��eŢmF*j�(@_4U����]o]S$����ė��M?�*g�j�ܺ�Y�}���Ĕ�c6k��f[sR1V����>^��S�e�E�Hl���Y�Ҹ�Ղ%��0���)�9��$�Y��hkFV�&��x"�m��N�vV9��#�����>o�lҐ��-�a>f+	�`&�E��A��.(a�˽t����>.J��
���.�*g:��sk����wW��5S]]�Fcѹx��Τ�pp�VD%����k�q�b�ʒ٧��%�dZgFNN�&��<�eQ`8Ñȭ�?��^�u�A.-+F%�۬�CE���i�����x�����">���q��ޮXGF�q����cp5M�V�5:`���N�$��'�
UfK�%o�"���M���hj�fLD;_Wi�#�'ݩ<a��y;�vٞ�,���/=C�{��N;�r�����*�O�N9Ya����~k��_��h�s���?b��ӈ2b��[�X�F��t���I5q�l-t�_�EƪL��qA�W���_޴b�>�\&3�3�zq�Ja���y�"���0��=9��3�C7m�%�ׄy�.�U�)q4��� bg	q��ѥg�����@�DDy��%�����n�~2ו*w��_�u;�����7:I���K�c�p.�a>��/t�1\aW��Sf��|�5/Vx�J�\�u�qiv���`{|i�$S�F���S��x�� ����8T��t1H{em���u�$�XP}�50���r5���u� ?��4Rf�+NR����2���v;ۂ��1��";�w��y��p)��-('Q��	��� �y�G��D) ���TD�,��D���z�%F���8��Ѿ��IH�k{Q-kl��?�%�bS<�Z�H�M�~[���D+/��F��=�5�Xp�ke�����1]��,�,��a6;���Ta��:�3�]z�V�;IVs� gk�Ven�U����
�C{��j�Q�tF��n�nG�$���!n��u����W<� ȳ�Gtٗ���D�Y�y�ll��'6V�~��s� ������}�Og۔i�l�ZU� �P�y$�u5�_כ)�Ǭ/ p^���KU�9b=�Ш�Qi�!�O�q83�V{Ld�\��+(�����{m^�+�NFX��m=$�v>3]��ߝ��%��,V�t�7��zne���!K���UO,�y��]xK�f�C^d���Q�K��z�P�f�/K��t�Tp���)$�0�0ᐇ�	�~���FqMB�k�h'q�n沷�4Y`Z��GPM��T9-�+����GK�Ӟ(����I��ѦW;�&���]C<Fj�q*�����j��}�qH�:f:*����t.�/9��A����:�����xL�\�>�HN�(�`
O�����T(g��^��3����]¶T����".�jه2��T� Gl5�&u0��bQ����g��T�|���XU�vl����l?��$�{� �#-'���J
����Ѣ��*!��HW��NTR9Tbai��D1� m�,��g珹�l�\�x�ﳤ@V��{i���n`�"�T�ˑ�a�Z����3(�Eg��[�@DK\�y�y�4r�"�Ź�a�(��;W$ڜ<;,\�g��$ǫ���^L||)X�n�s�m��ƚp�۠�⫍zt��ô7�������fW6^)�8�c�E�Ԓ�b�*�6D!��G�yS�w���`'�
���)�Fp����Wͻ�����׎ޝ��ל�����aF� �|W��g���% P�z��s��
�a�`N���X�B���J��΍�a����z�#L��k�f��M�4�M4�<��:!0�7�;Dr�<�UQ��?���'c�K�ҎR��n�����C����Ԋ~�<6�`D��_��Ar)�n��6֓,�J
�����Z�4M/��B��[1&{��U!�V�����X�҈��*�6
5r���'�k�7	�XY�k�qiv��7�T��	�������ݷ��^��6{�����"(�� ����(XF��γ����~�����e��D��IN��� ��$��p��	F
�F1q!�ο/�~ls��g��I�,|�Y��(�ئ�0�
���>�^P��&h<��C8�Ƙ�!�A�$Q���c�Z�x�y.������霍�r ��q��ɘ�0�w,���[�Mup�
�U"������)P�,����3^�$o�b�2���(~���/���{\y�;��?�RC�>�6T]���۠l-R�����eA@����P{-���LOt�)�EN���9�5:�G����EV��cc�<��hx�%¼�M� o�#�*_����`���A��{���S/L���G�d2�CQZ1�4�&vgX6]y�]��0I�1�n�>"��^+��꓇ ��?>�ntISu4*��̖���ͥp��Vs�0��PZzBT�f��ⳑ�|9 sw�/
R�XA8j-��� d��~h#R|��=�O�
�ɲ��M����n��:����զ�6.�g��	���d�����k��2�����EZ��A���ey�rLpP�p���Z���zuρ�WKS�1K;h��裹��.N9."� ���E}�����UM�EQ�q�rJ�(%@���&�p3r�?�P�_	(?�M.9�/ΔUQg��ڮȋA+�����'m2*{������Z��7�`���!��>R�$��:@���8��%�/>+ʾ&Ѹ��lE�⪰?D�W�	��Pq;k�6����ʽ|���ŁCd��'�$G��R�T �M�$]�I��/���~(棎u��-Z3��	@Uue�����)��
�$0˓+���ȹ΂Ŭ+�i#iHs�����w�hK���x${�Y6f���11��٤��j��?�D��)���ѿR��eNێ�M�<�:/�Vj�!��M�kYj}a�ils�uX�A�=������~��O����@j�"���gi�f$j\���& ���?ī� 2�b�_����uO4CN��cD�
�m2���ΰ�2�6�+8�_�_sw�z"���ߩ��RU?�9�sT���L��-g����@��<��(��R�����Mg�H�b�Ʃfz���[�%)��e�9������� 5I�)��/�0���YK�\cL 5~��o�'��nt0�TZL R��~�����|�������{�7x:SjU�e�EUn�i���2za�1F�ф���PU����Ŝ�nV��}\)�g7#�Dg��S��N�Z1k�j�s ���B�8�O��x�,�i�h���v{��-��0O�?saU�C����|8'�>�>v ��p�\+}��	��l�e+&vP�c)��8e��Ɵ��baf!"{���:~l^��ݦa2����a�	[�=���t*�Њ� A�$�*G���X��=^�M��#e��F*�D�Uv���ٕR���Z1_4�h��j(��I��zɩ:z4v�xg.�8(hP��:��fݓ	�꺆yrV!\ݡP	�����s@2��v���{̈/I���T��#� �i�]�o���-��߯�%�[��F����O_����սc�=����`f�-��]�I�!>O9����u8�H��v�΅$�Q��j0�w�����a����'7���#Я��is��̒	��p*.������؂.y�o���iz�����Al�hC���M��H��p�vN(;3\�r1��YwO�J���	�|�Q�VN2�Ӊ�7#�K� �g˸r ʋ.%8'�բ�0��
�ׅ ʾ��B�Dq��@�f�g.V\zn���/e]��$��j	oj@aj�f��L[����fS� �c���:�-�t�f�(Y�MGg�iw�Z�S�L���7��*�Q�4+�����#\��}����u=��sK&.B;k'?a�Mn��Un�S�����s���>qz�( ������$t���;�����%߄�l�K�̺@J�e�X�D��Б\�jN���e)��&��]��s�A�W�oE�p*FrFQ*�3`]�M,C������T��W�w��$�<4�;���|I����c�%�ÅSPQ������®
�6TM�m��ȧ�ֻQ�7p$��#���H{���+��V��d�e�kb�4#JveV�����&v�O^8[���Zi��6}	�,j��;�솇�V���"���!��Q��|�pn������C˭k�ī\]1��bA�h��ks�n�Q��. f�hو�����k�J���$��e���Y��*м'�^�_�����W>����Xg+4�OGO�lu��Ux_Sq����aa��H:��ClX]{֜İ�w�<�|�F������!��D�J�����;���x����ܱRFPH$4~�xN��z��,�d*�t`I�7���l��ۭNV��ng�~AlT��]ڃ̖x�+��5R��� >:y���h�Y5��}�(�5!��d�|p��`H$Qh�F���swX����?oV�h��`�k��FNaM>��ns�X�k�h���@P���$� �)]#�«�H�5in�� �P@��hΨ<��w��Ů�ޣ�W���տ&u05k���#-�ĆQP��{&�/�F<��6�O�]���=4��,E���Г�Ť��/�mKZ̺�7n��h+B�?�7ߥbEC����:�u����u�G!��{�z����d�m6�	��pC�-{M��P�K*�iE�2 "P礶F������u�<0��oK�Z����Ś���#�]A��i��[�j�M���3m��[�C$'0��4|"��`���q��eSGn�
z� ;�\t�6�5s��!�ڣ���DZ ��'��Hj�
��&)�1�/��y�K�1$����7�M�?��m�XW�8��?���i+��nL�t"FZ�r���1����A��&��3Ǡ�tԴ�����;���Ki�/���i�U�%$��C&T0g�m��Ԕ�`�#���[�:	z�>�}荹M���n�OV�]t<9�s�S��W+s��vݗ�d6V�&W����$������d|E�0rW8���R�X��]�tN�Gme��d4��;X[��Q%���\��f�����U�	3�i䜑mkO���腓#��X��PWQp���y����4R����ˡF�a�-����c�\�׍��9�����]��{a���.:�?I���3�25�l8ɏRm�Լ0��z���2NFR���Ċ�&i�X��t��z�N\���~Z#��S��<W�R�T�候��J-�r��&c��� ݣI�P���tq⨊��	�Qȋ���Ddȿ��5/P�v]턼йe�֤Oڇ��8��R��ϕnz���	Պ��wV6���S���E�;*�����r�k;<Y�����ps�����O-��7$9>0�����F��Y���q��p�־��<2��M#��!���|�����t͊�.�x&E�d�@^�qC�і�&>�����*t4�;J�j0,�؃ǍWo/���3؉%/W��!B��I�/c���``������*�,1k֕7�"�*`��3�� �BM���]��H�tV H�cVP  �p�����F�(]f�8H�b!_R��{��W�{Y2��1�d(45�{����� �xj;���?�O�6?����n��8`�5�!�o�ڠ��jd)�2ٯGy�ebL!"\J$aaH��#���3����m��DW�N����N�#��{Jk��.w�˾q���Zz��7sO���bK�8 ��u�"�Ť%��Y�_	���Wk�s�}"iW�(�����ܼ:��irr�����$�>ɰ$����1+;� '!��P��@�Q,ߒS.��#�S*n�EҺ�}d�>���m@ ��Y��'��/-��6�N;
y�*��_j��FY���J3l�����t���z�a�a���4A�51������h	ƬP�osP�Yv��F�B��-���ؕ��9ܺ/j82��4ݪ��%��9����m����'�;%�Vol�8��� ���«��"���T��4��+R&X�L�R��V�c�n�7Ȗ@� �~a�%����:X<�BX����@ρ#�2��bJF�7`�(�*���KQ	*���}H��vd9EU���Vd&Q�� 2��p����i��`>�^W�=�N�iGz6'�%!�vjH��N�]L^%�Ro9>�'c��SC�y_�`[�JC��Gs+�#j����*Rq#Lv�Y���~�dB��� 7l��2�0�l-�?n��T�V��񽶺��,�R�� 8�v�&m�ZV$K�~r�\6�OB�f�۸���T�9�{����*������r8G��n�X'wh6~�"=�nS��R����w&��(^m
(c,ly��~�_K��g�P�Uo�6�R� �S�oJ��&�K��B�8q�OI�\�[M�/��%�I���������I��*�}�B��A�6A��]Qa�3��q�KA)��mH3d�+M@tXC���e��vl �k0�-���M^��{��N�S�'-Ȕƌ��D�
���)�c^]g6����s���an���M�8��wKvD��f�?������3|������	����%`J��;��a�g�_��7w;lS��\�]�:�9�= ��r�)A���@����	P�D���(n���hg0���O�e]��L���~n6c�H�S.�$����]���i����KE7֋%kZ ��'=P||/3NuU�������K���ܸ�通�]Uz �����Q��E�e.�{��#�tSd��t��&d#ݡ�����r!x�c�{^�"�h&�9T�y5y������U���"��O��D���>����SH��JB�3��+!e��;�^�
�W藼s�������x7nҝ���F��pNF<��0��gC��-�X�|bf֭�I�j6��b^F#.$FJa��e����"�M�[F���q���5�ȅ���ELU�̂M�񄏮cނ�����W�VFƾ,�6C�*��'*��&ߝ�KQ�=�.\B<aW�k�<��L�W������Dg��db��5~��2�����奼kI�5��M�6�Q���͆SN4۳��iL'��=o�+�m���'�>�Ϊk�mn��x%L�S��b_�xe���B.�����+@�;��w�2���C��!��u����/ݭsDN�'Pkլ�q>�� ��e%�%�7��J�|�@P�IW��[�.#Cs�	N�*�Z��ltN�,���Mg�G�,��s���	l9��,����$W�0E(Q���K�<u�k�>|?j�W�2�@�GLz��X�Ss�D�F��(9e�������R�����+�3�r#��?%x���Z[�+�=�l�L��NI
2���#2v���\UQk�IQӟ�j�0�����	o�wM���"Z��KA�/�H4~zZ�J�iI�ہۣ�Bf�@H�)˕�߁A"��]����:����fO�*�d��OZy�Z,���4�˓h^���#xN������H0�#t���aT�y%^H�]l�q�3�;�BʐN�������o9'=�Q:��:�9$��Y𯍻��b�D|H"�rM\����"�pBG0�V��IB���h���,���O6
��}����)��JO��t;d� �f�Sb�17����n�A��N:��r�{Y�[�rʱ�"�7:"��fpJc�-~�r���	��$	8�Z=3��k#-vDjӔ�0[�X��P4>e��n����(\��F�|��"���/@D��5�Ǥ�&��#���)�mb�`̼�7�EB����i���e΢T�O���6r�-R@��@�	�F����ec�9l�Z>�����.�:(X�H�d]' ��V���&<ݢ��QH����Q1����ʡb����S����C�,���9�/��S��@U�������u�vSK�r�6-ܥ�dm�ax�T��Id��d��	��D�`�G�Hp�ō���T�]���[b��\*{B¼ʷ�Ói^�=����N>RCu񍵐A��_��^c����z������x�V�N9i��A'#l������`p��~X��v�ۼ<���/8O6��ph�!��ɝ�RFMӇZ��Nd� p�bҍ{@V�,�g��Ņxb���%�A�a���	ئ�Djg�,j����Y��������	�bF��ii-��5�յ���O���)�n���Gq��afq����ڵ� �\g ��V	D��h�����l�09�P�H}�ɾ���7��ƕ���Y��Ư9w���4-��>;�j!	��U�c�/�#�AP���g�����X[�d�����_8��J�ь��qq]=64����$�k��kBR?=�&���M��L��h�f\8])/�f5-�6��P�r�n��V��S�z��9���T&,��O5���s�b䖊�"Ք7y�+��-+��D�0:6:%w��/�l��T]����~SFŚ�_P<ǪAU�:@����7� �P���v�*_��hr�ז���g<�fYӮO+��\����sju���yˈ:�J�|QԱz�ϭ���E��u�����vJg����H���B�%Y��	Pd��h{鐆lR��ju�U��ח�Nb�̻u����y��)����/FΤ`���om�U��"s�K�RV����יO���lO=5S2L献�>-8��d��AoҼG2��\]�-XA��]�Z！�~k-n<Z�����K\����n!z��?N�?�^��N�F��q��9H7�p �s�иj�]]��)5�E�jiD�tl���b+b��t�ؐ�:�*�(Q�g���,�d��9z���	ӭ>x���Yy���`�gfI[�*}�c4߹�$Ru�JtУ���"z�;����th��[`�"���
��)��(��~��J��M��F(�Nv��u(���M���6<��R&� �����$�o�V$߬ۦE�g$�Ƿ��%��Р���-*L#�V���w�5T��U�6�9g&�!.��?��>p��bA��o>WP
���?5��8�;����w��)�V'H%{�Oא;����hh��_�eǬpʣ#Ϋ,��.S�/�mأ6B��@�~��hČ\r�#۬�yQ�B��,�9M�niA��I_;��co�(I�C�^-��
�z�ث�ʑ?#�\�(_�ObO�6hY��|ٰS��I$D���ռ�G�jo��O��"�����.5S�^&�-lpl�BU�z��w��=@�뭧k��e��b>���Y�o��~�N��}$&�if�,y�e �	�_�''�n�#P~Nd΍�cf��2��(X�D�ޞt<��
�.�NH�̋J���)��
\�~xؾ�A'��?����3>�xg��   6�N~��C��=.a�;��X7/$�p�`�u����ۗ�.��F�qEL^#����A��:"�P>C�n\��H��,���T�#�â�e��z'D�y�8��޻�u�%B�r���¨��ʽ�DJ���\ZĎ��ڰ����7+Z0������yKi;�3����ȋ�q�Q��2XI���Nۣ�"���p$���Mg����O��M�R�g���t|��rr�K�X��|�E\,�V�Φ~��������*s�Y��|��ނ7K.]���ʡ���V@�6�3����I��<s��AE1���<S$9V~l���1�i�WFXo*^�?�����s8 w����¦X	_#D!�-��)?6��7	?{��f�Q|��OCX�_8e��m���|���O7o�dN6AAEV�4f�@�j��{u{Pf{{;fv0�=7qF�v��`)�.3Da��g��&��r���]^ݳj�a1��v���;`ز �	�J9����Ȇ�y�Ce���p��]��"���Y8M/�q�Vc�N���0���0t!�-�##��nߓ����R��A��BWZ����b��һ�vE1��4��a��O��� F	X^�g����}�p�@�w�e�!�g;w��D��c���`l��nO��2��+2�cƻߤ<�NEћf>��uc��
�h�EC<BH�Z�V!��{^���ۖ����i�:p:��։�W�7��B�o{Z���c�4p��<��'x�^��r0�m:�d���J9�v�3% ��fǦ��� k�����,j�6.V"�`����GA��=��Ĕ0�W?8���"?Wek��C�V�grWѭ�5_*
�DJ�NJZ|S�+��l���^	�l�6��#Ч��qfMi��34{T|��a����*n�U+mP��A���?}T�¶�5D:�_�/������vG�A����#�@�0�2lw�q��RA�1����)�?2�`/�]�sQo&�uE���I��s8i�r8�E��Y��h�%[Y��m�A<���+�i��|nm�����'�=& ��ـ�I5)q?��3���$��`���g��u �x�l�\����Дf��Ԧ�C�sPPLW�P+7{6Mo��80�+֚�EF7A�u��({��F\ ��=�mGQ>?��4N����拸Z���x��Sq��T�1V��kC��_����!����� 'ģy���A+��}'�iF_#�F�o{Ə��L_�_�u�]��ҥ	JD�NŖ�#*���C�k�-��G��x+�(w�|-��Rl"�7��VOn�B�,kֺUB�}��>�Tv��C��o�g>@����¯�:i�t6���?�>�;+^�#���<��`j�l���A"d��'��z�١ Z�{��Y�l͈[�J�����eBH���b�h@�s�C�sFx�p�T�j�4�,���6��k��!"R����#����k�� (� X[���:��$��w�4�2[�C ���!���&�yc��j_�I0�<�T�ĳ?Z�Ʀl���k�(T��m�^�����{�/
a��\��£"sh4�� ���9V��P�bh��Ӣ�њ?옎�=W:4��n��ħd�H����|xí;���z�g{���OW|@�M���yh�-�˃��*Ib-����4�	����6�_���/Z�@94�yXJ6�{���`W;֥�5Pn�v��3�;��&Z?�-�������I
@�U�7#f+#�27�í_��tg��	
y���'�	��f�tS�E�O��-��[�9��Dl~�T�����ּ���\V�1�6�=�����s��wr�8�a�&r���S���b#��7���KoȘb\��:�Yݸ6���Z1�XnD�3R��w���G���9�5��R��w�Y�W�_�?��\��h��*����UO�K��x(���1a���,�#�W�Sn��]�!�[�=��+	)+c�E�XK�J�YS�H��fQ'��G��Y����'f���T�z�h���vW}���/�ǋe})�vR!~l�6�%!�����ǁ~�l��\��<uB�_<��~���9�5�C�������9��z�_�Eʻ�Fק�8vQ6�o�����6,P���϶v�E�6��3�A�����g����a<���g8;�Q��I�����ư���~��J�#{j�ed����-�U������#�2D4U��1F���ѓ���J�JrBA.�n�@��,�2��ӄn
�������\b<��t��ܱ��PN�)�|���l�%������"�v�]L!�\�^7�ܴY�҄`g5�x?J�ޔ�Q8Y�k�v��P��Jm^	��&�ԟ=�2�䧦�%���֟�
��B���:�ج��j���B�5���������9߂g=���$�с�#гe�3 R+�n(ҽ�r��@$W�ٳ�{�jj�X����<"z��{D��6�@�.d��d�.����!N\\y�4�����S�п�ɒ��3�Ex�&7�0<�xQ�	+�CN�%l�z���6�;#w�j���Z���~���z	 �_���e1d1{}|0^ڞ��IC�A�uR}{#�`&")�A�d˹���=x��� C���rA���Ǯ,%�(�ԟ��u�pz�?��1�8%T�A��l�p������,�1e6�����r�C��zl_�����Y��)Dvzx:|��:����L̳o�a~�Gb�!-�~ڙ�ˑ�Ѡ:�:\RׄO9�����Ф'��O�ÁB���#q
�ڡ����ۿ$)R|��Sk:���H4�����&���!7�C*<{�{��I8��E� �e{s��|HFaB_D�a��3![�x?���G�r�i�7�͡��J-b�ܑ���o,�S���-G��D����� �6�3����BQ��t���vt��}3��*����oZ�?��iÕ�ʢ	l�F����	����n�v|R�n��pÜ����!)�Es��X���y\�%h��s� �64h�OX7:=d}6P@B*�B`0����>��~��;�2*v�*>�6N��`������햝[,z���S5�V�I;i�^=,%�6�w� �&����Ss�#8Ԃ��
�{#��WLz��u��\���2|E�JO�N5�Yf���M-��m�P;0�t2E����2в�W��Gw��mt�#ռ�����z�_��mE�L�ya�����##�!��� ����: $�8�V�ϛ$�j:x}�
�����8���������^��y��������C/�bNx��V\��䏾v�5�I�8��.Pm@pL$k�e�ҪnI/����-�l��~	b�o�~��$��R�q\�d��Z��21��)"�s�e��o��z�9{8��25|5�ɽ�R	S^������W�p�B�=ȫ�UǇ�����ن25mD(�U� >E����RPr�O�I~ֱU��UU/� �]�@���Bݿ�<�uq�l��j����d*9M�f��l��#i?z��Ha$�����ȱv�Փ���������b�	r�^�)��
��x<�}��qK�*�9���:$q�{w^<�ٮ'I��:�k���@۷����>3u�]��;,��X��7w���y�����ņ����1�w��P!E�#��"s՝IpT�]Rgr�,[�����
Xv��,#R�/W�F8wv���	󺰎����N��Z���.�Qf�����O���vCm�˪v# ��������:g��e��"�&$�l��������B��5DI֬S+�,�e���D@�[��aN�!\�z����ƅ�XI�f*��@��&'�����
��;�o���"K��@l>�ő� �KG���[xf��vPd%<8�\m(�}���A	 �W����?"t���4�~�;s�0��vt��0$�F�A�X�.�7�}�߰��wG^�+�5僺Z;���UJ��1�:׳%I*¨]�۾�~h[�n��S���Ј�p�H��c��;��`�<�Z����j�������8ʅL�Js�n��e7�+{��d)b����s�k��b�ɭ��Lԅ��2���D�`�V�GVT6�f=�n�T��ث#�@p��ܟ/��/Uw;kTYc��Wk�d��$y��1��x9�/�"�W>_<�?�xpI�Y��gc��@a~H�u�$y�P�K�[r�z���re�6Sn@��[��R�d�k��
�`�D�M����N�h;�	+������ǡي|ĥ�I�'���ػӓ�"����6B�1�)~��Sе�$��$���.>�t���J!�l�x�Z��6�D��OI�E���~������h���z~���T�87�p�{W���k3"U�)G̖��r���@��BL��}�'��44nO��@�C/�� i�V)'*$�L�I��l0t�pw
q��z}h�����$2ѐ�=L�29
<�R��1ݨ���n�[��+$� �y�O�R�-A�;�54�vm�D��W��{bW�ϖT-�璡ROl�^6���Eh�v��܃�x�Q �S�yN�Q��r�G�ڗ�*��|$�>M%����\!Em�L��Y�y��O�|�%$����7�y-�kzpE>�T΄i��*��ȱęg�rT��̊v�ହ+��ዛ=�1���E���>C��az�ON��{r���f:�i43Wx���nx�����7�����ߡ�B|L�Ⱦ?j23H$.���	5�%�^�T�����K��C�Z�4ğ`�:��j���-�'2�̹����nxZ�n���%�ɔ	ǰ3`�c%4w�;erˡ��p7��{m�c�x�I^�������c�*Aq��Ts��±_8�}PiFn���ҕ)�{��l���=�$���ń�\&1ٞ��֊M��������	�	�"��3�E��J�����;�{�O<!(@7�E���dϽ�����d�Ql�
j�W�RL_wz_q�"Fn�d�_P�Ո���R+�8hg7��y)5���SR��&$}�Ŏ�����=&׬�W�[<ǲč���mz��k��X����� �*�����9�2�䝕�����$(� sW��n�\�gskFtp�q����'H��8�\]��Nb¨�:ҥp;w�EBp�ش~�I���]��(��/�Qa��.k`���*��iOz�G�0ә�Fh�+�6��.�G���i���RS�W�\_u*)���f����6Ю6��e�Q�,I�z
܌�.�C�Rl�%�<��y"��{`'�^5��E�p;�GƦF~ЛLS�bL���n}��yV,�|$[�p=��Pv�S�8����C,{�$u9ZZ!�g��g��4y�k~	 \K�#���{b���sMZd�+�������K�%]�(Xց��r�^WE��J@�_A�ݽ�О�S��d��'[��'��َ9�����Ԡ������7K,��!Bʉ,1D�������s(��z�NLW� ���ww8=`�����ۆ��f�O�D��|�� �Z��n[��7�u֯@��v�IE+n̢Dy�ͤ;Ë�Ix�e��BM;*�4���h�W	R��8S�:�-3%��Q|x:�R4`�<͎i���ћ_�O{� ���s8�� [�'�JaG�êM�>�SS|�Ծ�_ا�
�vK�b��	��N�m�
;E?���?o�p�����g�L�0�j���~][%��?G-~�g-�:Ï��!	k- �Ǌ�]�����o��8�j�e*mv�U�c� a:�����9�+���"@,�/���Z��ϔ���?��|6�V�n,C�bPC����)UI��f�y.�2�3:���aCm� [6R�nA��U
�ּ}�jXi3Y�%dd������E��6�/��-�h���ڣ{��e��y���]#Bc.�.��bUӊ�j�#�|�)q�m���v�y���lqc�Ӄ��+�=���aa����_�%QoQ�]o��d��G-q����G�z�f"g�v�>�9�uBi���e�ʓq�G�-��s�4,wln�D�(f̹�k�֞�ڟ��f�z��v>`�����bZ%>W{>���o>��+��y;!:�pi�H��ӥ��%���A���E��!�6����]���G�3੭W��xi�.J��OCXxZu��78�ϵAU�!�Y�����J�Ӹ��P��/
K�;��0��$���_�?�`h���Cc`��Bhq�����4 �ޘ���o�@�������I�'�RY��pP���Y(�����;`t�j���T�8\���_g�V�n{�j��x�;�y��t���j3�ѐ���f^\bZj�*oś��R��o6uE_I"]�6�����[o�	IU�i���]�݁~�e�D�%Ξg!x�^��C>!r�}���8䥱�Af�!	��hՆ�:�U��AA�"�{���M���Ҫe�ت�"����j��
w�m�־k��N���t�5$#�j�K��~I0�\l;�G��6�5�� f* �Xp��:���/^�⧜6���W� ~;��7�����3np�Z~�c=N��u������b
>��Ow�Z'��ݨ�J ��(���]�2@�b���Ô̿QsE�ɽ����=}��� '�6��n	�=;��i�x��B8�Ū�@���]��#��hɖ��Vl�e�gw֚p4�E�0#�ŉ��W�t���(���4^PG@e4�T'�ܱ ��5Vv�랒��D���'`[� ���[��l�H�*��{~9@'��C�I.�d�T~�NBot��e��8:�g�w���ݽ�j��C6��i�]�=/|�+B3��!�O�o��ؓT[�]1EhT�:��%)lV��K�)a�(�YNʇ���1tn�_���m^�"#%�-K�%�N���(�E��~�#��)XLCX�"�(�8q�%�,�a|�Ce|:�>j�R���%�����7���e�;�ߩ�%v��W��jTg� {���@�U#aQX��LO�7TGG������%�5]& 'Obۑ���}>�Dv�Kpu!�Y:1�Q�"���\,-OSq�b��q��"���FYă�Z~;졽'���>
�0υ�e��C�����dT}2д�Wߴ*E���X-Z�������2����t��e�y��Lո��Ȋm�0�:u��߰�.T�ND��������F�Fm��㹩P��,��v"mˀ�z^�4�o�{J�E�9,��^�ct�TJP��4�8��ԛ�T���˧��,��N[TVU��(d8=�G���q�C	F��΁Ӏ��
�hE�	�
���Ӳ]�KW9��N�������]<�P!6J�O���͎��1��rCM��|S4��˼��������ޮ���@oR��-��'�o{m��v��Z���p78;gř}�nr���M�#�U=��M}x}ƭ�	w6�Z]Jٰ�:`�jPI	�h���k����♟���c}�AG�B�O�*qzj�NL�| �CwV6(�$��?��h�+����J=57�t���d�/���t��1G��%��m/2�T��[��4���M2�>G��Η����{���Vv��������y����[�o@��1�q#>ǽ1[.WUЛ�[AK�6�Շwb&,(�]�G5��4�@kxV��_����y2������7^�:���@�@��w5��j���5�^hkZ�6	Z?�N��+<EXS��d��,��~���m`��	>���F��m�K:�D���Ą�h��z���I)��V7�=YV�G`�~�K���
���p�9�6W��Pp�w�/�~�U�ɜ�Y�',�=�TlC��f����-������2:d���s�1=��j��6��GG�$�J���5�_�ޙ.���o/�e��x(�ch�����l|s���Dh!�L_��ǫy
k�ߊɡ>Yx��ڃ_P�ջ�p�����e/X�@�|�f��	�oh�&�{��K�u���F3�F��]�0���&-�%I���R7�`�7���c7���q�N������ �����R�4�)��Ŷ�i�S�Gjy�B�B�{g#Z�0:wϑ�g�dDL��+��3���Ee�e�$I�1Y��6jج����=8,�z����)4@D�Cq[����W5펣1�n�W�A���M����>��R�?{�2l�ί<jj�#�����f�p{���i 5)!���U��t��=�ra44$�g�����*������֖�q�v���v$�b(ko���䐺�_u�t}������q�?A���)��$�L��ϐ�s��afW��0�I�P�d�E`VW3�j�ֿ��ŬY��1�%�%n�d/����t��|Ά�W>N
u,�#[�(��M{CaF�ſ�R��0-�E�!�X�E��3C�qi\�%7���k�����.}'2�9�o`��"$0�׻;ʊ����Y��dT�W콾�"�f`a�����岑C��ϼ���� ��q��HA�8���D�i߻0�������f�ם��E'w��ѭk�$����y�VV{��l�J�O�&[Q���l�W���@��yե��^$X�j�ښ���vt�&(�������A[u����r��{(���*���	�oN�IIa�YA��u5%!MXa��vO�D�,M#손����|�),�N����fWK���gQ�̪��&����Bg�vp\�M6��������yH�'���������0T?��H� `���CF2O�|���	S��72�;�p�fܘ*��;��,s@�k��'j^�	��%�[F7ʐl8�@�+ф`��0I �[�I��9`U��K#�%����/w��L���E�����Bߠ_w���(��	��,;:�O�
�.�B�%���*y�����UW%Vt��>_l[�GVs)�㺳�3�g}Z�[�-G��\�u�)�� ���� �l8ȸW12kA�a�`�X3�E�~k��M�_	��-+�:�*iԍ����H�	|ժ��%+0�.+���J�;�]�{+Թ�����_O�&Л�$�'wҎ�cnT��>�s��NNF��H�����i�?:ɢ$�͏Y�X�2\�%�W�u��-=��,p�&B/�{��~�&�e+�S,�$����ߐ�i	��(M�BU:4#�1 ��=��������O��WS%v<�gn���������u��p��	�t�\�$�P�\���^9b	5X(�r8⬠�8�S��g����͓�E��z�,B��+�fy@��R��M�{� zc�h8�:'M%ՍÌ7V�A��֣!��ANd�B�T9����M&q���p�v�#�$����]�ЅMqB���H�bGK,���^�u��	b 0P�A���x�=oC�f� �qpp3XF+��GD�l�y~�Y
q!�tQ��gÃ�VMh���Eh�RQq���ď¹'��t�&���zѮt��Z�E�� �FQUp��w��`���7�mG���n'zf�Q�$:1�15%�<��f�ޭ���S�2�,���+��yZ������{�qZ����*Vt�6�&�D�M?ĬC>8���}D����
FL5�h3冸�^m\����� ތ��^�疽>D�(`~�߹6Ss���j����
x�ީ��P�,����!E :���i���F��z��F4�t�e�7��H�q0.UcA�>����޳��z.eҖ�cFh�!䳉q�5�W�/Л�#�z[��c�J��
b