��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��s������\�Ἡl-�y�f�����f� �ѕ:�nA�kb-q��_���ѹ(4�dê*���7��N2�ɐ��+ٞ�4Y6Mx�ejǴ�y9�����=���D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6��\\�l�����r9s��@'�k~�{�<���y�#���i6`#Ɉh:^[����*`��Z��|���z���N?`q_���ר�Z���FLe���Et *�mk7���-��fP���� A��׾��o��Ӡlv�jj�����#�5!�����Ѿ������Rf��Ȏ�����ٺ�:G^7�A'�8�7��������J���А���W����i�k�d. �58+&s\9��]3z |xkbm�F�GɤD���zSl��x�za{����D2���5!���
_���c���E�;����C�6p�$8�mc	N����[$sq+C�o��:���vc9MR�|Z����;`+~�;"n�ԴQ@]\��R�|�4�ː�бÂ{R��O����)Z��k�&�O��7E�yM`>��5�m�"�^63�}�����8A��
+<�%��M�g)�G`:2�[c�Dw)x��y�'� �����m�v��DI����O鈩�0���R�5@��t��㒦�9��o!@& ����v�W���s��mnS��j5�Ѣ��lѓѱȦ��-H������t�	�&�k�M���4�!��X��#�x��V�p�$��ɠmsܓ
Y�A��\RS��H�
��}{s�~8�`��_b�f 1�a��9�E��pi����x|�&��A�8����:]B9/铪DpRqSxt��g˙��t�"*W�\���+��:�Ac�$��Lt����>k&kX���4>>:��+E�)%:���Dr��I������
h�7�U�-[?��Q�L���{� �,���12�(Йʌ��~k�J�����j������`�Ȧ�um�J,(l��ãM)�ׄ^���:PR��;`��2�@�i���7T��鄺5<��*,�q�H*ߎ�HR��I?��AK�t�[�N�d��R�l�v�1U{��X0Bx�g%��=d2ڜ�WLt�b%�r�-e�x�m��zlE�W������?��`ߘBl�	�vw�@�pnn��	%��;�PdGWO�Q3b7����� ����B'�Y�ډAy���&���E��ZX��	�u��UR��u�<m�����.�������dH�5�����[Bl�&�
S~Ch��՝�^"�p�����V<��.ӕkO�����
X����R�����`�����]�ݻ�M�HM
�X�6�i뢚52�2�J��@�cۡ�i�zU�4Eu8�S�� ]�o�������b׋Ao@��ѵ�>� �"#���ǽFe�����e&���$��r2��x���)oxV]Ȅs�"��1!|<�Ͽ�iE����D�V�p}>�4��P/�"ʮ@���N�$eM-DRʌ�)8!�"�ҖRPH����QB�AY�������9I�Hq��Gbղ�ہVl�4��RV`�׭��-�X�S��6���T�$*^�w"�X'�!�ZwFl)z3�X�@*d	yM%w嗂�٪�I���$��v`�5��gSb���� �T���`P��0���B���ה��]V���fa�=�l�s��{��	���:Ε\}������Ro����DQ\�uP�%;�̏��Ta0r)$QVݣ1���N��M{���*~a�ybF�kZ�p�vb�:E����x�(�ţ�L7�����O0K���s�g)�3cV1�L��q�!��Ӽ4�i-�N*n�/i$6M�������f��)ѩ\d�)�5;z���۝��x]Z[��p�+��U�>=�Kuq�a�I�3	�U�y�5u�k�Ѽ���{�����f�|�$C�� �~� 3�U��×a���fgO	��	����m���A	�(p�J���l����j�/t��R4�x�?�k�1�G]��h�7��&x\5�˩|`����~�Ւy6@b�n�k�.]�������P�?)�7ho2y�&��� �	��m�b<&��2T��^Dgc��}�5X�y��|.af�eA@�qŊr��5��Yw�]���_�5��Er��>@t�RC"+9P��r��q�7��le�\��8	�e-����P&�o?�}i^(�V�#P[�O��Ѱi��y�t����Q�ǟG��� �_��T:R�S�/C��s[��d������θ��`j���s��L���̬�y �Ϳ�9��*��W��/5j�y;3rKHm;����Z��$�H����DJ�$�,P�J�F%&�ۖhƫ4¾3����|kx2�����LQ�Z�W�T��v~�0�!�C�������07ס�TyW��iR��J M�A^��I��k�B����p�)������9������`y5���9 �ـ2�gd�R-�^�^Η��:�sG<hv��p�a�Ļ�,隸inN�ExOp�	v�M[XE�ޱ3�?.��! A ЭG���wVFޘ����BN7���Ń�d����fTr���p^B�j�N���Z���q:��ٜǣ �!�|���_�ϴ3�}��`F��Sz&�#�m�^
�S �Zu]'I�c���ɔ�d$9�AN�����Z\L6��A0��K'IX�H�O� ʲ�Cj�	�B���ۄ�ǎ\��(H"^A0`ل��46��Q]����b�)���7���f����Z��@:�*˚�� ���xM�T�b�~�ll�P͘Fs����>�%W[�@Ja�!C/c� �Ŝ�F�,�R#B�BΔ��Y��ۧ�T ��1�,ɩK�1o,��}F�u?���Zk)R��ˋ��+�ÅW�-�"��g�����Ȩ�}�?��Z�㩪!?����o���E�Q0���2�'�W�!�f�����I.�Rc���g���e�4�e���%j3�{���g]6�ޮ��$p�� �)�x4�Dv#x^�X<��Q��y&`�J��!"�lJ�@+��b3{�h�E�d��R�9�"'�r}&���Qnz�ݡ�J��5��>�b��B��֪/4(I!�a��ơ��G�Ђ�B)��exx�z��i�<�O��)}��������= �+�Vr�f��INu�x�k����*���>YG6Y��+{D�z1L,S��	rI��Q�,m�I2��۝���}�էm͌��}H�nI�XesCU����̋gѻ��lsm<	y���F=�)�J�%_\����J��C��/���:*(�������`����1��됋��ظIC���s
A:M"��^�I'�̸�DISh!���B<�U�u��������[��@k���� K��pm���<��&�в�t��Ov��#��l<it7�Ț㖗�{��"�t���9"O��Q�`.@��T� �QА�`�N�"k� �ld�#cUP1l���y��9h��R��M�e�%\,�Ir}mɪId�KU,V6\iNP{��g��B]k�i��U9"'R�K���Ĳ�=l��{��.����5ұ�d�1T�u�1)<;�O���5����t��M�}%�?�d���ǚLz .��Y�!cq��I�n��M�RQ�6�(���O�R��Q�പ�F ΉI�t?M��&�:�Ь���Obpz�9��=���e�� ��8�
��sy���U��32��<�O���
�&uI��h�?a�U֩	���f`E���� ?��zӐ5��8XT��7�H��-�a��k�,c4IP_ow��/�����������6	#\�4����>;�L��s��Dh�%�\^��m9�[���W�ks�P�(8_���c���bz����#�hM"���� {�,�1�Q�`�}P���N:3iA#kk�0m^�/>sB$Qs�n���!}AD��<�Jyn�`�F��T	IU%��fQ>NTH����(T��3Mt#ֈ�D��6}�A�Oz�]�۪ˠ�m��R��b�����Br��qJ��HVXP�a£��ָ }iuI`=G���k���)d���4E E��K�։zk����
��ٷ��^
��Q�5�,���$����\g�Aa�r&PL��~2J������)^�&�(9H�/���U*�z�R� s����ƓK=X�S/ߖ�Z�FwK�f�J��Aq��j�9Mr�xf0����,�����ӱl6ck{q׳@T�}j�&Iͺ�n������Od�v7ze�r1ӽ��\#'�_\>5b7�w��[v1�1IN�� �e�z��~(v�c�MOk��@B'�tT�x\~]G;�\Y���4�iDk�L���lk�@[-�L�����S��?�&j�S*�Zk-����(�&s�:��c��
�7Y+��c�(��K��C�g��-�����;�4�ʉ��td02��S~�6h��=���,Of0��P����N+���S��_��w?����2Y ��@���n=�4�GwZ9���M����[�߽`�]�勉���R2gJ�~�xNׇY���݉#��2#��R�I�i�Ḱ~�ΌZ�Ø@.�����9iU1k�>�
�qۖ��I�^s2���H.Q[6�
R�//��!r~�3� ���A�	�l��h8����}�ߒV����q�������9���6���0���3(�.�/�7�p�!���<s��>Z�`���2�pa�@�ٕ�9>f��&��n�Z	�v}��
;S�m��s�����)|��bA<+���)��A	�Ē׏;&'[c�2^�'��촣����v�9Č.+W��3ژ��2���D��ó�8�z}�~�5�5��bZ�\��i���N�[�':Gz����j/�*��v���P^���$���N#,���W+�e�,�n�H�k(=B�q��"����w��3sO. �s��F.�])e��O;���ؚ|� �\QԔ��M��<v�Q4%Z��*21�9���{�ϩ[n�M>v��<\�����(�I kv0i�1�5vd�!�k��ے#��!6%W?s�~I�'>s����$Z�9V۽�F.qv1t���s�J|���oVůW�2P�cPvˋ��#GS�6q�k[Z��[�]ibЍ&�K���Nd~',P�yW��+�;i�-b��R|�6r�I�����pP�k�������z��Ӭ5�Y͸c�Ǯ_'���q��ĻFg�g�Z j�+�2tb�U�F�+�Bӻ�-Y=;�v~,��\�"е��p4���S�X�S�>��/� �+�ϰ�l��4�B��8��!�P̑��`T��0}A�����8��@�Ŵ�=f�����2@, á�tx0>)�O���7�P�����y�*�(��=0���7�YXU�Lj��-}>�7�/n�s`Aa��B�8���-e��!��<��_E.|�N���F`�UJ=����ض�&�����>���Y��}	'�r
P��|f۠��o�H�Z�@�H�5JY!=�;CL�j}g+)��!��QT���S��i�Y75��5��{;�"p�S�Vx����_S[%��wcm�w%�R�C
�m�%ѣ��uV@7���6OQf��[��Ws�cx��K�[��n�b�?=�b�K��b@a��(�����r �����{�w.���� �T���9�^n�@�
�Y�X�)�	��pi�/l�d�yL����5�?�Ϝ��d��@�Mq��(w�<��;���z�;5�SP	mZ����X�d=8����љ����ki`�!8�\�����K^5oϐC-�}�Eto�Kh�����P��8�aRct�!ُ��Gp��V	��P�� .{0�dd�"��=n7jzιֻ]��{R�ˣ7�v�D�5r�� �R���%�;�[(>Bh��:n�$bN&Г����G�����Α�uԤ9Tp2�	V]�e��?���u �^���-�;���f)ů��?n̾�B� �]`����qpg�x�Ky��`!�=��W����#��=
cFu��ԄV��~�Ǥ��~�U	���8��3��)oG�<3j��Qq�;+�Zwl*W�ZL���H|�_Σ�B.�t)\5�;wU��E��6#�|�\��$B��%B�/����GӔ�>/�-L0���9�?��t�ݬ���>
�����{f���	~3��*�����&S3�p7�����8��"�#��5F���}K�츎{��#l]�a�H���+*�L�U�l��IBA�Y�����<�-[u���G�O�9�D�1^W��m8Ȓź�G�$b�[��_���ٵ/�e�z�"\��iE���R$׳ǚK�|�O��o���msH�~-�)`%:��t�?\Eb
��t�����P4�5X��i�gz8 �]
zk�O�t(8Y#3��`�r��.2r��;�HG���j��~@-�@ ��=�g�yf�ӫ{*bs;�r�GV���Dk3e�ow���b�H���)1�$0PW/(����ߤB	V	��ޠ�T2��/P����4L}�*���Ă(���U35o�G`ĢgW6E3��ʾ!{��J�Y�6BI�rݝa��A��5���y�3D�b���6�P�����tJ2��C�W*W9dG/e֌�|D�WK�*M�ĸc��o��K/W�����"G''��p5����0ջKr�N6�"�����֑����#(��G�����RĞ -nd����������FMP��yV�_a���x\ �b_�=��f��-o+>�~���N@򊽚4��u��X�!�yVpa2�u-tWX����"�y!z����`�A��wq�In��*�8y��Ѻ�䣵0�1*%��5�zl�׌0�b�֧R�]_Vd�q�Ĳ�Y�up���q��j�R�MǉZ�K�,�a|�=A�E�*�B|Q���Ӛ�Me��S���Jʇ>��nj�=Pm8'��󪴲
�VJ�FILH�1uzG�/>�����DS���2L᫈��3�+-�������ڕ��e��;f�z�$HӃ^K�d�������TV�҂��w�JL"�����c�3���K�P팇���Ib_
����nVA���O; �G^>C'jHHA�ָK+�^93��҇:��������w�,�T����9�*5/$Q��3;|���0�����/�m(�rw�Y�.���F'۵"�Q��dߣX�G�X`�Dh#�MCt?g�*e�-Wr��8�RE�bRYaB�m`�'�!�� �+r�NV8n̵&�9���8	��s)��`�vwOl��ܠ�sI�uf�u�ql!L!��}���|毸;� bR�ܽ8G$��ó�U�yM+��휍%/��E9�+�L✫���͓w?�Xd�S�]��M��K�<�z�6���՚�`�I�
SFOv��/a	y�"-Z��T&ބ��@�U��~��.��_m�z� C�%"p�wJo�S��o]��ı�������O����~�a �J� Y}���2����HS�?�"ս4c�$��4��߆�����I l:�;몉_�[`���mP��q�J�1��!�W�T3{�M���q���F�I��a2�����*�B�u�C\��i7`^W��u\�N�I��&e��$����4����0��bj�U�-
��I@���'zP���VVds,Q���b*k~�O�������8�I#���+���aӾm(������9J����G������w�sd\�wTYx:��H�v�_~�v$�.�	��ldg&e0�p�-2Ly��P��̓�+�"���+�E��O�����p���� VW՟�L�@����8���kz��c<��D�o4y��S�S5n���#v�H�ԩ��a��5����p�{���:�5���b��q�`��w�)�y>φ�Siڇ�ڳ�j�Y��Փ�n_�+�1�|-�������䎋j���pFI�lD�����կ�=7���$���y[�G���IVB���k�õ��<�)���xj�2>2�}��a���*No�a#hKe[X�i��P��dߴa�GU��-HlL�2���{ܳ*M�hγG�I3}�g kӰ׳Rrs�ݩ��J���.G��ix1����4{C���~�!�xh��"�^��#m�ٷf�hgW�NN�i<��/�p�[����Z�{x䃶�Ae�����0M���4jP=/��Ѳ�/�𞏺q�|�;�j�l�_�|i7�cOZ�<�ݳ�M��Vأ�:-y8��h�I���9�����ɻ|�6�?#9�*����ɋBc|�T�&o�{��㯐�[�*g��@(f<+Qy?��k1�s�U�:B�'�����ߏ�/T�b�$�*E2%��'��pQD(<�(I��2��k��w*FEN�f�'�A�(�R��XK�u(�)�K�H���_��ŀ�O���G��n�x���n� ŏNܬ�k�4��Y>��GQ��&��$ ���5C,�?�;��T��)�Үi�R�/N�7��7�#@��簇��w�Ջ.��\"H���AIFޢ\���wЀL�,#����oX�4�A��l���bL�Q�C}.��{t,���zJ!2�9,�h�I�Q�t�2C������=�j��B�7�`WP���r'��	*���޸�jQ:��x�wm�M#i��.�U+Ύ����V��=��'�m�NU8�s���e��t`jƟ[&IM9r�vwU� ���{it�h�A��X&�Z�R�����PA�jX��G��X�5y��Q�<�t��_�1��{�g��{LxT;��nW	��x��eDYbz Sq!Z���!L�]�\�+D�n���cw �����zca{g��ә:��>�SA��Gsy���c��}��=���G��]�k@@��HFX���:lH�\�nV=�K>�V�[a~�� �$�a�1�_O�H.��a�|��.��|�M���A`��X�C�(d��!9�`-�AAc�cR�pv�g�)W�NR%vv����Ma
q{��g�"�IV�Y�H�UV� ��}���,E������pLI�e���z���\n�i��"���٢�B�]sp�ܓkb)��l\ppA
�xW�y%by���O�lyk������	�C�Y)¹/%uh��5s�p*%���^���հ�	����@`Q�b�$���*b�����N�i{S��7v�_���0�E��3?�yj��ب�ʙq�| Ϻ_�/�	|�D���9�Womm�P!���B�3��ih8��h?߄>Yr?Ν�A9om���P_�ݚ����`�h���W������8�b�W���gK�d7�0ʄh2��a����oB~�[�=�|b�1Ϙr�I�0�(Ҵ-P=R��т��E:90F0�Y�ȼMT�\"hcQ�r\G=�[Ĳ�Ո�轗�ȱ�8�����O�)$�	t���zs�ӿ8Y'�޷�;O'R��3NzZ��X�o;����vw�N��8�䷺mv������?7?�N����2�f !;W���7A�� ���I��^�x�5���u�ӠrR�I�7؉	D��WV����k�7w�nE�B{#�;��^��篺�<$ϨI9�iv�}�n�T(q~�$5��k.�[A�ʧ������w�f� �r�dϸL3Á�VK�#�1�õ�y�g�ʭ�7�2ť���N�t�2���I�@�'��ca���G���#�%p��p��ӗWI2�:���vY5��vtP�]Pն�,t���)F�iK���Q��b7����ɷ�m2����D�5�H3��"��)��V4��X�A��LW��ir�Q�i�_�˾���;�l���hB�M.�4�Ox�c�Y��zD���~.\K��*�̔ ����W��.V��q�#<O��؁��U%D
�_�� 2�dQ�3�b�7T��9cd���Ala�嵠���>=��h�������'nR!յ���ʘ��T������W�s��"/
B.��6׆��ܸ���m��I�=��29s#�2ήom��g�ۗ�l�z;$a!�b,��|z�'��$aʊ�E��1ly1;;OH�Z{/B��N�[#��ǐlL���+`�
_��t��:���{Zi�	�P��fc�$"�Q|�M8nx�p� ���Q�����<X�4�d�@X��e�� ,�zZ'�;��4F�4���3k+�|��huH��6<�B�ǌ=������Ҍ$3üi�L�K��*����oʊ�.�a�O��R�+f)m�F�q@�9�|��:@Ғ3����jBi�����f[@��--�$0�5�[��w�qb�V�g�������L���uj��x&!ݎ&T�$J �7��d�r8���]�����$;������S]��ғ�t������".F��琁�����K釲Mg1M��JR86R^�v�1��Y�do�O���?�(1���dm|����B<i$���~y��0��Gf�W�ֻ���
��,���{<L�'y��%���U:�_����v��W��y�!�/o����t�lضw�~o{��m��8{�j�7M9��B[5�e�^���If�2�����ƽ�7u�t�~�O�1���R�YD@�7a�X�M��H4d_��H0+
A�`/ǎ�`!|dKA��@���������,_��R׾Տ���W������,agHw�-�)��s���u� `���^�Xt­��;���� 6L.������O����\H�S��8�] ���]U�����kcg��=3�U�e[.��4�T{��.ii�ɉ�s��j����Bu���qq:l�.��AG��b�'_�i���2@�-����3����N�x��6�A��0�+�k�a�݄^7��Y/�L�؛�t�;��]�.��·I�/�{?b�t��D���a���>o����K,�NJ�S\����x_d�ĹYV�J�PQ�IL��:A�b�<�^_
�ќ̑YrC;GU��H}�R���D�o��ZG��+^��9�
U��%����'��8��<�������>��t��ZV��JQ��lap�C��}V��
6�/97w3qC�=@��lvO�8t�`�y�9�3�D�B�#<�v�Miڌ{*��֊c��0B\F��)�|��.k$|�1���Њ�HFrΠL�FK��m��˿!1,;�/'3r�hM�3�*�L��e�;����eA�2����"�:�]%�:��UppY�fh�j�j�-_+�|������9����s��tڙ�#9r�3L�46�Q5��_�!�olo���8�c��LO�ʘ�W#f�U�{YK8X�[��v,�cu%?�PE�����~����X~����w���I�,,� �E���mo�fL�q�:�w<游�e��'4M���9�6�n�W��m�;(+��
0 ���<�t��
��lOl���xq�ї��rk:�f���`V6k�Hn���]����d���S�� ���G�e��r3���$�Bt�����<~L��ڀ��
���N���:�Ǵ���-$"2~�^ �~cZ&��<��|��c-/���{��J��Șo�0[����:�A��cj^��+F-�~�ͮ�����bwX� �R%�3�绉5�Nf��㟀���AD���>҇�Ym0�$T�����_��2ԕ	O�cvmf���k��b,�3>��2���R:j$��}A&294�=*k�*��:�}���<�K��[v��d��z�i�-Aa:�㺆�o_��Y����i0�ކ��e��.�]�������,d���Q�`���Ʃ��K��:j��s���Jh��Q�$*;�"�����K��;;�
<*$�%��'�,plQch���������R�,��h�k���Ɛ�1������t�ȼ�{������Oe9i<���>�Q� -x��O����u�øW�69�y'����3���q_����<���~s�&�9C�b�	�1W<�$c�5��B� <^pR��u`�S����bZ�"Y�I���qCT��L�HA�3���Hi�H�\>_F
�y�:ff���0D2��ŀn���\��y�R�c�G��:H�㏛?���5���^��#Dir�	��і�>$qȘn��(�I2R$G��b ���E�F��Vn��;ɛ��4�,[BH1$X���S1�>�fB��k��M�u�(��$���㚺r3x�O%rg�����e̦;ʜ�j��dm�}iӓ�Dn���n�[I�N念��W��2Z�kJ$���ǋIw!��� �ww���`��h㔾xp����W�}[Ļ"�6���~ti)^��>��0s�ڀ�Sh�#��w������2������P��<i{7o�C]§��Ǿ�ұyaK�~�,,�����V��!��c8F�`����ėG3��U ����a��ǆ|��'��J�R5�4ݯ-�<K�-��Œ�:��`����/�"��(�~�pQ��@;=<%qf�w&϶stK�u.m�3���0���k��s���_� Ѹ.$/��}(��c�D�>܃pO��i�C��M�6H��[�/���ңQ��O�,�+>���tNv�bNp�5��Z�7PGI����bm��a@��K��4:�H��&	FB������р�(D����>ؼ�h��6��Sת[ X,�����#��ԧl���iڱ:::�`�`�f%�.��{������6�&�#҃YGk]�+С�Y{�o�\���$��i)w��CC��P*��'��(]�3�]��6	�x���Ƣ�+N�B�����~���ʻ���Oi<^!㣥�"�0%n^yW
��o�n�ӝ�E1R����IJ h�$���t�3���D�	�)3ʶ�|6�uF=�EѭG[��*w�����A��5�1Q� ��;UO?������,�>��W�d�ֳ���0){����\��X�E������!�<}�f��t��*��zS�)A�V8���ϥ1��_�t�<aW�d&�$B5f�U�=�m\�����+���S��@�nB6��a�q��[�[6+�;�sfT(:��3	����4�{�{+��04o`Z���LtD¨^�r�h�6���ǳ����޸0!�ɋ�J���yA�X3W�'��o�{�bU���w���ٝ̀d�n�soǵ<݉�0o�44_,�A�t�x�<!'�����s� I��X�dV�->�NF����1�LꌙզW���َ.I�ռ���q��n�븛�<����Z-��$(�����~��b��_5�'�ҟ���m�Tdx��� �.���Z��V����ča���Y�����߈����N�q>�n��m�3�_p_�lI,�F���G$��m0|�v5�-�!(۷&kV�FB���:6�GP������fJ�����A��[�%l����j��Ha���k�'�c�^��m��3�n)Օ_�r��Q@�6�"��m���>�����E2�>�5h��N���	e8�����3뼥�	p�LB�aX���%�uJ�P�|����,;��~2��8v�׽��7lh�R�}l'F���v�`��
�q䔔:Y*=�說M<���ݙJ&�1��$��������iS���>z��C��B�y�_M>�ty��HI��	���f��@Kuܟ�j��FX�r�蜎ީ����	�t!U	7yT���\~���[�9RR�۰�Ď��P��r��ОB�X���=�aηy��>)�b��<�d��F�?�Y�����/���[�t����*\iA�� P*�#+�����[�&V m�����>)�b�$�Ο�F�2�����f�2����ӝ�V��y�u|+�L${Re��~w��'��iE�MUUq�n�A��W��r�Hc����@ﮘ�ܘ(ַ�;�{8O������X�3�i$ab�@UN�f���$��N''��M=;5�Sw�/��U<�.S1�4ճ���dk&c2_0@�9*]B:~��I�� �S|�^)6Ў/�6c�����_P�\�y��_���K{6x^�R��=��O.�
���A�~U���E�-��.J��8r���O'7��o%�Bz9;)�f����7*]Ԫ�[��45( ;���V�>�6Fɬvg챩6��^��<軌�A�z�lBh��1ua�&+v"�*�/��X�Dz��]�� �:SM����x~�[g��{I川�9w@��o����	u^���U
��OM?Z4S���V[�e+>�s8�F��Y�v��S3�t�=�(�鮦*�)p��֢�}М�s�0|(`Ĭ�qm�!|Y��6�n1�c��V����W���-4G�R�P�j�ԃ#�@Nt�Q9H>GP�`�,㜯A�&pZ�b�z_��"-�PϠn&Ƶ�ر0Νf�r�Z��":�\�5��s\��M����� ����~�[j�Zw�ZYIӣ0���v��_��a�/ �T)�t�w`+H�8��H#מ:�'��!�Vu����w�l8/0l�M��������a-�"�_M0��Ū�*$䟯w�^��������#+��O���\�aN ����Z��h�d��jg
X��c6����(��*�����EB�Lh��>
��X\����g�{����!/o�MeT�f�m�{3,s�'�� Y��v�H�����+��&7��=z��ǼwX}0%ɨ@`sUVJV�k�j��y?��+l�X��_J�j�9�*{�m�i���c��_�y��zKsh��
�`��t;H�Or��F��VG_����mC���NT�!�ɘsm�����~m,��~��-�S
�A����Jc�y-���qOW�,���,����	!�P�3�i���C��?�Ni�қ4��*^��T�%�V��u r��:�1W�[��[��ۊ���}��;IRԮ�V �~Iu/�����(wU9�$��q�j��X#K��Lڀ��"����4���2r�=g/qE�|/�e���F�6��u�����l�d����_��\҅�f� ,�)X{x��.J��Π�c��M3|]��f��o��x�w�1/=��tQ����j�+�ݦk���Nm]���XԪ�#iAI��;}K�\۹���>v-V5�	5O
��i�U��'% )\��U@�X���iֈ���rH#��em(e����;p}���(�9Er{IG�8y����}+�V�Y*A�3�a�LY����F�c&��3�[�y�\��8;zT��=�W	���|�?D��0���Q��/�{�E,vf��R6$J�Α�K�0z˳g!�)p(�L#�[N^���
oϟ�7�b�5��B���+g��4�+cɀ��Eʎ(1ۜ ^�$E��a_��S��/�8�Z n(ܞ���~������/?�yD��t���|H�M4c�P�bc���@tѨp��6�v��ub�`�Szw-I��ԩ�C|5ln�����-�10�bJs�i:�٤�9v?��@���X�.��_�u2F�pY��Nx�ޢ���D��$��ü7����Y�Oؕx�A�@grs�2�E������m�c{�̰����VYL�!Tm1���I�r� 9�07LU� ��p���3�;)���R��2g��/�=_=�y͙y`��ad�r��"ԍ�1˿Հ*�YI���br��u��.��X�5��g���r�I�#%�CY¡�}�x���s��3.���D�q�\I��R�f� ��Û�ȝ�k.�o{�h]Ð'vĻ��PEC0Gy��-5��/����e���*��V�/�H�w�;�)"c����������6�Z��g ��L��(�f��z���!�6����q;A�x�h�C�{�@�)�۹c�)����bh�s"'��ϒ9�����׆��m�>�u]�&�Ͻ�.7��И���9b:��tiLq�
s��OC�$�~P����I=�8FfEں\T�`�-�P}�k��<'�p��P.*��+ɫG? Z�(->�#�Nlr@>�2/�wg��tB$���ʥ6�F�UJ�@�پmW�CjMT.���s;D��^s����Y���u�+%m�i>�^Qm>�@1��i�F��
�2�o$��w�G��k���H.��0=�Yԩ��Y�N�_ �
TF�Q�6�lZP��J�8���� qς�k�Vq�q�=:e0�QGWG��߯B�����0bjpN���5L0�vMT�^�����Ǝ��磿T��-�Ɵ�/x�結�t�r<(:`�@�ˡ1e���ƍ�P���p22( Ǟ���є-���^���Hc1�`���'�ț
 �x�]���~�I�[^��إ���͊Qxr�lus`�T_�(I�r�QB���<�.�ӅT	(էp�Ko�L���[�*����d�p���!��t*a4f�K����.ħ�DæH*4(�Y�Na+b%kV��P|t� 7D�l(Iഃv�SP��N�<��$a�r(�.2nS�4n���f�F���Z�����������mB5tE��jIY�l�E�[��; تX�>VF&{{��ė���"��;J����&	rj�0	�j=���o�Ζ��n9����Ñ���ڐ��R�1�c%@�>��T�Qhj&�37)-F��8 k;7[L-�3�%��X��c�b�$A�!W	�����~�CWʔ�\̋]�]�h$�L~XSe�"�%}�ϛ�V�?�/�S����>�>8�{v�.^�0%!3���t`�7�CmtGE|�c��튭3�l5������o ���3����|����tOs�B�oǱ-�����9�j�Ni?�$U�%�������].a	�9 Q��n�D��#��t_�^��\h[�wy����k�����VL�9�p��w1�\�뗭����f�Hj쭉K�����뗧����f;��ܼ�k�o�.
�@Ђl^�O�25�i�����`7���_l�jv�����̳��T�yzO�I6�\�\(A=0�⨉� ������aR�`����BR�k$�5���n�G�����ac�ItJ�ۧ�I��;��?���_	�����x�^�2ꟵlM�3���}����cG�`�<�dg���M�R�I��,;w�N.N'U~�wN���S��b��Bǩ�;��,�4�S ^�*;�~��޴a*]$v�>�_�1O��/��F���+��}M_�p̓��O������]<�L��4�L0>��B��n�T!��-�|����w��AB	7�c�=ԐF_���.z��r�$}�����z���A�V���*�����<��!#Q×�)0�(�td��W6�a¯��sn�=],���=���s%D��e�5HcC)n�K�]�w��=�4dRs
�;ޜ�$�y
{p?����� ł��唤)���>�"��=(յm����;�W�8�.@*�Iˆ+����e�.��/��������G��V�:0��-#�|����ث�VI���;��\��bD�Us��������p2Z���|&V�h�'5�s���Kl���߀؝zS�r�Y����J���2au��[���#6�!-Au�ӑS5X	��u��?��$`a�88�f�h3�	K�����̾����3V��2#������$\
x8�C�i�Kz���&� `,K��$�(���>�hI�U=F�?��|j�q��x�/X��"C���fT�n`�-�K6Ko�G9 ��/�Tb;�ҏP^O� �Y�F�5֙E�*"F�dv I�)��S`�C�ŧK��E��/;�[��m��D�ٍc��O���v'� ���\.7�,fv������@����a#�	��h^Eq/<��r"���؋#W>���Χ�6��~�[����e��C�e���͛bm��ͥq��o��
�/��D]XdhS��Ri:+Q�5�� �M�AƮ�;�LU߸�T#�u@����م��dU��ʙ����W��Y��
yy}��ٴv�ٟ[������#��,�ജ3'ygsu���JOB�l���#⒚�]�9��c�q~� ��3�F8����Zk�d��uBfɏI)�5_�%��*jC�6ubi�<��w����#	D̿Yd�f��h�t7a2�����!Z ؼ� ��Sn�"����<���6%mrg]#�o�nZsh�"���t�+Z������9��7j2�^���A�Ȱ�����Ϻ�F"�՘Z�,�?x�%�k	Q�Ұ>�?�c7~�a 	4l��je
�~ܵfH��\� ��=XH���9 |[!�F����1���9ts^�m�3� ,�%���@*(�f��6�������$�N�.N�xaZ��}CY慗>�hYٕ !�O�ޅFxM�b��،T���ˮʑ�[�k�x�Մg�c}��)o*�QR�r�u
(��S��/4Yږw�F�-߬T9�p-	�s0�#�|iں�!�����/���<����
�.D�U]yt�YP�tlܕ�Q:�s;
�w`��)Ӊ1�R�������M���1<�k����&���c���'IQO���XsJ��ҙ�:=��O> �w��?7ѣ����A@ǋoj��ځI��X[;�I/cF~?Vo�Eڜ���&��m�ީhzq�B�@{M��l)����7�)P۶���<ߺ��!��3��Ab�.�>]ͣ���'|¥jF��<�z�ˑ���dd]�;N�BGHg\���ZY3�(^8W����g]Z��-�"AE�%)��,���f�r�`(����F������:	��.����Y��g��"�Nu���J>�ؕ^=��KW��6,x����y�q��߃e�!��Dt�`�}����K>}8��D��Y�D�6��F���_ʱ5g�/}��?{�4{���؍�k�hs���)��|;�@�V��s��ZeiK��l�%� �w��g��3�}�#�Qt�ވ!�G*М>���ݒ�1[}���0��U�$՛/
���È��j�JjnO�!9|�r�7ަ��rB�����a-���A|�a'Av**�r]בp��F��!��"A��kc�#��T�^� ;`8H�=aM�B�@f�]h���u�8#$��iOɀA�%blGi4�}��B��Uuj���rrq��yw�Z�Vn������ELl��$���.	jI��@��,�^��J�Ò�l�w�����hZs�Ԟ�/�ZBYC<�.��n��	�m��zu�+t��r11�S�JǓs�
������^�5չ�	��w�Ye�:I����S'���@�G��ʀ���{W�K¢���"Rvmsރ�  m�-Q�F���<�+gf�l\y�edJ�r�b����7C���ZE�uDDp(Z��N�H��p�X`Y#�gl\r�~��6k�]�F�ZAsʝ<�x���"{_ے��!��	����s.��M_�#{K�	;]J�tH�'�T]��p�re7�J\~t�B?�s�`�$)g�F��ćs�4��[Z_��=�;��k5�Z��lβt�|x�y����eMϚW�-����Ʒ��I~g�9��ޣZ�\5,�&����elC��#�(=�߆;Q���o���+s���ژ�7��h]���,U�b��Xh� ��W�&���ٞ��dx�=U�U��q�bP>��$FQW����yXtt�b�1�2@�oH�	��lt��26@�~�@�k�g,:�����(��O�����@x(*���T������ap0�p%�a�6��p�u�t�*�Q�[�m�GJ�;j��Y�߱���ޅ�����Q:w���d�A�ѳ6����mI���6M�X�]VwNi�]R����NpW½�xs�}�͈C0���M�kρ�;��p>��m�L�g9����I��N���&�4����1g'��Z�s^�sh ��l�A3Ή=�,W�L�\ߪ��s˫A�kX�}���T��q����$�-�t1� �Gz�l*���Jߍ�Gt�9�R�Y��	P�2�*�c�H�XoQ��������x�]�Ȫ���i_�at�x�:�ߕ��F]�t���L�����/`���3z�,P?���{��;4�`�}�Xi��L[�$K�![�N�,��y4n�/V7�d�ض ao��s��<Y9�>ݛ��8]L�ѓTo,i
>g�v��޴k��RĞ�JXC��2�IĿe<��˽c�a�uV���4��p�6pY5�1m����� (��9֒�৏�a0 �P��.N���;Y�\T�mY���r���>=�ܹ�^��+�5�Xw.���V��$��^"H/��ҋ�r�� ̻�eEèf���e�Tj$�:vV5��D��=#��8Ax-�`�^F�p��W���F�5��4E���j!ʞ���5�-�{���9�7��a���|���/�%���:p��J�L�?"�ݤ�U���
]�y&>�ċJ{tt����f~r����H�<ӗ5�^4�7�����m
<˼F��R��4�,H����'%�i�t�"&zM��~�0�Hy��#I�&D��=��g�Zt�Ճ㱕0w2��H|���~v�v�!M�$�T�R8�B��Kq�+٠�`Yz�BR��y�2y��yJ/��#G��]��e�)&U�Qꬊ����Y���e���|�O<�4���Nq,ͫg���Զ�^�6:?��}��1���%i�o�я��1�J���;��CA�ˎ���T�BAIi���;��ln�
jkV9Ȅ2���%�㪗�o��1�z������ ��=�xO.1�����HK��c�s��o����/�V����=o��=泹h��*'T�<�غ��c3�H)')B���g���4��;��-��i���f��Nϫ�B}��j�/��8��e�:H����:����(�,dP[�Y#�Rq����h�̽���;���H5>���
W"	��zbR��W���,�9v�YW�h*3Y�_c�=���/m�[���{}�0r$���i�йB�(]�Sz��d�p�y���'��opos�j��PԮ�a�e����&ױ�.��(��������^E�-k�	������k�q��T���Gkz�A�f�R���
(:J��v���b���KaR�w#��k=�B�A t�#�Qt{$=R�_%��ɝK����$Y3��~�0T�s�YxX��s+�E+�z'7]?ӄFn��߀M~���;�w^O�p;w����+��^l%�_H!l�-p��(+%4�~]oNʘڮ0�L���.�=�m���m��I�f��O���V�u")<`�G!R.zB׈:\A)�A�yS,��k󪺽�%��,�4�����/_���F�9�����Wx2mմ^n�����WD��W����Y?R,�oq=N�{�������EĲB��j���I�_�T&*t]x���hY����`���R0������l(��O�R����B"���w�)^��&�Sa��v�f�dQ��3\uX(��-M�o{��ӇAB9�����M�a���ue�Z�o����o���#)��P��y<���ħ�4}�څ?4��#]��B�o��t,~p:� ����m`�q��A�^�X3
ߏI
J�92�r������ ��;(�c����k���(�����؎Z�|s��qzΜ��ܠ܊�h.Z�Y+֭�Gz�6��*�'�Cq1�����3�5SшQ��W7�eg��&:�����>�YO�w Q�[��/�G�
�+�H�������;��&��S���[������Do�1��O�w7ň�Q DCR�V�í�f���7��` K��uCʱ�־�ݹ߷�r�̠�ѳD��I��m��h/�;��,#@j�(~�>Ui,m�"�"Gwb�><Jܛ�\��bڗkrk&*��)�]�.]���
�2�w��5K�z��A��G�����C�*$�.=	:�*�I� 5c��5p�l[���r�}�5����+|ƤF�{��7�v)M��k��\��I9�|�~
���a�
u� ��H�����޶������HHn���h'��))>%׻�=��O7��5MV�iƺ����݁�4�H�P��:1�%y�l�<�:<����V�NWVZ;����^{u��A��c��|��P�b�����s�؆����.��|?��M?5&Ә?|l���p�_Mm��3��绖ҹl�a,b#X�K�(��,��W�F���Iy�Y�9ow-W���"|Y�Ƹ��1*�Ґ���S�A�)�Ύ�]�� ���z�XҼ�����PAХˊX^�����"���5l�
���I��}`-K�\k���`�`�.�x(��Q��%�j˒}Cy$��l�h|=�:f\*ǜOok>�ԭ�jS{��	�N��=����A��%�E`s�&�3�90�l��\T�v2i�Nl��F���Z�����PbEG}�ج�Zs��J���s.�D������!j���+{���,���ʌ ʍ��TRA�ξeY�;7d�I�M����,��5�X��$��(@���W�N��bb���
oԆQ���9ssm#��� �5=9]vjA}��i=8�r�f�_&t��Ni@ �^(����b�?�b.�o�X�� �6��R�A�����-�E��!䏏�H��ǈ���zU�3~<�n+RtԐ���������3��*̓9�d�#����ꩅ�>I<�.z8#��[�����C΁Σ�Wπ�{��!�U����D� �����S�Ә�>_��U!��oH�{���b�wX3�l�vYg���'�,���#|�]|��펻2r�J�e�%wK^����;D�1N�ubڜ��i2�Z�#��8=�v�Ӌ�,��,�C�9Z��?�f��]������d1�1�x�T�x�0{�j���'�KX��lB�G�:U޶-�k�r~%E܋xt��ľ�xT��MlhJ�9���ee���ltD�]��6����L(Ovo���J�-�'� cE6�@���7�K������yg��YV]�,d|_����8�$s?�Tݏ��Uwo��%��ڏ� SÛ�Y��*n\�40T��h������t��,(M�ثv�=�G>P͌q7�A�wd����yg���bm������e��{�Q���`� �.���J�9j�.V�jn���%9�0�EK���B���bݙ$9w�1�^�=���M�%]�%�a�$��f�S���6#||���
y�+���0ɢ�	�w��<U��o�0J�]Şò�6lrf��ʨ$r�j��N����l͊4p/7pTK��`��:Q����q���sR�&o�����������u^6���Q�!��ףt'f����zN���Qq�B�L?�{��DG� �6����Y��d���Za���%{T�"�e���ؑp��ڒ�l5�LV��3���%���K�}��A�nng;.ز�9Ep~%B��~U�W�{�s)^�E�	g4�y� G��D��*A�ثSi�n�>6�-e�)��d�[�W��˽2��^]qĎ�����5B�[�+ �FIj����W��Ô�weM���<���U奊Xʾ���,&M��|��>���b��Y��~^����tOm�f2Qnv���пN�Cv>c�k����V�b�0�֏��8}��ӟx=�k��3�	R����b7'98�g�<fm�D�d[~�8r�j�J����ш�bI�w�5��F��R<��o�pQ����/K����[ �.�y�=�c�~�#t4�3�tP�B�b�[�;JcfcݑA��J�v�4�3�#�/x�zS�vN>ǁ�N��h�M����/DZ	���0�0kUs+���[]�f�o�Xl3XG��M)��3gw�����2���`����k�/�0j�Y�f.�m3Y@V)U�*G�d�>z���3%KJ�ͩ���.��Fnj/v�IC �}�x+J��;�V��8�^|3�3�g�x!e����l?$9q[�E������0����tD�ѩ�T}wkx��x$�ٵ�h�$.��I����7��r' �߻iF��.�vOf�.���08zT��I��ٿ�g��2g��jd[��b�"[+T8��q���a.�7g_�PfOI�C�)�����#���Շ�������Zξ�뽓�q��I�����G�z��q�W���f�c�	ZS�ٷPʵ��\=�*��;m�`k��t����c�p��u9���ٴ+��J��8�Y���FpU�N'yv/v�h�<k�`f;L�T����\
4,���܊]P��і�) �����3�W�-��I��q�8s3��@rP��V恮z����� ���A��~D��C�[�l���Գl�)����#?��n~�ՠx�up���r� �<gpB�I��6c0��ϕ+����q=1	�N�U�:תë�.�Ӱq':*I7�khqL^K������Oc��<�)e�a��ϓ�L��P�FA[��z��6��S�b��Y�1�.+���k`��:=�6���i?���	L����tV����	{�S�hf���$Òxv&j~���!�h ��c�M~���wz�����ޗ,�k%�'���1�*��Go��̱$}Z+k3�v���p��(�4<�e�f'M�K�kE�Lc�<�QM!s�a1@�~m؍E�{sz���x5�b�C%���ϣ����KQ��b}����1���&�B�Yt��j�l�@��S��nZE�4��#�ʻj�zx�\��lZ��fLx��9SnV�ܨʬ
�|��g<a8��o�z i�2 E�E���:C�`�f�d��(�a�	���UI�g }�^�i=Yt~"@�q����5F�)�6���)�
	��w�~�Lm�Ikp3��>h�Xo�i���Y�c*Q�
b��(/?�5�q�WMɛ�p�?�#5�n�\B���K�	U��c����2^%T#g�����O�C0~�<3ٕ$�p2�c��[_[�P-pR/8�a�xzR`P��Xt$6��+�'Rw�JeV���|�'�Ya[?� NT��f��?,9�Y�^ί�H?�7�wl��ms�:� ��)��H�^C�������e��x�f�x�'
�Y�%��'ǄE�?�u� ݽpDU�b~
Gx�8^�|�)a�ǣR�StY�G����fk k,�e� !nF���?��h aW^���ޘm+�z�T*C�R���Ct���5z�oZ�x�{:�W�|A��Ƞ2�Z,�f�ǵ={�c�c޳��˰6��d�wm���.8�G! ����TSw>��8��h׃���[��/xU�ș��9���ԧ�O;���Y\�`c�m�<v.��vX<Nc~x���@��Ipћ+��6�b�|K/[��)!N��o�-�đ-��fM��3s�s�:�фPt��2іXP�1%�-��!���s~1��f�����t;�:^F5�l� ��rŉ�g���B��y�%�*Ř�:��n����uX�I�4b� �-mTχUPAҷ��W�T�?�9��՚4(�Z��_��*�R�OA��c,cG�����c�o�,=��~����/��rs�P����=w��KP],&��㆑p\\W��40A�Mo�g��]�%�2�����_������v@���7W>$Zj ����}�<���/�B��Y���ؓb"Pt`�ŉ|b���IL~��}��Y�i������{*�C��,tvC�W�8_$I	�c�,�FRo��<2.�QV\
�; �%.Ec���������c�֥G\���+>�7?"�a3a��a��y�� ~��Ι����d�9yvJ�G~�d"{�A^Z�&��KFi�0%�f�j�į�E7��:Q�>5Jo�7ӆ��϶ 74+o�����^8���U��B��n��#�==���J�t�ID)Z:2S�є�!Ѫ�A$�8�*�<�1�B4a܎����⚘�}݃q�`�$�R��W�pX��=N�iM*޿C��i~,���6_MaR����?cYF�)
1�H2��)���Q�T���kt/y7�<���!�E�
X2 ��`�y�����TCJږJ���!�,"�Ƣ�t�M��ANα�/����J�!���,]'�o��w,3*�H�����%�O� �Q�}����'�L�_;,0�ՍP=�����B�?��7^2�$]��r�7����ϩ:-Ђ13K�ث�+���Xh�$���nݖ�� ��I��I�dt,��╷-�!ÃS���9���A�����+�_��_շ�����,Yf��ت-�W�ܺ��a7DtM�.ͺ&G>�O_$e' ��e�MY��x=��1��ҋ��x'A�g>7���Q۝�F��|��(6�|�>.�ܐuT2��e�*"�E��BX�Q��kTC֬t�2W�[Pt�O���i�����K�&��ʜmP���n	q|@փe�Po�]a�O�o�p�g�{��Ez��n��ޚ՘���:�c�lp��e�f	F ~��CT�iP?��l���Y���I<vE��L�M,�T:W�S �b�XE�z��Pp����*��1⿡e�%�R3l?�q��V��ڭkV���Bh-{��=ር��	�������V%�o����X$��tv�X�U�:���n �7�{�fc��-����2����@p�3��ż�H���.�yf�sƳ�(��G5g�0(QR]m_!U�:n�B���v�h�Î�TH�(N����$x��`NIa#��u�m���돠J�ez$��;{j`0�(��a�8�m����|m�&C;,�(nMy����e*-�o���j���w��R3zD?$��ߣ�mk#a����z���m����C �$���rr�~�Q4NΡsaU_ȇ
��%'��[�G�Iڻ)z�p2������+A�����<�`��R�]a&���S��3�T���Z�W��v� �sy�*��"�o�5���	��D�����l���H�T~J�4Ѵ��A
�t�i���I/�ɼK������Fj<�l�a�**�"O�������,Lñĳ��K��(�B��*%���o-*���n���φ/];�ٚ���V��<�P%n|g{N��r���%ә���]� {��B��̔ 񍚿�~�7lvG�)��/Pi�x�g	�B*������mbpt�o��y�A*��f�-Ͼ���YR�$X�%��|,k�c��(�(�����u����Z���jn�"�!Qr���8Q�F�0�R׳�U;a��5"��4+�m��.ؼ�f�*.>D�ή`�[z)h⣯�)�G�����2���B�Ӻ_�aJ9h�F}/9��՞�hH�����§���A
lx���jVW7$��![�����b�
 �dm�J� Ғx��.�]��EGu�ߊ�K�n�s�(\�r��y�)�W5�V��nJ#n�K]7�R�#�����8j��#K1����$:�s�2�@����l���,�����������33��PH�j�ٳ�/�x<����'>-֨�i��O��Ob��n�������(Lљ��
r�Ѡt���� �7J�ڜ~'�F!�˸�JH��j�^"�SC���ǟ�	xh�Q��'�n.*�eNÜk�,D��jr>�Ƥ���I N���n� -���NBb�̕[fƑ�"��e�@2�̬�ͼ��H���g�M�J&� ;�4E��[{������=�����d~Ԅ P��u�2��QX�����������SgM2S#���P��&c�|�K�m��,��}��Ş��K`q�(r�B�k�DP8�ß�+�3���Ʋ�3���S5.��!v�-o�9�^�����+BHP�I�1��	�oKֆ�M�&���l��>I��Vw�sC�E���
`�.�z�@��y��dǺR���\zv���0�wBt�[��T����t�"8�=Y��8U6���|G����*�X�X	�)�ٯ�'i)Ӡ�|��J<��L<Y��W��W8�LW�V3�HI	�� go�~�\�����J����̲T�*3�	��.�]�t���Kξ���]©�i�k���D����߭e;�?裐�"�f�4��Ժ�5�(|<\�q���e!�DM��$:3��Q�d읪�p����h~��֭��Z�ږ���'Y/��[��Yf[@���2uzb9�@f��@�@n��o@�����J�n���GX�>q���z�
A&�S����ӏ{���
M����`nB�ze�#ψTxda��V���R�0�*>�ʛ��d��+�43�!!v:�\�X�/=������0/g�C�f�T�;G2trs�2���r�|�YRn��]2FkR(�fI���ҵ1x���<��[��mk7�ԉ��pn�N"b�ZD,P,��|?��S�q�g�X:ߕI���j��J�^)}-�$d��AA։�����z!��:1kx�+q9D U��dAfpvo�t/*�<�]F�Ʒ��ݗ .�U���D���\�/h��K;%����\m�aw��T�Ja�A�I�u�m�ic}z��5��d�)�����A�߻2l���g�����7��ԃh�l#��Z��[��}h6qF�}pp,�r��J�ߴ��{}�"���i/��HN�'4�K�ޭ�& MC���F�0$�Z���A�pH0�iJ���۱@Τ%d��%��2�j�0g�_)�2قZ�P�1���g�;�'�qGV,�]�0%���
��\�������h��vg�}��~� �ѧ*�o�ٜ$��lύ[�*	&k�cՎ���6����s°vE����/����w7]����{�C���5�S�]#��%���*�'��)�$�u�� ���.DЈ��E���N��@'%>S�@.b�#����&wlYr@�4@.d\bt1��mzzi<#s� k p���4Rȱd�9��ߐ4E��*뭨K v2B6���ק�=��<�歾���������<I��]�'��t����[#���v(����9O�v����2��ɶ�8��Z�k3(U������}%��qK7�(ɣ Vw�7�[��N�g��L��ςn�-%�\aE^�Qў�Yj���]Z?����n��3a6�1aan���(�KSz���أ�D̷�0ע����kl׬-3���@ܦ:J��mT�Ad ���Þ�m����ՠ�kN$�):���3�"�����:?i\0���O���3\~N��~jGo9G����������3�t�Չ8��$V	̲�Ƶ�!����ɖ�_p���g��S`��d%��)9;LB��5Z.L���zY�^�iS�nP4����v�1����2�f6I5����+��ײ�S-ŨC����d=T�� V�C"e��*e*�-k,�#�tZ-��c�gJ�F@��/��/�X��6�c�-k1<)%���zJ�nݑ�L���>����/*v�����ɓ]�6/���B�)��i�<5t���<����*��55A1�Y1l��R�.r���#�2jb~�
)i<;+�Cd�J3:��X�D���O���k���_� ޥ�t��[T�M���cI�bvη�-s���c��˲�����LZK&-Ls2�Dz�L��?�v'sB���?6��j�5_�����W5��`[����_6�0�Lg���qq�H��n�"J�k8�U�0�/@�rS<����&Q�K��d�]!��o�� I�Q�`����e
�G�Ne�ǁ�R_*�T�
ϓA̠ 	m����I��y}�鷭�S&�yVz��� `Ye������T�}��vT~�7�
����{�8��1T *�4#R�z�l6�Z�bE)]���Y0�M�~���6V��8g��ą|�
]��8(�Ym��]���S�CPmS�rIK�<��F:N�6�t�ח�%�/����7˺N�᩵LK�����ԙΰ����(�п�����̊��E��F*|;qk1߬6�"_�q�q12�I�z��[�9$������3��NԼP3l��-<��H;*�a�N��ꀠY�lx}[��c��v��o$�Yax�q�{=����Dʬ_,�"��4Q�8Ǝ�M��uZd�b>����	�7	�»Ey�����ϱ6�������B �|l�a�6�q6���h=,���+��'���[wK�ڪ(���%v��EP��qQ!��J�u�NpP}Q����"&*�K�#,)�]/kY�ws8RD̆d�5S���K�7 7s����$����yʚI�+.��X:�P��&�i]h�����+G��1f�9a�fM_x'��E�{ i��ٵ�S��=�S�O�x8fo��O#�Y�菛��4���F$u���4���v+)��%��������'��O7���֗8�; q�gvVS�^#L	��
;�>�Eh+̾�����-C�]_"S��<�p���`���3"5��]E��L@2����� ��ء��=f����Z ȷ��~�m�����WZ~����t��ޔ��/��`{X���9|~�=�yÆJ�w��>J+*vG��MQk���1�ſ��f g!�|ˎ���P�D��ِ.�n�"|�6��g2g���u��2��	�Ɠ�I��-1��?hځ/�ڕ< �����_xQ�\������{�^��T���\�[�~��hJn��؇���l����R[�)��O�|M�I6�6>`PgF	���;�	�T�T�S��sj�l*�v�0�4UX���-���'�,�S�wS�s�]�Y��+�(d?�l�s=ь���I[5��q���n��&ɜ�6���x[Ă�9b�D��9یȧyȆ�lT��,-	�םw`�ű��Q/��Շr��m3W�'\��e��[#Bt�#��Z*����Ǚ��W��`8)�<�(fs��2�}��1�׿��lRr���K���=���g
���f���Lt�*�0�u��*

��Xx�|��S.���8��bZ���e-�_B|P7Iy����vAU�?�X�S��9U~���EV��m��9�8�g��Q*ʬ�t�)�������ܪ�<�v����w�b�%�(Y��&R:_�@�R���8�D�ˮ����\��C�S�q��d/G�:�iLٱ����-g(UE4�ڶ@JĚ<<�I�6�#�L�u���S��"Ո����ks���h����� �Y��#@�R�:^"���\,�ǫp�R�}�	G r9�^9yC����;],�<x����!���<���Ģ�PJ`�'�' 켊��;X�X�s7'�UНը%�c�KP�v�=CwA�({2�1�5Z����a���P7�*�i����
�_z𣼊�E� �ȧƪM�3vMH�u��nB�|������i��TfTqM����4�BuG6��*�� R�U�2�t ��T����%9�E0����q�u�ɘ+1�E���������@2�^U"	��|ʲ_#��~���@�e�}�E�Y���
_�� vt���pA����dZ�(p�u��`�J&�.]����_�7h��J��	F��T��������0��{r���̅*H:�O��VitJ!K�GQ�3ڡ��Bk��O�ͭ��]�h!�BGR��W���6�O��-Aθ�yb�JЍ�{Y맟��U���{	����R��J���)�3 ~ ^���uA�+E�&0���t�A���I���N0 ���J¶���PS�����O�{���Y;�UhU2���gG�]Ԧg:�b�g�so��>����>X��ɣ�.�4U����+麧�Y��a<�d]��Ⱦ�g��Qf������A>r����w�ߡ�'���i��*z'�,�&���[��!��IX+�-e1��̸��>������f�C�� r�K��t�o��Xz���Wƥ�q1Z30/�H����SH�i�M ɑ�.�܎�W0�]awչ<����ZjmtN��7)����
@����L��qJ���Dgٕ�����N��i����m����������J@�Sp��*�J{��b�� 
ѓ:��!60��&M������L�$�(�fx����������I��w2o4d��@{b�A�o6�s@��y:����|&!B����:/*U�{swrc9d~���Q��cZ �
ୡ�N.���y�����Szvb�v�������f'��k��#����^�çT�pn�.�7�)=t��b|��"��y�S�y���?�M���:Hl��y?6e���|�`��ɑT�.����Պ=
(�2�����4I0���������sD]�����Z*bk���F� ޭ��vuó�6�w�woGF}��!����T͙�n���ւoau������SVj�̡��zU�VD1x���G"�;Q��Oޑ4	�A���(c��ݯ�6r��]�sOe��@/X~�T<���?�&?�
�c����	N�M�w�_#��qE� ~�[�)Ӌ)#�($�(��=y���dJI|����Z��e@������_�/Xy��a0�>1��b�C��I�~��\{�_��}��䥜��4�9B����%h��_�8$�,���@����iT"��N���q[A.��F�gL1q���w�e�EX�� �fb�z�y��h��3��	���U$`4=aG#RB�`�i�!�YD[������f��e�q��Y̚r�Ɣ�������s �ڇ?S�pg*��
ZN(N�b	}GH��PCwƩ��I�i��z�w(��MDqI���Y�m���{J�)	������Jlg���CB0�'�7�����H�]����׃� �L��\�.ȱ�����{��e\{Lޑ���b�~vD�xS�ʝVb��Ӹ�Y�얤��_bdE��DrFu\n*,�����?K�"%ѣ���c�r�/.�B@l��A����+,���$X69�Eא8�B ���U"�/���/�3@��a�Y��`m-t�?�0ͱB�C�lX��0����ġ�:���k���j���5Z�q��Gs�֓��}N �C\ ��D>p�BWW��]��=
�t8��hh9XF��9�=�W�6���l�:��d�
RF�&wʐ���}�(=u+�t--s��0��?��cc�uȃ�ZY�*�N�Y$7��	�$��S|�h���g�6���a�"��4\�0�"�MTr[3r
�X�g����/v7�>�Fk��vun�|��vg�V����o�.�ڄ��*���Sm��g��k��d�-��WyKfDk��Ѡ��ٲ=If|��os���@��:�Vv��Pkc�U+��7�f�'�U��j�}�����?��*�2i�LK�}�����R!ZC������w8VcJ �ڽ���pG�<��;�p55!�%�!*@/�wN�YCg�LA^�^�iY�M�6����R�d���&��j������r�s4G*�t�2����JC�D}8տ
d��6�`F˨�n��y�d��au���C>S�>tf��p�Q����A��d����x`fu�jB�r`�����ዳ{e�|PJb�W5�+X��4�Դ� �zG�
��6t��6y�s��]�� �v�@ߌw��b�ଞ�֊wr�ܮ�w�yIܼW>�$[�,����ݓ���9�^���zO�1��M��L�qy���N��r4��z�΄=+i���w+#�/R~�<߅Ӽ�hk"}����B�p��%I�)������pJ��?�ބ��=n�O4C]Ĭ��f}CU�R�t�xb��y�Л�g1�;N��c}���b����\{m�:g�
tl!>L�"ǹ�Ͱ�D"�/����eA�2'�4��v�!�!'��oM4>G{��1�෾��	֝��x}296K��y]�@����v�[.ӣ)Xْ����*��h���+E��|��������[~��2�\��#���8�~�G�z��x{�?��b�x��{�p�G��]��$5 ;p�Or��<�TzWm_v`���m]4�O��Y��-V�������j���k?o}��4ޯa���~ż�����Τ˵fS5/��l�����b����W��^@��ΆX��� �/W�G<��.PgH-
Cs�'��T���2_��_��V�ps|S���g�*�Re����r'��UAv�$F���Kq{Tԑ���عX�`�φ�s�]p��BV��T��;�9_�|�e�b|Ρ|���kR1W�K�R��j�p�Mp�(�_zc:G�T3ߒN�[���(s<B'���s�7���Gv&��T����b)�w�=�g������܉��j�-Q���>澫A�)�\@�Ί]��*$G�|���pS�ʒ]Qy\;�x���������Yr�!A�H�� 0��nM�Z[�Oz+m: T����2����C����&6m<�� ��2꽃���a	�5�εѣz�EK�0�0�<_
:�.9��Ov��A�~��� �ު��ݒ�TC�l�B��m�L��4Z�`�H�#�����R6��[�di�;��*���U{ؔ�={6�Cw�1kυ�$�M�X��2;>��,x~�c6������c޿1�OS�; �J�EO�(}���i-Z1w&�����9���w�%�]��K&����U�'��n6��fY )M�3D>j�:������&�YW��d�J��(�xH��3�c��(.��L>DZʍ�#���h̬]D26~48�-ݽN���������S�aQA.,��+ɺos�8�gb	b��*� �m�ߜ�z^O	.�"klt�� B[a��8q�X{���c�|��z�2��g��ξ�FȷG"c�w�2 ��煔������Z������Wyt�3���q��O�1�AʬD 9J=w7���p���a�0��Gd�}O�&��6�6]�,�.߻+���3��o{��D�J��I8���X��>Ƨb�T��u�A�b�I�$����g?yX��T<���o��2��Eɶ�I=x=�|�;uވ�)m�D9���_��&����|h�;�����=�uɛ�	o�_a�J�Q��f|_�Yk�;�,m��}�����-x��1�����<E�s�93mޫL����5��}�؉�K��	�`��K]1_��X�E��x���~ĩ���� \hU@�[3#�o��J-�YbB����a����F�gV��]�5l���3���r��c_�!�+�=�4:�$��{2����ġ�t!�<�
�1)C��'!�8?���N�:�ΠJ�*�"�e	��\$�E��#�i�)OG�CY�'ҩ���n�0�mWD*�z>���Ԏµl�~�[X��x�c��3��\*;��b<&>�VU��Ս�7�)��k��`R���# �x�YLT���_`6�h�V��
��49�rvx�#v�oL՗� �B�t�L�H����#�c0zɠjǅp�9h1���?9�x�pqU�;����&�	���1�gZ�N/�H�.��s�^E�����N�;����X�g��|k��b':�AGRE��i��(z��Q�[^a�nER�,l��g�n��C\���=��Hu>��ƫ�N��j�`�:Dn����ѕ��"2
V�g��"��
4����\��f�Y�:xЇb17Ҳ���*3d������F�Ƞl�����,�w��	���{�e�K^����Z�M��skz�=��@3�@1�:SؐrF-�F�c��;RSIY�{���*��&E��RV ���t~�֍��ղ��kl�dr���pG�wQ=����;z�/���sG���s���\�%Z�mL���o���yK�VA<�}Pt�s{B,���C)	��b"	��f����- ���*ͧ��c%��H��Gg���j ����e�:��,Ƿѐ��B���9�g�O0���a�v9�^RP-xȼjk��9����qM/\N1�#������a&�ژ ��i��E���~r4xG�C^A�~�R�,m��
�S�K�������=n5����*9q0T�r��7d��cqޗĢ�JS�7���^I�H&�������!(�����t���Vz�8���!�X�N���z���S�!"�Q�\ݍڶg�R_����x�-F���]ǝ��������$=|�^&�!lY[���-���j�l=�;oh��%�,��Z^��^�n����I���' �R�`�K�
�Uka>����O���$>d<Z���ʡ�ѤF&{`�4��=�q}O�c:׻}����[�1�2\��n7�.q���� m#��*I;�0�8��cC6��ɇ3S�;%�Ɍϟ�*TU�;n����Q���/�ߎ���;~������a'��+_��ͤ�[-�Z�:�MS��Wòp���a��<��n ��ܥ,�4^.��P9���2 P�<�����5�kx�vt'��^l�D�N����*,W���	?�)�6��ߓ�A03�g[�{V�\<QS<},6��4k��\>�t�-��i�9Ŷ��(�(����X�K���u!��ǎ
Q�{3 �~O:� ��M�Z����ɱ(lCGU1��,���d �ܙ�=�q� �q2�gf-_UĤ	'^��6�l��T��N�]�*�>����^�^���nQvP��ɿ�:@^�ͭЈ��th���g�����w�D�	P�ŋw5ȡcW��0���^V������ q��{II��_�9[��>�Rz��k�9!^/<#�P$���5���(I6�P���	{M����h*c�
*��<Zmw �c w!���j,թJ���A��$��*�� y	G�(��N�'�6��-v��4�47���=7�9&�D��P���-����"���	��]��T֡�`;�d�4�����l;��ʂ�4J��(Q:�1,	�u�F\C�o�z�o��!�r�H���B.�",��_���B��4DM��j����I��|�?����u{Jث��o�B�`����]�o;R+M������Ԭ@���@��U�=/�]��po�K{�}�����F�M�+�
G�u>`��j�u���}-�$f
IN6��u3�m#;�!	�_�ʖ���i����)���#F���NH���j�5�q��3�L��i�g[�Jx��P����.������'�J�wZ�A����(��`�/�������bSs���]D���=]���`8g���ٽ�j �C���]6ہH{�! B������Z쪯
�&����تf���s�����>9�f�TV2��#G���rp�����z�hTR�)�)*{5z x��D�8G���eB��MpQ��Q�f}at�d�G�k��Rs�Y
�Iª]_d��c:�Q�뱓����v�G��kA6�(K��ė}������(ƘPi��D������S����g��i`d��2Գ߂Ǘ��������z��[�e<���jh�z,� �XM^4��ML��X�@Mw7��+��}��W<�G!���Du;Z�W��H�,՟�_�M oV���O�J9��m�͍3!ȍ-��K��:�(��E��n/8pKO\����Z�L���$��A�'��ľ����r�/��Iޭ\�<��l���`(�c�f�#)c5�|x�2�SBY�Ή�st"��@��H�aHEG�U|/���ق .��`#�I�a����ԯ������2�s�8�Ё3�o�.(1�;O��`,[}�"��4�S#�D/5�=5���PdI����V��&�۔	&�I񶷊��d��iD�)%�l�Z��������p�~.�7
���^;>��bZ�Tnr��h����s�g��$�Am�����o;��_y�ֆ�T���.5������CI'k�.0�-�:X�_�o��C�8���9�٧��&�p��� �B\�z�L(ۡO>��6�f��]mے�5Է�\�d�	��畡͉Vk[�U,��L$I�`�YL�q53't!�/���~�)�Y����`$@'�d�mJäW?���hߞ͉�HcI K{�+����Sr _��
�!)���h��7?�Fd�$��!FGz���� f?��$���U	'9�EpUԅD�T�.B��x04�[_h�x��u����MU8�;�&�y���ʜ7B���M"������D�p9fo�|8@����]w�,��	�_��|8��`�����(aE����6ed�u�Vc$�(���	iJ�O��y�:X�Hq:*D���5մ�)�B���%g@�5H�F{J[}�QS����_�O���\��ܲdW0i���R����S��:�C�� ��Rtg�t,�U:И��8l��܄��ͭ�����63�{�c�ҀE��cfJư+�yp��3V>%�� �[�y���-��I$��-�����dD�b��H�p�Jl}��b�5`�J�:�!��2��H��{�Q�k�N	|�LO�5�'�j��|�p�,KJ��*E�5�лs��j��<5b���%߷�w��7f�D�����)�#��<r�8nS�op$&�F��Af@iCM�c�d�;����'�	.XkX�Rdԧ�6
�0+��vb�M��f���������|��Ϳ�bdY/W]��06ͪ�o�ҩx���o}f��b������p��m�����INL�G5]SbƫK�$�C�0�>7>>�������'����H�34u#��J��h��Y��u�^z��#x��+�*�2��<З������E�)��h,�zS �iH���Ȣ��!��v���x�IK�S)��Ի}�uT幵'����=+����#,���(.��"O�ߡF���uDs��N�rӵ�+N��fA��la�+Z�S\�=SfO�K9�X�*v]Hv�q���a��!�����Q&��}���d�X!17|=�,�Xf��|���H`\�O���ǂ�����O�*�֖�3"��4QL[[���A�+fA�64u�<��V�?�L����-R9��z]ޠ&m�Cհ�ކ��φ�/������a���g`e^���?H�� *�����=T7�P���7n����X��-�ĔN�rlr�b��+ێ�L5���}�����k6���p%����ti���=0u��hfX���3_�� E���'V��?*�@���X��3���S�U||7�xhm�\�+�M�0���U�:����y}Z�v�	&$�pύ�G~f��/Ɣ�4\��X�� ��tb9pF�C״�ӣj���#�8��}�93`H�k��>�� \�89Ѡ]A����iB}�.?���%�v�y��~l�S ����KۚU�<�D�}#�܇�|E�S:|0e�>������\�03S��*ǁ:,j%jC`g �+%TN�I�Lt`�*ӼA�w��+�t�����'�B�a�R��`j��3�M�����aL�t��GDiZ��o���'&!w�	�ty�d.�{[���UH<���<�a=�N5�{���@��p1]��wH�g��4�e�a�� �{�M>��\\�nqʰ���4�=�8AS_j�8K]�i��q^�S���D㨷�=�h����#G�$ZA�Rmb/LOm�Gr��I����K�t�ݽ�Z�pH�&�����f�SY$�rUW~�����I%�	��ك�9ql��r<�v��%;fU�����U)�b�2�'G�vl��;�:��?��l(>�%}\^�G��֥U��/�^�S���[R`�>[}VY��|��!���N��F��ƒ��2ʛ#A�yA�X�ڝ��\"T���ʓLV��J�T,��Za�u�<S��N�7��T�o8��,�#�����Q��C�.�&�hd�|ae	���{N�5{"{��&{5�V��]�2��xV39�[q)�;�P��G�
;�;��?b�p5ώ}�Kۦ�Qf���B�5��f� �QL��?����C��JT&�5����KݟVs�H����w�=�"�U��K`���nG�[��ׯ�?�L��h %��}+���1��z���R�w/���`l�uJ�Y=@F��͹��$��i1^��Z*s��FC�|L�׶x�c�Zo�`���3��v������_��]?�j�<2gT�������]�%�� #�C�~��ˆ-�!r|�fae� �{$݌v7��~;(�Ç�-S2�������8�2ŭh���ـ*��梭�A���eK��0���R��� !_q
���ekΛ����B#�L2�؏O},���xy�u��/�>�`f�z�Q�b_e���EF)^?� ��VK'Ǧ���PUv�F��@�� ^ފoz�N�jw���7yN�G4x����_��[�����/�m	���d�m�u�	Q�%+-�����ǋ�ܲ��]��)=W��M>?��P��8�'�����p��g��l�>݅3o�cǌ������^�EMo�XK%v��R�=;�{>�F���%��#^�Eh�Oύ7����j�LC����eFy��gL�F����('�Q/h=�~��^6\��&�T�c�V
>z�0掟�����EP��(N�=
[���|ɘ(��m���/��&��O�	@2���vpa]����W�xc���2�o��;	q:��Ӷg���t� "C�J	��p�d2&c���j&@�����Z!< �O(�	�`�o4��h(��}��Ѝ��p��0D�)	�n�Uf���wbpb��_��vt��|��2�+a��^���Y.�"K����}�ђ�3�/��N�3��t�t����޶2D�zu?1���PAT���I�{��f&�-�}�g���ڦ}Ț�j��۬zg�<��i?�9���Ԡ�Xu$��4����d�t���ݍ�6��d�2�t\���m-.)����������w�$g�<l�"	ȷ����%5"6p�Z^�
��=Ƣ)\s��n�W�W��o�8X���p����
��Ѫ�ޜ!ƨ��8$إ�ΦgP��x�v�_�^�âB�=4AuZ$�d�l"v#�ڞ��vG�f*Q�	,R�j��f��,��_�6qZ���5c�	�) ~���ߝ\%fi*m�8�|?��m�!��BB�����9h����!e�t��A���TZ�����4�a@�	uM�`��0R)%_,Iw���_r{�U��eyT�Wq�c-(c(� -��l��879w&���^�4�͈��$�I8�Pϟ�껮i�A9��E�m(�u#g��4���`��᪖�
�V�,LƳ�vУ)Ӈ���gZ.ۜ�p�yH�/�ٌ:�K���4����1X����?q@9֛]aD��VxU3��W��׵�K8>��5��n6��K(�G�|>7ĶʎSo 7<4�C��	�¿~���.�@� =��8s��ϖ�d�yK�D��p"�6����>��u����߀�N�\G ���"T�%xL��ͥJ[����2��

�� ����p�JL�;�,��#�E*|���� �I5t��ps��?�~a�}2���P5��QFC�
�]��<��+���q���b�1�)�տ�гl{����r0y�3ե� -;���ʹ����!KЗ&��J�u�J!���;rp�Q�^?~`�_���d����{F�,Xqv��1=ikj��n�Y���@F��C�l�MQt:��)�.�?�fE�1���s�=�xy0�L��cߴ��B&G+��u#&E���WT�!gl�p����h8��E�u����N@Ĺ-p�x����9"��'b?g�x	��-��W��Q��ڍ�-�i�+��!>ζk�F~�g�M'bZ�����"��dg��t)����TB1[��<e
�<�_��kw�n!��'<ϓO�K��"c2�Ii�����t��ϡ��&G��	���=fzNRX�U�e��3� &G�������C�0�m'*м�;U��H�Q�� ����wƂ�&Ň�ZI���T4�+xI7=�/��D>��˿A�_��q��$���w\?������QR�+��I�|������_K�X6���E;6�,�%>��[�L��
L�T�i�:5�ý���BhË�Bۦ�{��z�q�mQe�L'Yx?�.ax^�$��OW��o:+
^�Ŋ�:���z��6�����e��#�6�b��а���Pݪ>@�est#�<�� % +�ԉ����v�m��	�<���Q�v�3<�
�n���3�.�'�x��CC�ZȺ*��ʰ���[�3�^��${H�e-Ӵ�L?�DĹ�n�&`��g���R?���:֕1�"I�����y2E0���iX-�{�j#�=���`dh���Ԁ�7��O��W�^{��8��̈́-#�תBUq?��Ń�`�^������1���&?� y�&h�f�u��|sG�z�0�-��KZ����`wN|"AT%Z��[<�X<�F��[�L����&P��	aq6��. s-�V�-	�eM�5�i���$��]V4�R����'�qYԠ�G;�h�����i��t�*���%D	#��KKC����(� �-�����?y��q Q>Ε^qid&7�d��uQ��d���|��<#�&�k����kQցŎl���[~'�2��A�+ʛ&uĈ4U��S�H׵K�Wy[3��iW�n��`��;�C��>&�sr'�I�,�XM�����$G,�󽜾���]��r��i�dU�q�������Z��}%ד�St�k�0�Pꅇ$�a(�ݗ�HXm�6�{����JC�G �pOuї���[�A�����2=kb�J3�ʄn��I^�l��a�0N`]d���[񨨹D�1}�۳.��w���ۋ�_�%�Jx]��s�:����m�yZO@��1HDS��4ǝA�'�T�Y��P��:CW i��l�9���զ�챹��aWY�8B�D�!��R�4����w�ܤ�H���!��R��:[�;Ș���� -�kl�r!5��0F��LӍ��)4��U�S���l��ls���~&�V���_�"��s�D����*�%�f�1�=�j�1$|�����ޭ�LɈ�2/� sE���𑧑 ��0D���>�NK#{�mJ�G4"�,j���a#�f�i?NI.�j>z�[4��~_�3G:��)ƫ�m�}�b�ki \��/�麫I���Ty1�\ڿ�^L��zFYwBcZ�#�2��`�\5��d�#	��e��ɀ{(/��;�"B��N�B�����I<�F���]�k�T���ϼZ�Jo�Cx���Y�|d��(�H��Eu2-��66ST��,?#���Ne��r���w�A��Ϯ}WI��)�&sG`^�A��p��N�"[u����O�& ��e=���~7��T�y�M!���*6	��^s5\����F	��&DS����M��H�S8�5��I2]�u�I�&��y�<�*:`�S7�(��X��<��lw"`�����^�W��_��u'�h��$����p����!�t_: ���װ��g,%�����0�m_RG�'��٣�o�e�=nX���۾uuϐ��������җb�y��^��-�
!�,Ù!��u ��m���0�-)���\��%+W���l�{-J"�1&��{����P�U"i�i��b�_����*�8TR��A�
�C��  .�G�Mp@��1(���k���eV����Ͱ�୮N]4?R��[��lEa:�-�.��� 8>xS�vhE�t�q�O.i"ٴ��U��8`k��b6��Ⱦ�lk�}~a�P���HX/
�?����JT�.��$�G���מ��C��7� 8�YF�?�7*�ɉ[BI���3o��Ɍ�@b�����n��|k`�c
�T]g7i_�yT����c�h@M�Μ,�~��~�D��$�2Tg/�D�-��'��r%�7=C��c�p�����~.��v��#.Oъ0M�N�-l@G�Bot8{� ��=�^u�5puG?�!�����E���OG9�C��B��؅�{>��k6��a��k8�f	�X<�m� ��ʙ(��ĭK;xcs�9â@�A#&
mT;�g[����ɣ�z~d!l3z��ݧ$C�0���~��ֈ����Ԟ��G���vC8}����U��~z��{�O[�vJL��x�4^s ����:|��i�Dkn-�`|	_iU9W)4Ͼ��Q��XBK���>��`�d��4(��I���	
�؃��m�G���R�x׶mTfK'�su�Q܇�&@!���<�D�ZΪc=5$���y����(;�c/�m_�9i��d�)(ߛ�v�`�o�5�4U��f��ꢣ)}B������*$�Ý�a��^��k�Vn��r7�X킐d϶S�Ӗ��W�Lx�.�@)�g��c���7g~I��z_�i���$I�vGH�&W�:������'kQ���u��/� .{��;��?�y8��D�l&��[�c��ld��_o�@�l����y,�>�5�_%��d��5�
���T���[�=�뚶��!`"
��s3�}�	%�M�_�l"��kv52�O�ot�"|�%D��~%<a?=w�9J瓩�`J=)�~�T_Mv__i�;�ʒw�Y67�Mn�J.�?����q����hi�L�5�YyYLƶ>���n&��4����([�>b�Z��Ek|��ɵ�����Eh-V���im���M�s���B�Ҏ��U�[^���i��s���h$N��24g,+*�X���Wx���8/ƀ=*{"j�����і6���C&�+ޭu<���=[1@��</}�~!X0�&����СM��S��3SQ��lV�&�+�M����"ޕ$>�3�}l����;�͏h{οj^���Xk���Cfܨ���$9�A��[���Z|,��8�UD��7W�8WJp��׎��,�+��sH��io�Dzm��ۂ�%ƪ����L�&����3|�<i9�O�t�JY#�D�m���S��XH��x�e�]�L>����cȪ�~�ny�5+���ΕI�m�h+���D1��l��o.K�e�Iq��