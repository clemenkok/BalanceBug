��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�!��
��%Y l�׾���b����Iws�h8&� B����.z!'�=K�^��6}K#��i/󇡜�`.��D)|�SbԈ�}Ys-��oYa��^��y�2� i$$�\�n����<3gq�cEd(�>����zt���Awm�	�f-�B�ѻ,ޕ��j��?~�Y9#w�l�K�*e�T��r}��5�٘�n�؇����O��U�xs��a��b��U�eR�`�+��s~��!k�f�.T��,;6��|�?r~|j�j�`���UܵD�Y�@�����[�7D�
aa.AA�nN����r���H��Z�y8��u�����"�������n�GbT��>g��I"�[:?\�//^������ ���|3YY�ʁ��E�B���:[	���9Z�'���<��.�%�#����[�~�W�	E2� ��&�H�Xg������H��}��� q{��Xe�%7 �!B�H�$t�I�Y]X�v�:�S[�WE�� ���#�3*u�o(з����#��/����3坙T�»闢p�҇�}��F�$���[-Ҵ/��
� �!V2�▖j�6�"��m*�/���rW"K�c�|2_;�( ������GB8,�[����A����?�/�+G��w(�8��P����v���aւΦ�l�������@))��!E}I�W%���G5��1�>�a"��"d��ϗ���o�4Nb3�}4��(�Rbp�q�D��!�s���Q��a����}�@�Ԩ���PG���F�=<�d�pİ�:�٣R�4}�3�Ƃ��~?� %�4�2��8?"�~reY�x�\���f=�n�!��xa~O?4���g������R�B/#�N������?�żi�*�/"&h���P��߀�&�ОG���G�"u��ѕ��(��?W���"��p��������]%�������R�5��A�aÁ��F6�4��5?X�5|��ʾj5<�Gw̮n���ܒ[s㱫��b�j�V�� JA���g7a�Cv���А�cp6�S��K��%���aX9 �+�41�I�Gn�0���>C�Bv1<��s���V���z0�GG�]�.a��.�i'�)�f] ޖ�-69��>dU��~(a�lJ5j^IT��6�f�RL0��� ��+\������cx��L:)kA��J֍��d�\�0*}���]`�u��7��HV_�M���2T���P�B��§�v�L(�C�k��5��w�Z�M�ܧ�yw(ĉv�L8���;?�_$ n�i�G���z�A84�V��!�1ǚ�I0_�Ɏѕ��_�"4�rf6�3s��cӏ���N��Z(6�����D�xڒ�I��Fǲ�V��3�ПmrJs�d%�lϕ�:�'�,lq�c ϭy����(��f �*�?(��,�-|����8yT|F"[�J�/TI_�ې�u
H�\�5m^��w��S�w^M��g�O�3x)���s�'34��qԫ]���nS�W��N���ܾ+������G�K���OQŅ�tu�_5X	�����F@�V!�5Sj�h����z2��i�L����W��# ��%-V�
����Y��	)�w�ڱ�������Ds*�k�b���J?$SMߵ�φ�!-��(n�n��>�k\G����"*TQ>|P$� be�e�bHr�\"�|���h�x���;G�yw��B�uL�-=�U+L�_�n|�^���/�	����dا(�
bь~�wNB�X rP3�w�vDĸ�X��>J�YK�[���i�Xu�%K/��HE�q��6s+P�I
��{l3�{�b���~����E��^�p�!:�Q��-k4�6I�i~�MN��=��lk��b3�6�.4��k0�D��R��l"���|�a俕ͬZ�/)�h��vt�b\�IG!�J+/y�xk$�)�UvΩg�ʴ>u��H��J��HD@g��,��N�o$̜V!>��yu�ehnR8�e�贯0Ϥ�ʿݪ�a�G������(��hȹ�Կ/q>����뀥c����#k�0)��K�
�O'�ɭϼϖ����|���/B��k�&%XsYɄd{�h�2hr���7t�Eڀ��2�\<>/c�уB
�ëyd#�φ��l<��rH�O�A��� �E�y@��� .�3쳠�����e�{���J�� Y����*�id5U"��k���g*�^g����zG�b�(�����