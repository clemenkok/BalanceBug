��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�!��
��%Y l�׾���b�����:��@��\w5wu�S�Z(j���!*�����UxA�@BY*ޏ�4��{�Hi�]��
h�J�O��f/�dY�V����kEHn@<-K>��vf�e6yx�o/A)'�=wMa�T>ΏӠ��w\t�����v@W���U/�?�E�q�ЧVN�(�z��9��2���R�o�8א��D�h�'�ߑ�〞Z���b9�i4s�|,��e���C_@����U����H��a;S��>�\��6t���H���:�z����Qpn9�=��G�%�H��S�|F��\ �֍$�_$<2f��_���uO"3�sAY]��eq��6�aK�Ht'k�`4S}喉.s���lLu���8�ϭr�~�fj%���+⡀����`s�v��| 8�s6�u���c6:���#/)�j�%�m�(G"����ϸ��Μ
Th��&X�_�2���YT~�B�m��4���{;�����q�3��Dzp����9���c�g�v2�8vI�+*��c�ul����'�T��`���m.�Y�X�
 �� �)�)*���(�݇N�/9���		ʨc�h�y�bف�OJ�;����������)�o�uu��}w}x�q�b817$:���G/�?��J������$}�G����ؐ�Qa� �/۝f;���.��oa���a
G,��E�W	tT.z!bb�ʧy������@�.�|����ʁ����tע���uh4\��)�(I�%������qy!���Ѐ� �M�8u��cbAш�yc�lP�5�L*�U��<��ͪ��I��^�[U�B��0Q��A}3n�G���tu��%?|Q�s�|��
 �w=榌L����"(:q���IHހ���'w�8���$k��Ď5�:}����խc�^�ಪ��T@��l!�Ya����L�sC*G�>%�D ����;E����9�RG!,����C��N�c��p^��]6��/ݯM�5�
��u��8�{��?��Il/�Q0qs�b��,�3tC�dP�ѐc�턯ϻդ#�ysc���x�4|u������%�"I�$�(�A_}.������bzs�Z.�_؆�Z�����nri]��(2m�UBv_S�8���ė3PGg�O���v6렎���X�^�L�J��_P��q:JVMk��D"S�5�&$Z�6o|�U4?����ձD1�A9nS�zb̓� �Yr�?��z����֌��6QҎ[?°���5>D� ��=�Y.��L�t���B':�*U�5y�B��g�����@(j���N�b��t�G��8������4�ׇ�I�1�X��;kl�M�L��P#�T<�S,�ie	���輢zs�-�Q�{�=����H�2�7k�W|��&wճ�g�ŹI<�	7I\�)�� `e��"Tt�R�e��LA��+���+��P@�1;��O�`�y�&�tÏ�m/K�Y�I�Wd��l��|t�[T���%�i�*1���lĈ�Q�3F��c	w�,N�`_���B�p^!��yE�BP��]���8n����Q���l�L��8��`u~����q[)�em���s󺓘�NJ�������_�P9= ��t�m�k0?U�m�ϵ*K�
[ɡC�a�l�4v[���ۤ����{u\�� ���n�d�Gy�aZ�h�B��o5쨜^�����s�N��
m~��Qj{kొ�)�%�w��G����Z*�q�`��Y�!�ve.�"J��U��36Z\D����&6���������Пhv#���)4-^[�,4�%\�?+���׳�c9��
�Jd�tf�������~�w��G5��V77P��=��(�#����K<�Nm	A�w����Ja7T��W������$�;7�d�s��/�ް��bJl�.�`>hB���\ԩ2X&�! �u�:yKB�7~E�j<�@z����Z�o"ń��[�� }߈#w\w@5ш���YE^��ʼgB��ş�鳱ǚ�b2<2��~+���E�Y��B@���U�	P\�U����H����ͺ�{��}�����B�~24F\�!�0�L�^�9/}�%N�g��W��C�e� 	�6�J+�%ji8���M�g��ض��r�K�c��L�:�]���cr.�P.=�g	Y��عl�����e������D�Yl I~�<�c����n��bT���C<(�G*�[��!�Q�X�
]]c@�C_�c|�%_؄d�cدk�M�@��:�i�nB� Gk����-��"��j5��/��dv�;�[U����4�vu�pV����k($�U���s����=�����D�aV��v"��M[6_�hD�^���^n��Cu#:͒k���&)�+��tg��Ib~u�]�e�>�@����ʏ+;������N�Z�����:��9�Ԅ�^FN�-c��}������]nv#2^�f���w )v��?E^$ڃ�/����`�-���dz�IC�)�ayڌxt�h��dNv�Q������É?!8Y�u�T�(�� ޚ�vy�G��q���V�~wfː��]�K�F��/��1嬃aY:�I�ߍɈiD_�:�����|>M�৽9{r�8r-�ݣY����,<�Arj�	����03��^$�)��U��/.+_ �7
|��_l �D���cC����dyw���O��
}��MDcBT��ՙ�H��Q�^/Ўl)�dCԘ���Ag�����lɒO,�-X>���i0�6b������,2̱`wkZy	��!����
o�xM���<�d�^M1?�+�����������c5�C�AP��F J�b��a��F#I�����\��Ѕ�_�#�p�X��gi�{���T�n�qf�����0i�ɐ�u$Mn��_@1k�"mc>� ^c����wДpF�}ۗ|���)�