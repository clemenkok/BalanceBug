��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�0����L�A�Sd�����y8L<���/ `r�����|Mo�<	a�g��F�J����P�%�0���7��]m��4�x�BC�g�<w�ў�l�0���q@�ugQ��b��o���h�L�Ł:�^�Xד�\�S��k<�*{�G���Ms� ��ΜT�翀�12�Hj��c�UĆ7��.�Ύ�uA�DO�U�;�mQsʆ��W "���	\�f5ނ��Ę�>ʲ�'�SI�t�2��80`�	j�&�-�͘�ۭ2��f�`:�Ԕ��?�B���X���J���'�_(E������F���]3��(�)g�,�	Y7�����a�����:�e� ��n���`48Tg@���K#3����H� Xg�4r�ދgJ�e��U��y��͚�:��:������x#��A��27 �o@��{De�"
Mi����5:�vH5�Υ��}����6��+�e�]�|So�ܯz<�?Z�d��a����go$5Î)�����]��yT����M2��F#��D-egc�S%H�q����!���]� ���(�f��&i�G;5MnYR�o�g*e��v�$�4�Gct�`�Bt�<0�=���AX�)�*q�9,u��t��V��{�&hbV���;��AU�a��B���L�Ⱦ\�����
{'Óu>?uz��'/@�[Zo	���6�RjÆܽ�P�0�g��|�����a���3��Tm�L5j���m�H���=,/ٔ��Ko��O0gfcs���A�X4�Q���`���><������\�e����0iT��	��RW�d�X9��nS�aUv�=��m�,ew������;��}Q�=!A�t��(�,�� �Y�{���)��m���6�z��w�"%X?��Ķcn��\�Ʒ����=�6ot�2���\\�=U���mh�8V��%��
|A�����{�{�d��l�N�q؇�+�N�.��>�ܰ��rP���܂2��,G7v1ԇgmLW"�<!�ܞ1���C��Y��'��!�n�<:�����}$i J̌h;NR��rU/B�v�����I0
���Dw��N6�O7ƭn��9ȀEW>IH�2�z	)-�4Ydj�����h��g�yF�v��J����8u�kkWt�����6z���0���_�.;f�-UI��m{��kdpxw�ۚ'�yҷЊb&)� 6­��U]����\�B&�]����	���W>�<�������L���5���o� H�b�vk��$M�6a����t҈l���_"�	�B����Ψ֔Ú�6m���G���.���G�YWL�Q��u���sY�	HT��b󟳯��o�K�g�34��d�ž�.{�_ΗY?g�ba?�W�#V�R��x� j�B�[Ҕ�o�q@�ħ�-Pj��2�/B� ��%��0&ږ�NK�V�͋ń�C�9G��(GBi� J�"C���ǉgQ(�9V��̮"���G���z��i�Gl�ۗ�.ttA�WQ�&w�Z:�D��U�=@E�d�CoD�� �ϼ�J���=bf!T��._��!SvoY9�X8.����7u��ͱ�7�p�ɦ?qԚ�6[�s��c����))G�)�N$R��s���)���j��������Y� ����<9��']0��N�����j?�8�t[V7�f�h�ߊ��J�sQ201��r$c���#"q�W����uY�J�F�7u:e��7�g}�ڑ]Tڲ&�Sx�%�U͌s�nHTD�|Ya��[R���K�^!��ޖ�YS4P�`h�ѱS^�ib�C��υvaM}-��g����
��-�ԀF�����SC���I>!����4p�����E�m$�cs�ˬ�6�	����\3$	�x.�tq�4����=p/��b!�iN�P�7d;�+�?vl̚�L�9A�!� ~!����t����3�Y��|-�����_m��yԖLdv����$�p�1����s��c������,d�|%���A$�<X�38���~�rҲ�Z�
/$�Vܽ�:`��Yg̛V�D�Pg(�.}k���0��Loe�tS<�HX<�Z�Pg9��@^=�g�� 9�wQ����@�B�Ã���"쪚����Vt&S񖺂G}����+�i0�p	0C�Ū�)��$)l$@m�i�8
�j�����|2w5VX�~�7�iWj��\���]����P�&y9�4`�>&��`Y���|Y�Pv����~���ꝞP�W���BO�Q���.�LǕ�S�*�R