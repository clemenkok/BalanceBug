��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�!��
��%Y l�׾����|R�b�~�I[Gb|Q3E�_����=9��Gp�mv
�D�G�x�ol�'��.ͽ燢7>ߏ��=̾��~D(��~j���N[���i���t�V�~�*Fw�t��	��,�[(�k�w����Ri���[D�e�Œ�J�b	i(�'�(�����
�i`p���xtJH���~J&��+�"�
Z����V�S8�ÿ�MA��E�^���s����=9��룼t��(�80����W�N��Sd�X�ދ�j��4�7�f)J��X����mEC�����4T��f�o�}R�q7���x������)f�f�8Mh��M�rM>��O�!db(�oҥ�x_aA��zP���U�$!��m�YW=K����V,naۗ�G��B�= ��3����1��1�d�1J�!�K��1�JЃ�7�	�`���E:�_���Y3F֠�ԵG��.��֧��}֌H�M0����X��m���믬NG������b���Z����/2�r�{��mn8e�_M��))rɶ�?�3���E)�c��aj���Q�P����2�۷R�+��o?�u{����}g�)�p[v�D��y���l��ƴl�k��-���m���~��aovU�<I��ø�����f�f��+=J��JHOt�Q㾦]`4�%�OX��a�6����h��.]0;*�ٍ�ö�h�#]xp�@�m��='��f: L6��E�{ܑ:��v;J���՘g�1o����_\�A��o�gH�Cj&o�Lo�!�O��l���=1�5gGhqqUxp�i�_,��:Q��<��*r(��)Į�C[%
h(��%U��,z��O������7:D�Y��eR5c*��n���q3��9��zz΋e6/:�+�����Z�%-Gɱ�P�;B7�Pȭ\�D/g�ۿ���<��j
��V�OR;U^�SG�5�?��:�Y��Y&+e�� �O)�?���?�{�� ��$ܑ5���Fu�%��K�Dy#p��M��Ku>���~Ӟ��>ZQ�c����bEQ��ϟ@�C������Ro�[Zقm��cP���1�����{Cq�/"fBKz�����l(%�4*�:�#�9EL�_���D( �:8�e�d�/Ȁn<� ��z����K�IB�Z���15��5u.=�jG���`u�?$f�*o�X&y�1C��7��*����WOЍ}~����+	���&�L�����Yզ7Ʊl�������$~J$JpV�<1���>FC�ȣ낋��:��F[2� c1}#�`� ��p��������R�ɑ��om�
�j���O�H��Z�&��8wQ_�����-�6����˶�ZH��� 7a���J��-���x�6�+|�ӟ�E.���ZA�Nl��XL3��n㭗u�	B�a_����T���rp�ԥ�d�w�腼�q$kvۑD�,�n��π�VqA΄��5W�e���	��J*�6Ī�8=�1K�ށ���i�H&�z-����+Y��2}N�'�5F��U�N�s��Nd� 3�Q)�
�Wn�!���kv��ֺ���Ң=�E�<�r����
�wJ��b���D�h��m7�ՙ�fYQ��B;�/W@��݆���f���x�fJn'W�����&jR]b�q��bl��S*D]�kM�w�`�N�l1��N�F���?k��W���_uiux��5�s�\���v4&����d��N&�\��F�an���'�����`{�)��Z��,�V9P��A����?���@�&S���n�M	֦C��Q�ʱ2���Fz�zfU_����@��:���2�&�S���QVV��Wٝ��5�>��
'�V��.C�r2����8Dr}���ĕ�/� ��A5溁1�qrBB	�|.�X�^����P&v
?œ��!��cM�x��D��/��;e�1%��~�>J{��AN�+yX&���F�)#�	�]�1,YD�'�����w���g���R��ή#0mGNA��Bҫ9kx� ��K1}u��X�E+G�����@x���d��EG5(��g#V�|0��L�W��,�{��ԃx�Fw�� �:�����z��@�e�"�@��S໶b6�0h��9N��ʛ������6#;ƫ�<)�e�;?5�bݳ�Ga;u{�P=`�� ��\�R��6Z��!��z��m[��/�H�g=���Bx��AS�W�y:d�"��!h��d��}>=����>*��A�G�Pyo9���څ�C�\TAВ�����A?�����z�3D�i��hI8,r�7�vI3`S-$n���|��Ӛd��&��}L�w��� ^�^2$H��3!�De�.wR+V��:�"d����h�h�b� +���{##���o0��HvV��`��S[A�=`��g^���}�F:��Ɇ!@4�$�٥v�@x���j�R�]�����{��B��A��U~ؘ���	�w�h
���0�a�}xo���[	Wb�T�m�:��N���ѕ�;�7*�u(Rl�
�x�z�3%�H�~��,������f���Cvv���4�&NϦҿ�d.U#��i��Â��|�['2ؕ�X '�����<�Gr�d��s�V�"��po%֠�0`�9EO��O g&�=*�j��I�ρ!٢�T|�4�K�N,�`��D;X)�PO_3;�٨�ԡnJ�9Ya� З9A��-�<�!I��L3���$�����Dhـ�I��p�)�(���b���tP�|�zl��Yy3�o�?]��"���r�����y������"jթ�ʹ/n�J�v�\�Pn�~�'����F+�SI�ϻSJ
�=tGn`�Ȼ��<���`.ȆW��G��2��F���]7(/}�6�����p��78�kb��&���S>���p�19�=}cE��B�^���u�+��G�*A��m���幋K�g�n�(�R�UH)���8fr���k],*:&
'����~Ug'F<�Ȍ��Ь�x�]�$��s�!�y��|l��"�ȃ&14���J|�h���4�^>Cd���x��v@!����q��F~��cf������e�()G61�>q��;+���xXCN6��"V<�-<`��*l9��CnmW�[(�����Au�Q
�(x�2:�P��(��=�ɾ�g=]�V �����F�،�:�ǡ�7Sߙ����
�� J���ꓛy3������V�m�DN{��:��	��h�U�+��/��`e�P�ˡ��E�	.�<�C`�4D@9����������4�����n܀���y�i��F��8�x�q�F�üqṂD��6�A���T@p��5!%���0Cצj�QB/�$=EV-
{�n	�gv��(\��ql��N�xY���fW�������PO�Ƿ�m����PsD��R`���A�h*Kë���u�9��(�Ҳ�@�ngm��7�qO�ʃ�������!���Ȍ�! �t8q����ɏ�O�,��'f#)M�}����]��.���sZ��!+��bu�i1k0�<v������MnԳ �7��j� P�N�贲/Α��L�Z�j����0��s��o�:�aN��n�5��8uѮ�%@��4M��?h�?U���-ߠ�Λ?�풴��7!�c��b�*!��{�8�XY<u�aS{�#��[���{]3pƏPlH���<��#8]1y�Z�J���(���-��˟4Мtn�]@�'ͩcopf�<a�dM�3@����
�V�\hb������Ӗ�2�p�痌�.)
7�Q�&,3��&��@V�GGL��y ﹤kUr��8�`*�x�üZ�����?Ap[U��=�g���2�EB�gn�`?��HD���isB�l����]x��J��͠���:D�r�e���z�qoF�4\��z����3 J�R�"��0�(-�*]��9�L���$�:R��?��8�ŵ�����nl/*Hz�s���I��G�a�No���&鴗�t���XaB���9��+��g�@��b�S��J�sݑ| ��:�2WR��Y����ꔿ;@����u��ù�D�d�l���ա�'}��������u�k:v9ǙU�ܦG$P��.jv��b�Z)�)�����M�6	PK��BIW"@�zhU����������{��<C�j�@B�i��wSS����
�������K˓o"%͈;���W�=�0�_qJM�
��B�32�ည�${x?����s����JK{��$�8&ϔ�ow	6>�%�����m�x�@�P�8qDg�R�,���~�p��Cp�匸\+=�ِ;�8�ך�C��.��~�^76(�0����P6����6xO�@[iR>ٓ���2����BC�>e�ð��i���+��թ�e�M��K��n�\�O�z7�j�6j �*�Q���\A�����x�#3p{��a�5��I��8k)��i+��4�	��D�ֈ$a�Y�'�?u$4dKSB�ÆD�@���V�Z:�[��#�R�ఈ�^�ў@_�pM�t����o�E�e�,x�1����&���?���W�t��Gz����>T���-����^Ӏ�����1�D��֐P�P�y0.����� 9×�v7�8)\�כ#�R/k�?p����E�̗tN���GG��v]:ƍL(ծ��2-�OW�R�'зY>4��+/k`Б-���9�S�t�3�Z&!9��d�d�D�w:)�M�Nq�9e��Aٞ����ӛ��Yuy�%�ĺ(���p�p�9��d7/s�&�闛{���`��y���j���֘Z�\������<�V4z�*����D�����G�)��E��T'6�0����uo���ɸ��A��Lޤ��o�g�hF�1��k���c��M3p1�IO���-~d�/�3��FǯIa<��V���_�ut���|�nE�6��N;T�%�Xi�"�m�ʓ�p� ��NiF��rw�P�b�?��(�*s��{�Lt�:�����i/��r�1���f��8�r����d�����%^��<So;pu�g�^@���z^R�+�e,-oZ��+Jz������J�*8�~���IY�U�z}���N
��y����	� � �E'i���JZY����l���aЎ��g��=+�Ŋ P���_�<"����qr7�߆0�`��0T/�:��Ɯo���J?�Y֓vi4�;?�<��%eב��(s%����c���L�+�!-�'�ea�z�4�@@�r�������K �b��废!0��~�zv��ѿ$.�����G<xk�K��O��~Ʉ]	��TU��?<	�vܚ�<�*�D���S�:1ޤ��|UF�d �I}@�ӝ�d�)�?%���!F|�Z/�P�-�.L�Y��-�6���2�	�$b�Ǭ&�P�ը^EP�qv�`�IDy���cm�P�箆gc�VM�S��6~�,��B�L��a[_�2���d�9c~��D��{�㇃�*�xuy,�x����ᜐ,�r>�7�UQ�:3�e��zΓ#� yc��6�k<�y�a{U���`�/�@�P�a�E��O3�v��Apr^O�/&�g�) ��_d��/?P�"/E���0�!N���y�r)p���Yb-��+1�U��Ѳf�eՀw�㶭����@�_A��m��Ӵ������;���_��d~  ���47P�ǚIj���UF(��Xp�����>@84*�Ç|->�h���"�_������>�L��C��)�T8��v��G�Mi6�ɟ�� ���I;I��p�#AcD��әĭ��H\�۸��2��JR�l��2 (_�#G��U�m*9{P�ԦߛS}��-��P�l�|�YSCo܁EW�_�r���?N .��� j%��kG�<XQ�z�3`ơZ�M���bmh�,E|��`aߜ�z��̽�jW O���lb�P[:���o��8ua+��S�^SY$HT~�w2�ӧ�[��� U��J���p�6ݱ�En��9vf�HWo�s��D��$@��X����*����&&�kM�4�9t��f\�*�������րI�ҜM?m�33ibR�_6>2�T�rt0z�R9$��	tVq�!�q�t�~\f�*&
}����^:�n��!�p���!R�?��c��b$�P.�X�_�Q)���D���ͣ�d�����i�)��@�oB[ꐓJ(�p�h�90����ǖy ��R����283�0��'1+®a�`9�6\e�]�Jph5?��
3��`J����óis��s��gؿ�R��9S�_����x{�-^V��Ƌ����1�5X�`҉��q�fY���k�r=�Bm�z[6<�~U�d��#�4rC���~"�κPj�W�靓1$�W=RC�Q-; �C
!�I͊�o�Ů�wv� �cS�`�'�M�Y _��
o��M�3`}�cEw�蛬�:��,��k3cMv����K<�{�~�?��n��en2��g��~�0���i�/�p2��� O��_�%%0�"�`�UW"��Q*E^��6�m�/�(r�ׁ� eT[� Y�߷a����$�m8c�	��2w���
cV�%.aJ��t-��@�rC�6�&7\��*����?���ce�e�+r�����GV:����[�Q��s��ꧠ��X�J�k[���_i�6��6Z'0�/�ݗ���8^4�震{�32-A��6�w�v4�+R^Y��˯S�/��+��	z�Y����Ws��["A8Jx&p�CE��C�^��V������&!3�/��L��Z��~I's�w��ea�F2zj>{C	����M^�Z��>n�vC,�
J���l ��O8)�M��Z��� y�m��K@y��Ϗ;Ps�b9D�boƔ#j��t���dC'� ֝M5��S�b�&�5��Cxǈ�Pw���]>���	c���.}>�,��m$#��gh6e�$	V�a.�)�q��y�F�1,��x*���o�-+Qk4S��'rK	�	��6{~J�QG�r�����ݯ-x+w�7o�n���E�KQ��JTL�21Da!a����M0�uC�i�X�ִ:q�����|�,���b�0��YB���^�r��]ҭ}�SO�ls�q����ܨkiG�;��mt��0B�
m"�W�꣓
����V�)��d(����YV���3*W �H�]�so�؇*�_���~	�տzx�~�(��!��<��e�yFlB�,6)סRD�&���M6�R9Xk	����j�3�Қ��s�ҏ�%������</3����g�W9ޕa��ry����	�`��"�E�_�<��*������X�L���Z�6���t	���ňrs���p���1������;�V�T�@�er'w�e(�U3i�|ce���3���QH�P`��~�a�M����|{Ҟ41T'�t6a>�cu��ȅmn� J�%)PB0�����}#,5��GʟR	�~�BP=~���ՇW(8����clf���1ڮ^ހ���D��l��\Ĭ����:�qD0���H����< �id��p�D�yg�LÔ�S�@-|	
6�z�Ku����`<���<��/0Y붶�Z Gj�Q�Ȱ������~���X�Wg����g^��WEw�.�n~̫8�3��"�7U�!����OV�vc�j�v��e%|$�SD2�h��9*����FD��닛E1Fc��И~:C5x�jт�y����i�&�q`h�+�����O���=ʴ鉂.ʐo�C�Rp�g���m-@Pc�T7P�"B���m;Ogk��a��<�	$���
M3z��Ą�:�;�^��fK�G���F�`+�-���)G�����ԏ�v`\�P�#K]���HU-�1v��Qy����E9�9��4,,s��*/��4~�)��O�Ӆ��!�ԑ��R�X�C�5̨�_&��a5��\��L�q�w�I2&:~�G��|����U����*���Bc�6X��U��=���.�Ӟ���o�u�*	�?m��^Rhb���0�2�?��1��A������YK>�Cy�O9� t�I���CO�1x�1�qlڀ�r��U�g�)Ep�ʤ�h#��r�J/�麆�;�����H;��()�z�<p|�%]��iݓ�;Ƶ��#�4��ɑsB�N#3 p�O`%����l}c۴	}Q��؜i��xn�����K�l�C�ڕa�r��agFpҤ�f��1̃%��p�|����E��Ī�>4)G������1K��\��\�<��A][;ං���Q�@��I}	N�y27t �_h'�2oܱ�iFY<��Z-�!O���$��j��J2Yy�MO����Uuگ�kñ��#J�,���e{��m���#���n��ǒ��]4�d�X�'ĳM�UQ��a�`�~茶L������k,�
Pk�f����9+/[mh.��h���8w��t��7�N��g��-F���|��>j�]cx**_�m�Vʦp(z_ҁ�ɍ?��=D��F�rߘ�j�u6�j%F�{gu��~�u��R��dCߐ�/�[]n�F�7zIF�ܷތ_�ݑ�Jys]�F��/�y�^�*�`s�Q�l��1I��iӤ6"��"rw��%El��Y��hhU���ʙcu�綎+���ꪼ)��ӳ&�.ТhG�b/qڴ���ck6��[��('(R7R�ڐ��+��:n9��լ��Ch@a�ۛp}� n\)�jG�$��)��W{�
z\3��B\��i�� m���e�
:��w��0��0�1�k�B$3�:�"�VH��$xC����^�VpMpo��W���h�FEE�SV���R�=�B�+P~A�W_;P��+f�Vǧ�[I���B���l :)�1�]|8��BZC5�/� նD�:�'x��YN��Q���q^���@Al-��z�͐r9�o��M���N�A]��^���K�M���3��_���m>�[ϠI�¶�!Dp�?
�(�v )�$�����ˊ�eI:���f�'�Ìk��fb��m����1��U��F�ء�Ӡ4K���^�	#�bQ��g�7a�.�T�Q�X�r���+�{�k�F'� ^��:鷠����w�/ƴ��v�^���&Q��M�
�u����f�W��i�Wv0�4u=c�����	�5CZ�PN����֪��:riI�
_��N�YR�B�G���τى����{7��5�ƴ�Y+<��Ѭ���͸��s���5�ޡ2�m5�l>Z0[9�b1m�����lBsit$�Nۑd���U@�!޹)�ŧ��?>�$��XKM�O��sSNP['��u�ʐ���L��~ Z�r��
 �󊒧r���H�t����7�o�!pL/�~���'�ͳ�.8����N]�
�P��ꤵ3oh[g`���֪t�S_����|�xS���H~��{�S�܊k����$�X�-��Ŗ�������|IhYҰ{1dsEv���L�ڢ���g�¤�s�/�M�=-Z�zF++3k �(��u�v�S~�J
�!��kn�|��z_t�s͝+@�8�ņ�����E���&H�� �g��Q	q#�LI�O�Q��5F��^��<�V8Pt��Z���-���)��B�g��(���m!A	�����qhqZ�
1���5��p)쾫����u�g*#�cu�Ĩ)���n9�3B"��ʌs�CI�X.T�8L#f��ZI��^��Za�y1���'X�v_����ԛPS�����T6R1lN%��|�)�(
z{��O�5�C�pWћ-K���������Dp���4��C������;����R�7:�����xǑ���8W�+�(k��Sw�%��t�8�`E����1
̋�����k]�eçw6�9F��q�є�
�m7G�ow�-"�^|%v���Į7�ߦ���=�,(����4��@��~g&, :#;�e�l������3�Y����ڋ�{�b-$]�z5��m��)`0'�^?����b����Uݔk�t5��p�?��&ً��ʣM�n.s=ӧ̡��̈́..�15!�J�96!�z�9���0�p��v?M��Q���j�P����`D�,0�1�1�H*�hH�xzf������a�����҇X$���28������v�L����m����@�ƺ�+V.�5�֡� �qEZt��(�=Z�Q��j��1u8B1X�9���+:�ǵ6����0��{�i��.F�4�:���Z�ݭ��Ot7wB4A�dQp��J��K�R`c���2 .��|�^ؗ-�IVh�	"G�x;1j@�{3���}�׍�A�nzZ{	h@��� J�YƞCW�0�^q�NV��QI�F�C�ƾ��E�(�ys(���G�zN�CG���oaS�����W8�uKX
��Չ��}�D۵���(͆���߇J�|�OP�HU+ںͳ�z�+d�����jg5����'����j�^�8Ƅ�}� hw�!�P�!�k���1�:�&nR���=��@���?�;�~�X@����Ϯ$~J��`��P�����׳'���m���]m�FI.�����_ɇ�$0���қ�Z��U1��N����yJ��tFg3��ٯ7I� �̒8%��S �T� O� �H���$�7D~D֟� �����ӌ����95&������GՖО(����P����f؀�`�ұ��n�e\�i����;f�]R�m�oD������3i4��%�Q��o�U��I���Պ����9���mUڣ|X�N��`ø��P������ ���7$T���7�(���1$��ܫ�J�h�A3�������r=��n`�s�#���I����a�(Z�4i��(zh��~��D7n&���*�U�{���܉|YgI�^�ƽ9�<��/��OZ�][Kj��F<�m�~���'��U误'w�5��y�j���_!ms�!1��]F	��v\������m@�e������=6�tԉ��Q@��7vM��>�?Nr���>}�K�$VU�(_u+<�D7�>N��K���]�GgOrg������h[Y�Tx྾ǥcE:_!>������`���D�=����h��'���q_�e��4�^�3ޭ=~�!����&k�2��P��.퐑5Ro>�P���]֛�e�9�u辄-���m's��@��LnM�	@�b�w?#w��N�"���J_^��=�����}��57=���_��U�p��]|Hc	�,�s�T��"��J�W̛,^����:�p�����p�z���u�l0W��)��]�ݩ�d�f>����*��(�D)�b1E���L�=)U�V�L"ܡ���#��.��P�y�ry�.1>�����W�R�=3�\B�FQʤ�|f�|������Ę������g��g�9�H���Y-��q�􍆕�&�D�&�$ ���i�(^������UT+�$�[�8��j��e��l��hӿh�������6_���a�S�;�����EpJ�w����&m�[�лs��圜�Q�a_z)��9��	�zM� �-vE��d��zC�~z�����+GG�3=�u�vK���}�ʷ"�YA==�1�G����?�I��~v�h}ZX�<�{� �:�.Br�$��9��;�|)u�6���\}��\^.��۷�ܲ�	��)��x�Y`��$9�X	��:�T
!��0�}ե���ż@J*�APm�ϱ���[L�� �c�S"R�L�}�N�=�}3J[�'&�}�������$VC�2�R{�£��]��u+	=	�E�,���.�
���*	v�,�FR���x)$�.�k����������F��i��B�b9� ptQ�����F,�,}STG�:�k��9پ��b����
П�'�>5D��iZ,�D����7��ɪ��f)�$��'��"eM����+����T�1R��.�`}��'�Z���4�<yOY3{$���a�l25qRݜ�����U��O2II��˨HuҧI0��㾥A~�yQR���Uv��ɤ�Ǒ����u�Ԁ����y�Γ�B���+L��x+��:�JE3����>ݵJ�?��V
�����%�ƛ�Q��[�x�>N4rD���R�q��&9���!���;�冮�1��i.���M[$�;��M<[�7кwK jZ�D4Aؗ� �Z�_;6����t�i$O��������c�a�PJ&��`$$ ���=�l�D~����CkZ���RW<��<��?�X��D��x���#=�b9ο�7���b����s���x{�ٯh);Ҏ]�eoY�"�������0g�P��p�/�G6�%���-B��u'V�/���kIP���A7ρ�zE�����i�`�T�4���������O��KX *�B�݄����%̩�5B܋�f��W��ψ�B�r,7:MjRq?X��n��
��fR�	v��&��*)	MN�:|)�
,�aH�a� 0ͤ�o��+��Z�����$#�)�2��u��][����Vc��<]�4c�<�qj |�B�6�0�ˊٞ��+�շ�����V�c�}6�" Fnh���d.��f59LfǊ�J���US�	�Υ����*�3�u��d�0����
�#p��:No�2�Oх΍�� �o�6d0]�����0I	��F��H�6I��8�E�������������8[�[g�t��e��>� �����'�Py��!��
"5f)�;:ޓn�Y��E�l�g���x�gEu���dR�b��Ǉ+%��Ԉ$����<w��ג6�D�����󯇚X�U�Hb%=fz�䨭��*L����-b�ѺD;�U�����胨c۷uQE��dN�	
[�1�M.�jX���	���]ʩ�c��^h?�[d�m�}��r�`�ac8��������O�Qa�卲��� |�����Q����ֽ4��S鎆6�#{cu�!�Kb��&��m�
��!�pv�Mo'�L���?P�sE�C� S鞲�������(gxG�t��{ͩ
��y0?]�����?Q�����eЅ�O8��H��a����1��6�������>nP� x�` �B��K��Q"���;�l3$�C��߇z�DP?%�A���~�#���Ë���(����g�+�/�1a�)s�L��*���S^��t��=��㙂D�P�f5n�#3y��Я�Qj�`���x�� ű�C�:���S�M�LF;����w�t117sei�D�ڂ>�-f$��eK�J`\��^��]����)@Ѕ��S�mi��'Omw,K��0i�򠖡,�_١��v��UnL�N��Eb]h�ASX#bD1v��x�0����������Ub�Pk��B={��_���<�b�h�B�@��t#���h�mxKҷ�3Q��h1�5c������=��5��أgn
w�׷c���K�W3�tZ�2�_5<�$��`�� Yo��:�g#3A���`���l�M�J�t�=`�-��|�v�[���#��ߜ���w��
���W2sP�&�����z2U*_ZVo`	�@������Gy��o�8�����R�r턴�����:�ݡ����#W`��Ɍu���f�2ގ�o���X�vx���|�����V���mN������ɈNȱp�p�:@���l�6_5@ǖѷw��Ҫn;��\��h75�<�{��*�%�;ڍ
�%�!7�v0��`uk#fА���1�1�N\�<g�J9��{~G�����Є��uE��"#r���~� ��H����V7�g1�ܢ��l4��;/�l��Q�n#��� s��:�[l(p�'K{�cL��(*�l1v�R� o)�{U�H޹Ěc-�YTV}�Ǉ��O(��8����;����'�dB`��a���H���3��~�ix2BN��;�븂����9X>����s`p{�G�i��2pVFȱY�ùxP���D�V���ѓ����l�={�'�����3�.�
�m!6�;ʥ(5Ӝw-s4絢�s:S�U/YsU��le�-�ɓ<%�6;�y���:a��#�KU���,t�G<�|=����uu�6��� ���<�"k2�nA�k?٠�������brR�F��2Ƌ��� �XYJ�%��,%>�Aw�Y�K����u�G+f�;�@�=�RQ��i�˙�xU��f�b���.���\߈C�q���������A�!M����c>��b%�VA�S[l��p���������0�3�\gݤ�"��ZLt6G�ɞU ���O�
?�!��Т�������Cc+V�[�;���M��'jM�r�=�m�.G,�� B7�!��.�B�&�K�I�s:\�<	�^/��1D*����\y[{�|�.���%Y��u�'�\�>
�RP{�?S� �|ɛ�?��c�Om���3)�>E!�~�ι��IƤ�ڦ
����1G$�G����fs�\'���o�q��0�R�X��߬�q�!;�)C�@j��!n�,t��3�\N��=0	s�KD�W���2_��u���~���+�X�`����;��h@�s���G�5��>"E�_L!_Ls1>���/0��.��C$����8��yM���
�F�16��S����?�����@�,��]�kAV�Ϊ�6�ٝ�{%Yuv^����qƺ�<%joO%Ѡ
Jy�[���܆^bk
�48B:�����U=��EĔ�5-�� �e��9Qc������f���b�(k�5E�+fx�%����G˽�w��. ^���O~
d�թ{�x ן��ߒa��9b�i�ǰB��S� C�jG��7���l�R���>�����-aȵt��'�=���~b�9��8�@y��4o��{�ȶJ���O����R��>�{���}Aj��NT�#�m�;��H�9��Y@�:���b�zc��v���W��<}�O[i�s.��ʙeE�y)��mp�[�ZІr�D ���i;�ٛL�[�6xx�*Yel�S��������c,������4���W��÷��rB�~܏�-�uH^_�.�%��j��+��M�T��������]�S��9�k|�.�����'�~y����m�M���?w��~�l��xщEM� �LxHZ��!��8P����M�~�:n� S���w
�׹>� ���ۉ,:2�hw�
Uh?~�զF1.��Aq��ݢ���I5���m�q5��@�Ԫ��v�c��Z#�pasW���\-�@ۙ���ˑxә�I�-����#m�SWk�
�|�����ncs{I�����%�`�[���M�P9�.4 �*�"AS@�����������Q��<�����Aa��X�:N�Y{����$7��X����9�)hnr�3x��B�Eʸ�>��3�	�y�!^�0�SEA�����[p�wl�`���u�е�k����"w���j�e��� �b���c>�c�Sbi�g!ݳ����A��/�����v����,d����cCݪ��D{�gW���{��M�/C@F�kwr <��Hί��X�9�NUr��[�Q�)1J¬�q��|v� 
t�v�{�2ȏq��Xvu��!6�0�Ӵe�P� �Ο6�TH��)q�zCk=��������&��7i����:a��-���V�-�Y`4���O5��$����g��Y�A�~�ꬸ?��Q[�ъ66B�RM"��(.tUU�O��4�u�-H��{��1��}g�ׂu��ˀfw�+|-Q,L�!��Y�	iUF:xݤ�B���|s��Tbe��o���Y(��/5������ e�#ө]nO�4�=)�À�MZVn���d�V$��s>o$��1&�V5�o����i���z�9KLM?���T[�XK?~b*�xn��Xط�����j�&�t��3Q����R��s
�m�'IG�h�-V����Q��	�U3��P���4��
��n�M�Hw"����=��_�w��'�ʳb�;�|�lݮ��5��<Zk~��^�e��*�^���턏E�脛�����Y��r���~������EM!Oʀÿgp�x���ˬ~M��Q=�(	���ׅ�ƾ1L"���f���p�v[�mL�������3K2�UU���ιC��`q{�`-Iy��c���g�q�ao>��Q_�F+�*]�s���<�4����vh��Ϣ{[F�� �
L����Eh�C�Ϝ��%ɟ�<��g�u�����8=�4�s�Y�߅��*�_�W�ߏ�I������d����G���D�)X�������b�j�J���vr�DA	��W�sfH-���(d=�˟�.',V(��8��nx��9t&�Dʦ��C�k���v���Y5L���� b`���ղ-3H-	�\y�Ŭ"�E�Z���n�);W�x�`0��~$n�������6�.}V�1���
x�O�/0��_�9�H�p�2�*e8q�ɧ�BK��Ɯ�H�
�h�_o�~<��vu1U����Ē�z��9T)vA����։V�äe=I>-b�5�N��R3
i�H� ~(��d�	���`?.��z��e�% �P��a�^��%a��;�H�籵N����H����ُ��댇�q���SJ	��%�Oȕ�z�&,�v�5��t����@���$1<U,������?|J�Vֲ�JiZx�������<�Ȧ옡z_I�D������$��n]w�\�Z�E��:Ps�!'�C�G����\�,�If��S�x�3cD��\� ����6UR�2Ag:�<��1`%�60��mE+�a0��m>�Od]�H�1���1��9A0�k��.Qq3��v ��8�xL\��+���GY� @������#Q�A���;�g��>�T��	����ɧwp\���A�඙���#�@^��k)�6J�1�Í0?	��1Xb_:��'	.���&9�ަ¿�l��Z��E�aW�at�0;��<S��*�<�����yz���E�qDj�&.���I�XY	��:�M�G�d"%���3���l�7���<��S%6�Ѡ=�����ef?��Tb���(�h�N]��m�$��@k%��%r�3f{[|�,���[�A�$�{C��6����h$K��r 0g��3H�=��E�y��K	L:~`��T1B54#i�~�9��w&�^7m�8���A?��9��f�=�굡0�|�����@~�+jZŽH ���l�CAW���{��9�ζ�֣��Ԭw��!0��2��O{���/���Wb}N�7�1�����Ϸ�eU�� �7�!n"ޅ@s$�y[ѱ~�,^*K�%:C�j��K�� (�uB�Wd���1+	ͪ��R\Z:��-=yp]|ӏ��[_��0�����o�E�*(����p��~���g��42�F	��8\򿠇%fՑqҔ/��LB\ĉ@0:v�=��|� �[���[r���jE�ms��J5�)l-����D�2ˠ���P���p�ї.�/~���d��@jΒe���������'��8N�Al�ۇ|5�� sMo���c���a���\m��Jo?�{l("��yb�oUFl�ٵ0��[�Ŕ�BT������],c$Ub���
Q��T�@S��k���K>����ݧ_6�9�1���|�[�V�::���u$!͏�wPX��eH�\��ҖJuPt^m{�g�5�/! 
ts}'ł
�߆����|���B��j�#���ߝ=�L@��q�Df��XI5��x��ၫU�(4� p#ɠ��'�z���XBDՀ��(����qt~���u�`w��y���>-9f	 ���#+p��.��*������JA*mP���w_��tT}-��>�I�V��9v÷M/iO*(����q��V��|(��A��wU3�ΙP��k�Q0t$�'WW]��DL:�*�At&.�D��4f�²E�y�W�?�u,L�ErfD� �7���F�;/�@U��v&�|��rQz�!��Hm��E��B��#�hh�X2�F���� �J��.@�@j�����W=��c��O��ƆYO�!+���
S�Z����#�y+�q�Nb�Ks���f.*!�oҾD���![�	6�t�z��[�w�⌫s:�e0[�F�� ���~�:g��J%�z,��+Ź��~�C)j'*��D &�����#�˜k������r��qt���t0q�63'�
��� Ԑ�"oJ/F�!��]�$�M�FQ���OX�d�r��C��g�u����{E��FŁ�i���}�1-��i 8�bD=�m�T�Bey�:'s#$�
J�!��W/��f�)�gW��;��J���*��Ô6Whc���%��8�2�L[=�-<��C`ۙ��vc��`���2�rg2����X�̀í�@PL�`��QJ������%�8�O�2��C���ZI��7=r�HCG�Dz�dW6A��y�Vi�Y�,tFuf��ݐ3�O��+7X��YZ�l�zD)?��d�F� �+�U�!/��QG�=߸������l��O����-1��,._�.��^Tn �&���Q�N��:���͑�T�Y��j�܈2o`�Jȅ�+A��#~��iDF_Y�eDw/
$,��Ԕk���YV:w�	�h��B���-�pbF�����f���5@��E�@D3��4!��o;`�ѐ��d��"�$��JuEKA�����5\'�g��Q��}Nd�@���R� {6��fDK���jd����P�E�����rr4vO�z��\)��R�P,a}�����*:�f��:��n�o�)8@^0�4מּ�5�CҒ/�z�e��XأV��k����Q? )�eQ�9���Ҹh���X1���>�#�/V�a^OP���"��1�hH�M|�g���\K	�8�K% ��f��/�����CK����NQ�lM�F�G�zz�kğ�}^%$f'0��(̡��v�Øs��N�'�Z,��uVSJ��+-}��>��F6���<��������mMdi%�c3<j#�u*��#J#d""�#$��{�A�ަ�D�6f�8Z�'(���'���@��JE�V����|�aF4���gگ���Ǖ��*��������H�Ւ��dq�Pi�#����b)�ǚ3��H���OlO�AũS�`7�����X���^�%��n�]�P>D�G�_��5��(8�}n�
�iڸ(�M���z���(�?�o�`�X�5���x��6K.�����tJ+��yOr>�'Ey�	����.�rj�����\��jХ�+���^$(�r��O�rƨ} ���eh�v�͍�KW׉�#.��Zz?��W�Y%��	ǣ���x����t!��̲�+�@:�Ed;={_��/eՂ�t��v�Ą��o�3 �,�MfSqe�
l�������*{FO�9Ыw�2Y����0~"�P|T��(�[R�z�G%�M��zK�Y��W���LzO�G�s} ���ʩ�
��XJ՗�B�B�����{q��R��Fc̴yX��E���0B2**��2Z/��Lv۩?zz�g���������&)BS=�2C��f�<���b��|J<M/���,���vm@A�w��NN�b�
t߷�Av�֪�d����/b�!�r��Gn3NV�^��PK�A9{�y�']�өЂOE�`2���G8&4�Ud�)�����M�t��ئ�k��_H������h�زc�g&�Z���2��1}(]��i����Nmr�;k���syU�S?��\��_C�Q��	���E˱�� ��S�f�^hG,*��f�a*���(�](!��0Z5\��&��z�;���4��$�Vӧ��_��Hܚ�k�Ou�\ �8A�;�k�?�����9$����U�oG��� ~[�<:�MN�@U(Ǡ�@�?b�Auq~�龃�ʨ�V:yʎ�Cb�t�R���������1�ֺ0Eїz9�T@�	����U�gW&F*w�s}�#G~�
F�|`I���IKҽ�l�a�P����&f�ێG<�r��r���E���p�X�,* ���a�AEg��Z˟R�dҭƯD���b]Nn��Q�C�%���X�Tz����G�JP���	|�@b���V[�}y�\���T[�"%��y�����^5�G�I}��?�#jMz�x�AQ_�C$��QOZ�����m�C�ֱ4��#'}�\�E�\�MVKG=Kj��y@V��S��1-ɷ�ψ�^�c%����/�2[��Cu8kВ���q�K��ru)B7���:���׻6����s��\"��p�B��*!�1x!م{�y�z��k��Qީ�p�Nj����w�,�����@N�_y&j!8vh�?���PO�_�Wy� �t�¡��}ȊYiQ��v�R]o�G�Cl�\���T8P�C�ސZp	��ƞ�"Y�"�n���W��/Ot�$&}� ��6�B�aNZ������Q�n��=U��5�{М������ϾW�<�f+��n� �#��)*D���1a����R�m_�����*�L_�7F�Fj��ݼ[j�'�P��#�{=1��LW�;ly��5���9�_���
eB�}7-k8Z�����7g#��H��&�ß�Ɛcz���m*<P�Ңs�U�8�4�3O�*\��}��n�ݗf3Rr׈��j��rY����8E�.)��P�wnP>k�}�</`$ ���T�{`���#��5���Gu�X�����`�6X�oO������{&sZ�;BX�p�%]�*����X�;,�_#�c�{9�	��rqQ���]���L���GAkU���g��`?�qB�5s�^u[��
�1����L:k�k�f�럯bz���.Ip����D��'خE��p��Q��v1��
u��4��% ��=�����ZT���fC���Ӎ���	�j�>G/����W�f �WoȜy��i��
h�v 1(��׫�X:�ݚ�Q>�XD9xΣ �]מH3G��z�W=<҅,M�0p��ǌ�������S���5BP�yU�\��x��l�����΁�q�Z�ڢ!\_���̴ҷ���(�K��e�b�\���!��e�h���J@��'����yCGW�8� *}S�w�(ë���s�V@��r�ת�]����z��AY�5翕�n����Ds���w��X�#?��3͕Wy&+�[l��
�R�f�o��.�S1���~x7x��"�;G�kS��z�!Vɪ��tr��%C��;�'ϣ4;��l�J�E!��C�jt����벦�ȴt+9�L���5���%�HA;׊ �3]X���-�Iw���T-�Tn�i,�&tѽ}�K
U��d�4��1�e�)+/z�k�-H�
���I��@�ς�Z�4Ȕ Zԙ�9�p9ҒK;s��b^e�M`���g�?��x�!�Qdk\|:�|UK�>�y�C��:��V3�=�)���0/?~���%��E�cya�_�Z�T�/���#lVu��P�Օ��8�en�G��id��5dG
!Yq
�6ݳNx7L�5/��\��ƿ�3;��ِC�y��R��`^����V�G��A��$����I��������	R}�~vT��(�N��q�>M�@l6�1��r��Bg�7T��2򕂐���vM9�j9�r��3�bZ�f����W�}�zq9��zV����üJ�}W\��6o���(x����������y< C۶�
�w6��.׷zc���jo�ء�ű��i�����%������6l8�%�����Ua�>ҼK���$>>៲Ԃ�J~�+Q�s��'x.fèq� !F󄱜5<�����?������ۇ[�;϶�! ~X����>tc��IB�����"����+�lV�|4��ߜ��:CԿ��d�ʞ��˷�����ȷ��v:��RK^��H\ ��
#��-Y��U�BEM�g��D�C�{/b85�g�;�P�U�1Ԧ��oƟ����rO'�<��y�l4�W�d&�HUz�KFR�Ӥ_���c��"�)s���Zq����4aA˜Z24��HXw�����ł�:�b�1恹x��єa�xu��$�p���؎/Ї�5��l`�g�%��!ή���S�>�%$�m�{oa=�2�s��5�[@E���ڵ���/�7�v�E*�W�I�4���4��g���P �ޜ�sw�\�&��l4�m�˰�,龨A�R_�C��5ʤ�Dn��<"(XlKB�T�����R���rx��>��vP��X9;w���͢�z1M�VRT��s+[*�3[�N/2�z]ʹ|(q�*@B�;��2%��_x�r��B�Ztrmz�i����KDrP9rt�.<�ң��mA���I�����$�:���X�G0��x[�I*�@'fߐ�7�-9J��r5"�~1c��Bc�g�f9����
����j�S�]0h*K���O:ʧ��hn�EQ�
���3�^e�&���x�ʯ��E�f7ǉy��.��ώ�p�^��9���f^u����[��!�ˀ��9���ݯ)&W|��^�� ڦm�Ũ*5���@�����x�uLWZ)�NŲ|���hV��ocT�I����MԛX���yQR8'g����0<bU��+TLv�\q^c6"�6[v��͂�#�_6����dz�js*G�5���Y{�Wc�U!Zz��ֱ�ƌ�*��
���Z8\Īq�����//��<Tñ��NZ1甑��)��x�!��&�f1� ;"�1����P�5	�G�g댻9��0����<F�'n� �h�s&~�KBQ��3u�R�ϲ�3_I�Za_΁O��,�Y_>�=Md�c��'��Ӕ8#�RU�%�,Zq��Nc��:�z]Y�]����	F��[	�2�o����b��4K����E!r��)-[�a������7��`@����%-�_�_�b/�3jؕ�Q;�Sp��Ҍ���wG����V� ʙ���v79j{��nb#��q� � ��u�}E��J�72����CJ��rσ�����{�3��6��d5) �+7�ttK����k;���S �:}v��48@6���ѩ>��_���}�r��BX'�V[h�Ճu��h�Z=).X��+ݍ.)�unO 5���L�c������z�pE���%jK�կ�u�%�Z�ƀ��w)��ӄ(q5*�B�����?���������A&�[}٠�Ђ�G����D@�+d��h�o��7B�����5y��j �q���r������%�������t%�'z�9��#%] 0C%�"%%n��F�M�jW5��y�j��\��d�awX�|]s��s"[��L����_|o�s���|`1�$����u߳R���%͢��w ��!��r|���6�?A��`:��uH��T��78]ڥ�"�*I�m�����2�(��ʛL>�x��x�����}/
�m���]t�R	�As���Y&�(*��*�ih��|}�/�vr��e�� �Kb�ߺ���-��7ԏl��U	c��d����Y�*j���GD�K�}<�<����c�CpT`��'T�{+�:�Fg7��xd�XS�̳Lt,�'
Ӫ��P�oh��{��p	�l�,ȸ�[F_k�
\i�H�7���Y��d!y��O�c�C`��P��}6�9��͐������}2ix��AS⮻�>H�U�G�eB9�纁�H�n�1H�[�B���1������.rA0�^�eDK�EX�C/uV���@է��[:6���7������p+�����}e��$ڑ</�9������M����"�XV����:����yF<�1��BC�=�pGI�9^Aؼq���A@y6���7$�<��!�}/��J�ׅ=���t:�	
�Wj[���qj�6�tf��6k�e���F������A��濮X;-���C��D��I6��1
K��(�*��j�%���u����@�	H�$��k��[|��Uq�a%>�W��]���ɓ�^�W�^_��{X�`z�̲��"��]�c�K3�m�z�[���q�G�6���m��A��M��*6�-f�3��_�Mt�U7�`��N�������n�+�1�>W���uqAq˃p�%;�P��P��U���D����q>�����\Q($ag�w3Uq�dc�{���[ĳq|�m8���qW���O�k��o�Q�jT9���Mٷ鈥1cc��v�p/ū��R.�Fk[���b�/&[�������\�?5��4�Ӟ٫���;�1�������� �"}�ȊV���o`�K ���eT��:�2V�!�J���er8�RB�"圂�X��L�/Zi�}��pyl"^&X���>�9�!LŇ���i6Gmqp���H���o~͜�{n_�L3���0��'�� �h��|�����*	c���������ѵgX>���x-9`��,wiHB�ř����X���m����d2*K��������ꧪ�'[Ya@�Ĝ���>��[���})B:��K�K9�<�r���K].)^�K�w";�� >no��k�%�X�����l�}��,���k��g���J[�x�i��e��X6��H �A����RY��RZ�ˏe��95D���t��$�
��NPg�,�#���n���9f��&�l��䮦�b5o]��$�y��md�)XE������tk���Fw��z�eE�0��� ��N�!��n�ޖsy�ɑ����J�1ݑ�B��b0�)��?�ޭTmQ妸VH*�~�{�@����$��BoM_�+xj`�cY��1�楢B��D�!��2�r�pb��}wr���6?;�3f�yD��R@�Z_����ٯ�����#��'ꖝ�i�M�A�S� �(\fU��S��,���+c��S��7��扚Gjt\�艨���Qm��nE�d<O�uT��<9*��_�#6'e@�-�@y�����a���8���P��8r�-�W�bZRln�K��O'�%���p���̙'��
)�Bt�y��ِ���{�����_����E<�9ݒX�]��u�+��p���
#^���n-p����H7s��|~b6N��)�)w}����&��߫ړrN<^xC���/���l��w��O+9�M�3�8��d���X�c3Oi�U�H~�6~�1~ݨ).���x͇���&̦h�A������D�<؝Xe�'��YN�����]�ܻG���`�������2~nl;�;c���$�g�+��<c����߲�W(�5�Q��ݾ/{� �Q(�p�>'�)�%��۷j� ��1廜�����һ�,}�|!kH2�r)����N�b�O���D/���7[[��-2u����W%�j�1�d�yBƦ��N�< �&r���+B�+)UCŠ�&�HU[��v�7�>˹��b�.�XQ1j�w|���Z�޶7q�I�^�"��$a�fB�lK�+i�<�2p�[��u��l'��� a#��#�n���ߌc�a*Η�ù�� Y{�м���(9�f�:�.gܶAgD)�E���2[�ZG��خ�ވv�7Q��h��Pu���/%~О���[_w������p���4�,�I���(� �8�&ī�B�F}��8��J�D����G/�M[�\p�D}pOtb��~e�54w�v2F�H<<V��4��%*�t��ur�nd' ���cz��)����u�5?���n�֙�5���lJ�ŹJ>��y��� �f�6��3AV�P��ڷ�����C����a��ts,�����b�O<�\�y�jl�89�Ɖ���SW	U7�N;A�u��u�Z��(|��= \��#ș��t��T'��]5��:������sN�������#ŗ0�����I)�������<E*S۱�M�Q�.hQzy/ű@Ȑ���~�x9۔d�H�S���%�4�3�����18��:q_�Z3԰��U[&`����}{���	�t�z�/5��a�J��M�Pb|�%ɀh��a�������'�J�U�=o����إL�*h������YO����)MP�K7�����c�HG��2�n ma���������u1*8%R��`�mx˞��7������q�G�Q��P�V���W	ǋ�r�9�C�n��x�MΜ^���LF�����z\ �[<��⛩�*�I&;��\��_�Vs�w�V3��aS�]�=(�������c`���J��Ie��`%�q�3���'Fj�2A:+�.�ͬ,�-��6PM�週�f7�ux䦗�x��/`pg`��~@3(�nUE\�-d���U^����!���W�.(zp�J�q�6rl7�0V�6p̩TQV!>`mzK�c-���!�	.@j=}�j��N.�4��<@�-uZ0��՟�f[���U�u�J��/�kls*F$��vR�\z����W��Wa���{Dʰ��9�7>^i�>l��G]�C!���\n��b��9<�R�[�
�΃�ߛ3fx
��<E�lWUF(��@ R��c�3������$h"t|hwFT��T;�&�(=���|���>���M��J�����fUN���Ԝe
�<�?���5��,��>�ꈄ_<��~�I�˱(��kW#<�'$ܐ�)�ՒR5���K:�A&�hT1RԠ�!�G3Ӿ�ǲ�kK�,�����Ghe
�}�t;kt�>i ���C���Oۑ�2�΅lئn�S�%��	�̛7��u@���
'v4RR�%�$.0g�B��S���]���D�AE���F��ϰ�C��^��� HﬨI�� �}$� �擧��EI��A+D�����g���,BS�-���sm�Ez���V<$hͷoe��ד��ɧ	�gfii�o���}ӝ�7���b�q|c�Xe��������E-�lt�B|�G�����+��v�T�Еsw ����#D�紷���#��²d1'�G�Ջ�=����:4V�>W�U��䝨Ro}?���w������۽n4P�B*k2u���+�/�K	�-RHWA?vܶ��Y���XS����"�f���x�H�JSBp������Κ3�hb��퀾RQT�Q�|��d,��DI<K'h#�BȘ��_�2e�ܕna�e�C-���V�[l%�W#�s�_��E������k��%ۋ�}ޯ�-XtC"��t�̧x*A�J�B�t��Փ}��۔�!�I�P]/��y2hL~`���zg��YMP`��'�O2]po���&��T.P����}|7�zl����T:p0 �������:W2`����?h2��'M>�2�z>VB�5tl��B��3`��C�2��	4��F�UE�p`W�%��ݖ�}�}0���?�AXOE͋%����H�tؠ
T��2t�>��o����T����7�����b���U�������jP }i�����"h����c��V���mu�{��lg��M�������w�����=�� ,c��ɑˇ�pd��m�O����)��]���:]�\JK�ūf�|����E��
~�+)�t��V9w$ˎ��vG˜�p Y���n���*?� ՒoJ"3M�O��9��P"d��e(l7�F�2�l��TVke�L�S���I�J>�*�5�� ��A��eL��OC@��'��`A�x8gZ��we]��F�]L�2���E��Дq�NG�f�,u����Eǧ�CF�*�����rH��7�:�6mr!����a�����	{8���34`�Y��R�����p~�[+���1�\/��=�Ǥ�"A�i����E����T�)V�D�8z:�;�+M��l%�d���20_k��j(H�S��~{�ϥ����e�g`�i>H�Y�\����}�;w�o6��g,qhAk�`$�̡��@äO[�$n`�N���]�Ǐ�*�+�I~د�Bv?#&���1���HܤՀf�d�|L�4+!�q��yX�h�L�)�zy��d��2#ͣ!W=L)��4�ը՛L F8�,��z<E(�c�$򁯐оz��}�@'D �#���ak��(�x;�kl'���@AV%����L W�<\fG؍���JQ����0�g�����Ϫ9b���nR����R��~@y�0Ũ̧FD3%TJ�֞԰$ر�7ՒnͣY�Q�G�0�
��>*��A|��]\����-���po�
�z�|�S���c9�"=�GL~��qr���1F;�/�N"��L�_S�}���>���JӞ�tZ>Kv/�G%�0!/�Vz�����T��WA�*��o�[fVŧ�j�4Tډ�C��F�C��i���|{�=�U���rM�M:[�R����W�_H��_�3P
���[� |���m6���Ԅ�!��������X!�o_����b�o	8��d+��q�n��˳�2K�ݹyЕ=)������Sh����h Gc�Jt��dR�wF]���/�Ve��g��ٱG_L��F�x>�Y�D�{�w/38�hyTǢ�5�>24��MC&!M��?���fC A�#$a�+v�@�}�U��QF�]��֩]�z�	�Z&l��N�����mf�P�O�G���*&D��*@H�{�h1�������PP�Ry4�Ԥҿ� �,�ВN��-|��(�z7t�w��L]��i������כ�*R��`55���2�u��
,\�	*�=Yئ�~��B���&"vZ��m"2I��I��pj7���{z�S�,|���/�}�V�U�Cv&�+�^~�A��_7��+7�[��,�֤9p��)eW2J�3y0�Y��%R�����A�vP�M�U���vH�p��0Y�G���I���!@���S���� �Ky3?�$d�H]��'m��@�A�����l� �~H&�G_�Tu�jP.��u5 ,H(ng�5"$r40�g�[YN���S���-�&�|�A�;�Nd�)�e�DD9xf�5�x�%l�F�Ƞbî�6W�t\ 8U(ч�wR�x�dK��q%� b5�A�l�6K��Е�\0��6h1+-]�@��E-�uj3@!���˝2�jۭ��S��ys��+�'P���m�b�_>x]&�f�%?�,Tb�l��(Z3�'izW�����1��-�msY��8��Z����BA�H��m}jx���\kT�ji��"#�R�;�"µ"X/=Y�oj���Ρi�m��m~=:5{�ɶ�i��ca�~>�,J�� �;0;@�jv1,S������At#s&}�.U��.e��w��>�G�T������]:v��o���ȟ[WD�-xE���OJ��{�7�LkBi���(#*I���v.�(�Uh�O�Z�'�M,M@��j�d�N�g�܌�I�"���!��� �RzŔ&���=�3�h�L�7$4.��3;~q��4W�Z�W��M�d��-;?ӊm��+�n+,��\�"ĠxT�\�7q۱x���0���OzxA�����3w*;<�@yMy�W�����dE�1E�#�~k�k܂/��7f�Q�q�l�M~�@�k�v��Ew�&�R���+V��y���(��t�B7�R���[�w���e[�k�'`f�/:$����K���*ګ.��I��` ��c�N�UI���6S��6���n��_R���T�xA��<����\�h~��_���a���,�ӯ�M{�g+�5n��3-h��+��ͺ������3Z1�-_��p�qT�|�<a?au�H�l�h����@�ŕ"	R�_8�px��`���l�p����]�R�y�Ѿe�G�V��n~��"��V;y�ɒ�?N�H���<�g��{۟M����f*li��^M '�)���A�d��3��E�^|���T=R��%�H@�M�5�h�i	Y)`�N��Tpzi��l���_$o^6��ұ�f��0 #�����P9����>c��6��:S��T��X�ʟ^"<�,>�j:ecu�l�!��F6�
Z�l�������y�g�J���O�(n�����|Iϔ_������eJ��9����P��Vͤ/N1��T���nA�=X�M0�rW�K`��L.&�Y*K��:��pI(_�]c~NF�S������tֽ�F��xA�ʞE.Ђ\
D�{�W��?���1�u�gO�T"]Y0#-�b>�?V��k����Bge�#�H�.%�4���p�b2�|p<¸Ns�gӟ
"���*�Yd��	
�g���z)��E������fI,U
U">�c�FɈ�F��n�Z����
B�z��C�eeh�A���'��)��;�}V�q��3$��'��à�~'p�d!5.*�~wЩe׷���˜eA��}폭�\8�_������I �	���V���v����If���Xc�QU�]]��@���q��G;�T.?���O�[��׋[��E�>Yi?bт��Yfނgm컩1auO�S��BԌ����	���r6-�Num؏2r?T%o1p'�C���,ԏ��y���������'P�����-ĠB��B &�Rj(9�m�������p�}i+���C	��9�����.�bӇ(��=ch����������lr���|ҿM���Y�>�=xZn46&?/�KY������B��B���zAoM���t��P������T(C���0NՀ�/�SY-GV��s=LI�՚L2!����%;쑩2�1����G����8̓G0�F����)��J u�J\�a�NPh+�`k�D]�mn�L1�\!a|��ZO�y�uj`7��D0ڹ�,�riP9��p��Y|��
�nYr߼b����`T���������`�ֻd#�c�-	ԭy����������7H��~T�1��V:�1=s��M;U7�7�&���/{�I��F� ���c;�·O݈����?�y�$�%�t��k�)�Djc��C�ґ������mG�:@!M��j�4X��-�D��1���:����?���5 #Y�L�C�02��Q�-�oǴI�F���	�2p�)z�є���P�����)h��'4���������;xkx��Ou�L�U+������ԓ�3v%�h��p�e{Ѩ�0��ZW��.3��V���#{WQ��J�2������IQ�d��
g2LkҺ �0��'�X�" %-[s ,��O�.�j��l�ǭ!��3H���i�W�hڃ���nJ�QU���p����+��$,����-P����܄q����k�V���F�1�C�Q�y����#�Dy�M`��~�4O%٫�����\��}��������f*�I �ePj�Tɼ�CKX�qCC�߅4fI֝�<K���[�zd@r�	���T{\��Զݮ�M���|��k���9�p�A���v>^�;zI�5��Ԏ��f� ��Y�\t�0�{	7� "���P��U*��'��*���n��OYǴGR�2�p�R�0�l�����{�ru���#��+�K��ma�e?C�P�3�,R ���x�7(u�B���xW�k�A���)cOG<42���G�5_�o�
]�F���;��(Qk7�8a�{���^���c�E~�ʖ�b��'_Jd^>*}���>j����z�dw!���~r��������R�.���7C H��q�/������ʙ�;�.��_RƉ~�g��z4r��]�i���5�D+��؇i�Q��L(���g�=�N|�{B>(�^��9N����߰9�8I_��-�	]	�OK������>h�� �>X���vW��9�����7�!7�	WE�Uu�<��m�U����S6z��E���#��N֛\�6�{ن�z�|G�#od�ʭoIQe�M��-瞝@ʮ\�ċ�Nqs����N��z"����pƞ�LJs����g���7h��@+ʬ�I�����(j�z��W�����j(�0'�%�y'�e5:{���k�B�cÆh(L���Wzw:���[��q�O5�lR�`����:��gq����U�m/x(�Y�DМvh��=�6�Ut��*?H:�\��L	m�>�����]���:� ��{��he�R��lH�u�E�M3��M�?�%���쫌���j)����d�ޗ��XT���NeOW=�8*L*	��Q��'w��N-��&�p�	�i����y��z�2W� $����y��vVN'�?wH� ���@��b�<�q��e��M�|�[�,S05�dTP���J8��6�[ɶG���[p��u."w�N?� 6o��:�?����i�.l�c{��V�	�,��G�(�ءq`������9�ή �U4T�x��@�)���T�[��O��n���9;4,�z�e|,/�8�՚��P?�c�D.AB���%```(vs�]L~=D�?��o�{յ�����F�
6�?U!k��}�F�u�[R@A�Gά�+�U�V��񵛩9�Y�췔e��2*����:"���V=�z�����2��ӕ�CFu��X@,ZGtSI�E��C�m��n`� �O��>Zr�g�y����� �ѯ\y�|,l� 	|�N|�,��b�T*A̵f�h�{�>\��֔��%��M����n��'�(ОU��G��NrV���AUR�^U���s�xe`��uOe�¿��t6���O�$\iMh+y$����K�t�Nh�s�'�i���?�^@֣��aФ]���0��L���h�����3���^^�F�][c�K��H;t>V�Dw���L0�I��s�]�,~&����5bW��t�[�?���c�<222���/
r�	:�7G���+���~$޷I��Kx��+q���萿���ѺU8Ğg���������[�$b����B+>������`<�$'���m���{{tX�[Ud ��d��Qϑ��h�J��mU;��x� �e����Iy�'��k����2c) �2E<j��]�|�&b�	�gKd�?2�>��7׹H7�\�������f8R��'7�`S��)�۩�����_'꒘�(;����Ks���I���$��n��YK@�ƩN�T��(��@1jK�]�6�w�����|��[�{߃�@yG�й\�Ї\�j������m\�T_EW2`h��tVv��`���k)�"�e|�H������)�>�*`���RY���,pE�M��h��j��m|�X��w����He�.7g:A���c�@����1gdr�ҥ���;���l�����ؤ+d��dLR�4�V�zD�<1�k��^='��xu �=-��a�a��D>��>`}�A��Q�ɋn�v�3#�0�$Q��E�?��A��ѰIs-Q����aJzw�9��h6�r��I��*��OR�		:믡�t��w�/�L�Ei͈��\��YX&>W���CYWo ��Њ��pP�3��f�>@º�n'���j�^�߳���s�A40@p����M,�_ɼ¢-�XQ'�*`K�ױ�gfOHw����$��M)�
�%��}$�	��m6d�<�+r�ga7���D?߬������s�Յ��&(/�<�x��1�����=�q�"�9c ����,����͗2hm����jl�D�7�\b���2��0���t�+�^�A���^�o�9aI�昪<�[��_�L�y,xx�$�@|!}w��_@x�;�Gp��n%����Y�O�J��W�����%"1�|j��j���tf�B���P��Ҧ�kB#_<�I�Hx�a�������nỏ;p���`����W��#�E�W���|��>�耓�����)q5�ѝ�."}�jy�}�� �-�̸i2"͖X��$�}پ���`�-k�/#D�4OX����q��As'��zLWj�Bo?J�k]�oZYr�]�.�N��F6.����M���X��1��fF�Ӽ�8 6�s��`�6��V�i�	͌�}�f������xd�>����S�T���إ��ڷ' K����ژ�yqk6$���Ml�~**N6�Df���1�		������R����f��-�b�^Z�b��EOa����O݉S������d���Կ\�P�V��� uA��B�	>�����=�b"3���`���Xه�x>�R��}��i!���Z?T�GD*޽�d���C���dԧ���
�>b���J�͠���x�)�@ c��Ҙ!�W �s�ଵƈm�e�Z�<��56%�p5��9%���:��׌3�P0޽z�~�0�����C�����
��έ��'�I�E�E����Zz��J�cA���g@���xX6�#U�Ơ�+�[_�9I���<f N�C����3O�̓������R���ǯ��Pz0{���j��>�v|դǻ��{7C�);�P���S^;Q����E����kƇ���Q���?�`�+~Z��	'Z�H�\�bčD?�}���<��!��:����~t�+�����J�W�$��n׾��(�̴��͞�+&ϥ�	J���z=ޙf�
���<����c�oaX��m�7[�w�و�ɺ��GW�^��`z{�*X��_m��Y��sHpw�}l*�\�뻀3�2��"�j�lʏ��՞�}�;�X-D�������2$�cn��`�����M���Y!��ҽ4��P�@�f���;�>"[7Z!����,D*���U���͉gV�$X�I1���R�a�h��l�D�Q�u��dy�
��e���ϨE��m �811P�&Jr����}h3�j�(���!ݗC]}xv�b��<���ւF����{.�wg�j`d� ���u�1f���+�����^�8y��:��t�k�p6P����8�2��z�c�����N!Eg_Gcf�~��f�v��+�P��i�$�
e���XW��p��gy�6H�N���|4��J�b��0�1F�^7��vC�X�<�i���b���Fݫk�����T��uM�?�q��h\��w@>��EN����	���T��\~�=ōV����!g;R�k���cլ�[��G�/���������gR:@*}[��i�x��>��?C�F����&DH��&�� }�� ^/�$��Z#i�,��c��������\�cN{#��9K�?�F�pxl���W�.��ȧ��V%��}<㺣W�,��?b��GH���v����8��3��4�d��Z����4���fMˀ]#���u�bL�Pd��x�.k���V�+���F^3�f	��t9 g��$�5>����m�Y�LJE"z�/�g��x�K'�����W�&���:�~������+�4��.+��;&���_+u���ZX�VmZ|�	*�0}�Ғ��j����WC�8�����ƆpF��5GAϑ܄>�c�NH.o��>�ֶń�#�����3�/8��[��x0�$�t,I�,�X
�0��a@�p���~�[i���h8���D?b��9U;p}�}�J'!�v�e�;��SLQ�V��j�梢��&[@D;78��Zx��@�𖺽2�>(=��3��t �s�_PP�
��b�P�{��~���"���Mԕ��0$A���V��'Q�(��?�@rį+��)��;%CG�*K㦄���ш���5�	9Mb���e�޵�:����X>Eg��p���.	���8R�<��:�J�*���O��!���MU�c,�!���p׶���HT���o�d�
P��E�O��ȃ7�.��'<[�@oL�,)*}g�g]��Z�Y��Q����ΐ):o�6���iu�j' 3x�� ��c��R�cC}!��ը�YӾ��}HI��ش�̧�`��+����0����!�5��H�e~�5Yr�E�v��M��ۨ1�|��?��|?����,\�S�Z�k
�+e��T}NU����]�-u��X�
��̙��+�C�X�&? �#u4����zx��2��nƉ�d.`�!As͜޳[A�tU��T-�|�Eޭt4�'"��U8���YsXZ�V�qT��r��C+�cl�Ҭ�����Nd�6�=��Κj�9��?�L�~S�V��T�F��M��W���x�����e!%,�G������)S��w���W��&hN��&�Q�l�3�c1S��JewH5
����EVH�M6Ɂ>����O��8���ؼ�x!���Fu�f�nd p��P�KTq�WY^1�@{jy�÷�m-QVdT ���n����J��J$�0�uٗ�� 'f�'��®��*� ?��:�3��,��}Bg8�4��M�<w��q�mܷ����l��ٕ"���p;����>`ҹ7ִm���W�v+uiX�n�5Զ5�q��s)�?y��eHY_���W��;^��F�Gu''P/�$��"����S��7ɳ@M��T%Z�Q+z���{��!^��$A�-�x�鋌(����K����ub���6�UnTWG����H?J*>0)����!u�y���	�t��#��%�������A�E�P皟0�(ƨ��7��)E�u�l�'ç��y'u�v}�_`"����
���J1�zjx�+K�&z�w�g��T�k�zŌB�Jf�#��m3�����:@�Sz���[��Vvm��D��ò������ų6+�$IP^g��qD�6���X���E!���e0�,��=��G����oKN��fq{���)Y(RK:ܶ�G��U�gz�ܡ	�;.�.6F���l
oA�m����}.���(�����𚪉�w¾�ip�x��M�ڬ�I$����v�f7�V[cPN^�ˣ46ƒ K�Ƭ��2&��(AQ�k���ʹG��>9Wb�z� ~Ioo`'u�!��
o�O��|��sV����ǵ�N�c�*V>�~8�=[ ��"l�3�I�ˡ��)b���'$~�R^�/SS����	�_[0�מ�8ud,:Ǜϓ+�?�Z!� LdTw���@Bx�ub#0�W2<�mT��O��`�9Y��|>Sv�h�'�D�G*Ap�aT�~��-�^;����+�}%�F��8*uBDuP@��-F��A���z	Ø�I�\�Ґ���\KjY ���'�X�0K_�F�� lYtTf��KY�dI�#���f* �o���b��B��N�ZI���F�ў�XA>�\C�����z��Yb��H1���*����_�&.��9Hk��+�Nq�%ݏ�szv����߽4y���}P �S�fz�Ne���l�$��s�5�&�H3�C���kya&U���蟻������5ڰ**����1j&n3xX������R�-;m�ǎ_��q�~K#�,�)N1f��:,B��')��rF�w<)��-B�7D��Fb���wi�2]��ŏ`|v��_��/�T6�t?��i]Ј^��x?�'���!���?�ӯ+��6���,|�8�4*�2�6pj����_5dē5�U"嘎����" O�?S�~L�{�k���&S3G"�ObR��#oծTϦ��\+�}���\��ْ+^&��쑧,�x�$e�Ӓ?�L�X�¤�<�n-��+1�V�Wv��]@�!��>�ҍ�kCG���(���ϛ�a-��a�T�3TUc�3_�Ɲ��;ƸB�;���ԝ�,��M���#nq��y�����#OY��`{V9E��W�b�c���,P�
	M��'�ЅNK*� cj�Be7�:y����>�Ԥ��gfO�&�=�]�Ν��<:G%�@NfԶ1�j��Xǁ���3
�I�|�OE(�ۂ�RU��^�2"�⤌P~?���>�H�v7�!�k Sȫ��HI������� �p<��8v�������@�,3'�w\XzeS��Jw�L�=�D��2w���c*�{����c=��{�o؊N03�RQ�8�)�,@�D=�Y�a���ʢ��y(	�6�k�@�gX4��?AaM�7pK���C��OA��3njtZɴ(�����xl(�MK!f�B0��_|�Of�S:�E�w���q���£���)U�u�*]��R����cCkq���Sm�2���	���� �T���dFh&E����p�,�K[�N2��{+���
�j�a����N�@6�Ct�
�������?Q@|�t���K���`2�b>�+�|��<��*YB &������gb�e�� ��2��9k0��$�_�D��q{��,��� ���{�@+M�ĝnk�/����?$n��9�w�����-��cy�Q�WX8N�&�T��cay����+��r
�WcI���[��=b_׀� �*)�(��[X����`$��B	Vv��A׆��CMbQ>�v���w��;/�S��=1p��I2�s�z\n��]��,�3���Fw4�.���]�ٻt��1� ��R~a������z�_~��KE��M� (8�A�.�)�j�5i���-�-�]#�CJ(�~Ȏ5��Zn�L����E5� �<-��f�K���u�B�:�eHԑ���8")�Q�� x�.}>z���v�XͦOQmMcT�yj�.�9h� 1T�m�<�_X~{�ֵKǗ'��o�Q�K��+�u7���3�<�F��>�>�v]�p|���}p��
�D�0�'tYJ��M�x��=&H���fƿ�\Gu�ԦdYbU�-���Ky�jca��E��@��roj+(9�n��O��F����n�����u���G��j�Mb�2��e�bM�����K>ώ�S��=!u�3#����y��f���i$�`7�4�X���X)x�ŶL����(�z0@y-F���c���x�� ���j4r7 ��,�a�B{��I�����/�LyM{�H�6At��<A��s*�g��v1PV}s�,,�;�l`6d��u˅��ci�\0bw��[��+7Q�z�"E(�g�t�z��:��w�L�%E8[��ϛ��4��j��=��r���X'8~N��R��q�ڼӱft}��������ܣ�&b��Ic���Y�9�$�s��h9�/�Ʀ#�F�z�hnr���^����e�d�Ǣ�w�9W����:�,a��!9�cq�I�#����N��p�*�_�;�GxQbؠ�(��$w�D쭮=SY:
ǧ=gE�ǃk�d�8-��'aYrހ�$��o�Cy��L�I�5a�0 �Ե�)	�6��Uqۑ������Z��9��WOT�V�7�G��!Bmtlr� ��z~�z�J�$$%qƔ{���Z�
�1kԲ>�w+0cS�>G)��� .D��j�o��Cp Qh$O^@�y:�]�(΋'Vn���f|� _�˽/˞�	�>O�c��m��,��ҵ��^e�J����u�O�$�g��y��8���l�@��~��p��3E(-i����sϒZ�jI�}�����5�N��I���=���R���9����6ĖΜ/d�j[:K��'���`��*EQZEm=��m'f����T�>b���'���P���L[��
��˵�U8��7*�R�9��ɳu��i�2����ͩV�Ȟ�1���w�dwH �$6��v:��R2+$W�m{�ZR�EH�7!��0<��?elx�ӟ}�׷�3�Q��=�o�F1�	JD򬏺�H���`����Y������fH��h�e��qG-�z�¥��"��^������)�<�I)�L���L�h��N�a�$�?�������)9����. ����'Y��[�:�7�{+���ort�?}
c|F�Y[����]�b���soBl�1�T�n�_�O�'»�0<��*���������\ZV� ?\\�Q��ʙ3��z-w�``ô7�����O��Qb����3�mR`f�2Y��l[��c�9?����{���מ��(5Y��ӐkលXYt:y����A7X�����WUb�h6�C����m,�DT��Ͱ�R�MU;$<��i���;N(��E�G[&%^�%�]��T��|d�G��)˩y�j��.^�=|3�lM�r8�wYA�|��:-�p��ɠn�.�����`��&Y8u���	��G��2�4)[�s�oz��x�uL��qj	���~Օ�(�5H��t�k�Ma�|"��GOl9�f<!^�`��j�ߝ��&�,+K��p��_=ms��n|��9+�ѡ�	��a���+ұ�O�5�
2X4�qֱ��2I�5�����=Ȗ>�9E���hI���Nz3tO���k�v��<���HK�X�W���O�f�,���(Ea�Fl<�+����5ټč�aW��Ӎ$ܞ����F�o�ߵ�6`� QP�nG3Z��vvg��<x���\�v]/��*��͐!B�P�_�?7>+����!|�#���B"��d���2�fj���2y0�tI�>!7G$�A����@��p�dE����Ⴄ�9�9�Z\X0r�yۘy�<J8G!i;A���{��
UH���g���TC����'�x�tz��#��Vq�������٢rT���²���\zx�+��Q���M�?��|��X+���z��v��{b���~�J�Fk���U�u� N�B��-ަ��9q��L�5Xz��/���<�T��������N�����8�(�ֈF�CD�_3���2��K(�;�[��,�p�L���,�dH��;4k��.My0�}d� �u��8:�aA�2�a�z(�}Aۣ��c?���bḇ�fL\���x��q�s�	�(K��Ѳ�;������P��6
���e��2G���t8��+!��H\����j;&uD�R���3��R�bA=ʨ�Y��$}�ͤ>I>��O�*q5@���N�TM��vT��=<��R��� ��zL���)|�����V�v����=ӉT]نj�;��b�g��b�i�ˏ�xh@[��l�gB��W	I	Y�
x�
�*&B��V�wҢ2��F��4����\�����r3�MK�r)G?F�@�@!U��I<�y�|�1��;�=��5�B���A�z~O_��/h@��!�K�C����~x�C]9�j�?�l�H��ܖ�t�=��O��{���L|�ݳx�#�ڒbX�ؕ�l�{������g�ƾ�m��׍d�����o�}Pq�O���4�l	�_3��Vx9	:
�p�1�g���p�f:���	��7���.l,��`��2�'�5��3�^	I;��Nяx�_,������\�D����/Y�ɏ���v� ��1�cߜ��O�_�L=1LZH��ꋋ,)3��wpv��0#Ȭ�=�&'�Y$K�����ƙ��dT%�Hw)3��j§��d-�$2
¡�0���4��C�n��"[@p���>�4Ǚ�+Fp���=��Sri��c��9���5kzO+9��-�7S����9�ݤs"m�;����l�y0��tz ��'���[�G�p��{-uR�����3�R�)6(���/9-��s,˺��{���+Ct��� ����3rX���l��K-f� �*#%����=��{��>��^�R�����}��3�o������e*Y�'�"�wE���B�lX����y^�����^���U�������%���e�[0?�;��[B��a����#�� 5Hb����g�I�����xx=W� 7R~J�X����:�.j����;������M+�D�X�5?�|��^��֭ݛm��:TŤ��i2 p9y`����7ׅ���m
�x���N�[�6��s.�y�nj�7�3��$��"�8щa]j�⍣i�*��R3�c�u:����a����a��M�/I{p��t?��2�Ns�������E�{9�@����Dz��	�-�T��	�%���o�zy!�Y-�2��z���"�k��J���w)f�+��x��$�ZW���1z�V��`���,/0mRN�p"�H�I,Q:��yj��)��^"+/ic\yQ�$� ��&Vx��r���,91C��uo��º�������a8�����N_!��It�V�m����	u>�Bj>��?#��@�T3����ۊ���W��(�DZ��`��p��՛>���f�@�
���/�e��w���
�'XK�hG�Ǹ9zQ�_NE} ����/.�!c=pf�{w0ze�%�"�79�?��@a�h{��b��o}�uԩ�둎�`�b���]�̨�kj/f"<��qL�����F���o۟��Xsj���g���U`Ē�2��;㩒��H�r'd��h3f�_X��f,e"R�yv��<LQ�"Q�Nr?R����N52���P�b��3�eg��1<�]$.���p����Ԑ�%e���xuQ�o2�t�	�7�����3`T�����"���>�	K*�B�qC+��]���()��XzL���pFq���M��!��r>տ��'�e����8��e8g������/���L��A/���B"�F��Xj�\@{5bx-`�VO�]그c F��>v掁W)B*��dn����t�Lho����5~� {��Jr�q\9��q���e��y�Q��&�4�T�"�`�ld��-gn��7���`)�.z�-�'\ea!�Xx8_�-0��S��A�$el�M��%��oTT%#��4��Sgޞ�� �B*� �l��Zo�ɤ��;�}��!��(u�l7�6?=-/����� B�
�"��+AF
��D�����7e*�����e��`unM?��B'D��8�.�Is�Ǖ�t�,�����B�Bq�<�f��M�6��Nj�B��+��������[z =�NSsz�YH.w�A�}��b{#�%���r� � ����+oR��C��G����\2�Y���A��0W63jq �����0�j0�0�_YN�iΕ�K�ґ��H#�u�s=�Ŏ�o�	�z������d%h~�� @�img!��v��6���:j��K���<���\����p�t�v�����:�[�v���4s�J��20BZa�=&���t�q"���fN��TC�>�����*�X0#��sD�k/!�N:(W�TR�Uy��c1��F�H��~a�������ȉY�'O�����Y���+��Cϙ���z��ITl���[���H�絤)5&	n>�A���������Y3U��<2aT6����	��m��������6i�z�1�k�!6V=)��e_�c!��,�ȷ�vi6y�W�R��@��2�(B���k|���@��9�Q<ćp�K2�����R�����'E��t�@��l�� ���c�<R�Q���%Իf��?��P7{�f�����F�J����	���=������J8�tcN���ú̑���DӴ�!Z���%�2ɬ��:⣡���w�~縶��]øֻE$������&\��X+'���0R��T5�f�~��G��K��nHFa=�B��5��0K�H������l؆W���6K7�TUf��w�'��΁�T���E'�LUCZ4�y�������
�q���G�u�N/�����: ������H�$�T
4w�Rv����́��|���<
�U�^����K��5~��4�VM&h������/��CA�1E�i�I񌝄��|�3ɞ��i �;�ظ�4
@\��Փp�z��ο���H�s%�T�a��X���7b��e��K��wG#e4&B��F˩t�׿O	��:]�~�'NW�]ykRϊ#����P���M�(���t��0�	�gB	ˣ�䙃���̫.e�m<�����|��u����͙Y7b�Tk�K�ɺ��{8������������6"�i.�)jʷ���urkc�/���\|�'8J&)*ɲ�@8�M��v�F�IT����f�)��i�M�O6���_J�k�3� #���xܰ��ބp��S���i	�?�g��Bq1�ntZ�P��61@�P]nO�դ���)��o���z�]l�.AМ�N!a�3΅"�g+��N�=h����L��փ kP)S��1Pמ.!J���Ry���4촪���=6M6Ҫ�b\G9wCf\#$�kf��L#��h-)�q��bBS�7�L l�CQtS�W1[Zc�	n�`z�N񋛘?���A<��
0d3ľ�M��f��,�J�/�S� ���>)`L�W��c���aK���VDc�&p�SH�J�ю�pvm��C�w'7���^�=y�I)��ɣ��TM۰i��O˞v#�nK,��*C+��x���Ӭ�\�{���� �1Y1߈�Bv��CVT�?+���j�P
�_�̯>���E�z�w�G爉�� �<��y��(7�gI�2���@��%c���z5w����O�R�|��	��;��NV���y�w�pR�~l�|�}��1wY����p�=l���)Qp$����ֳ�:T&K!@��Th,���i �TƯg��ur S������{������K��U�'��)r�YTVKDS9���Ł2<5�������!:CS���Z�s�ã�($ձ/�^VZ����繪���hn����m��>����ѹ�_?v��6��c���;M�Zb֍ϩ�����l 1��#�m���z���\�yǶ4�-_l�����ߋm*�kh���gf��Y1�Ɛ����MD��
�H��Z1�s��(��x�q�b�j��&qr��;.%ι�O��Ⱥ�U��ϸ-�\�f��B+�֒K|�>'���!��o���u݆@H�S�1������˛��'��K�X�n�䄲��~�
H(,�_�N���w��GP�� Ǳ��5_x)g+��'�
���[?�P�'����:�i��Ng��M\��f�ZˮZF�(��F՛���.��8!I�[m��#��#;6;")���c�%�j�"�H^�\�7�ﰀ��.c�T������7J
+q���x�0HL}x6�<`�苧�5ɇZ�o�Ω�@}׆�f��"&
q����&�O�8��>����\���p&]rV��
����E�T�*-�7'U�7j훣����_n��HD2o�����>�?�f �׹i6�VƼQ��{1ͻ��X��/U��$�e���(��J&�ss ���{�.�O�Z4=B���`�N�k�8�=��p�����PNI�[��LT!/(��o�䲿�8az�6̱B�  .cZ�=b�(��t��?J�j��9�M��#UD�T�Cs���s�oA��gJ�D:c��i�qF ��-IL�����������	t�j�rt�o��5���Ѿ��zH\��,��b'�"���_��kض2�}�e�+k���f�q��By�KH��ں�JH籀9/�=�-E��	F�2+�� �����9�	C!��Cb�U� ��k�jO�o]��R������ 8䴍�X������0D��y�Aw̔�����	(��u�Dܳ�9 S^�ؕJ~;�W:2?�34' 3~ܤk�/q�C�}ia+q�(�!��+w�h��O��<��̥�pAI����
��U�'5#�>��SB��G�m�.�+w�M 4��'%�#T����Gw�hKR�ᡳ�\���|
@s9�/�G=�ف��n��y�]�C5�$K����$� �@�t�p��}�nq���� ���9u��g�/G'�����ZFR�ɿvK�J�aV�U.w�.1�9GBf�����5��A��g<���q^V�����G���+.�*�K뜋hl�)��'}V1+��ڲ��p)���&���Ee�X0-���!����r�(ť<�_/��_��jt�(%vmf�$u����[d�T�l�Xh��0���y`���Z�$������Cĭ5�n�@|���q#�xV
��|�9���%�jy���D��7N��{|b����#2�vù]�Y�0
g�l[���hh�g^�~@��a^{���^H���V�����4|F��HO�S������@ʋUMg:���ef�D�.���N����e'�V���S���ul��T	����!a�]�c��2b;��&����h��m߻�P+����RYi�*�աF	�`��Z���$ثUd�bU�Z�l����)����4�P�k�阻����<�����mBy�%�L1=K_���_��Nl�|����=
��g[�.�&��+w���n��X�������A��īY>�(&��?:�O��o���%�{YA�6܎�q_�ko8�M�L�`"�g;
�m�@���OQ�qY���+�%���ٔ0�m��O໿�����4����4=�׍�l�4������Y�Su�B��TC����~S�*cu>}Ez�to�&)�bi�^�4����f��������D(r-@Ѐh>D�C�gxv�׹��Ы,/Q
d}�{�T~�ܹD����BXL.�!�Ĳm��k��G"�5�x���g�Wùf�9��xh�\M��5c�����j%6A��A�ٚb�(���vѫ��qmE�rϣ��ey���0}��1�h-��Kb��U7z}�����C���'��D�$��{6����Y2�o�Y���o�(V�"?�A�k�뷦��=�F���g^)���~�M����DPn�V{E�kl����vQI25�r�@��6��r�]��Ϣ~I����d.A�; |�����!��Ms���p���y�l������[�����-�E̎03�`��t9�KD��ܩ�!��1�va���S�D(͂�?'�m���B�C��nE�Wa،`�R�1?n�o�vC�ԯ^@,��#�v����8^K�z���E�ῷܷ�h=��r2$#���8W�Q�	kzR&��d���������lAf�#�M�M������|��D�9�L���t�E����M�\�l��i�m����UQ!۸����?��,����Q�E�Z_��OY2�����N�r|�V��D���~iT��Z������!�TR�"
y-}y:�'�n6�r�Ő���|�9�uUJ�����`�����	fz;˹��_q�_�(�'�[n�@5�}�_f9�Ź�f
MP*����ڦkL�J����#�␀䕫��Ca|�6r��G���Q�^>`��nb���c5�R�`���:��\�������]���R�-�fs���D*��p���k���fI�j�'��z6(�I�"�x�,��K���4>���	���v�,�I�f������3��ᔈ��t��2g �\�d���C��C������9�����G'�f�d�*�� �5��Y1�O���Y��\��kó�E�<T�b�i=���3g/��:�b�(�>��iF��P����u�����"�&JO�uܧ/�E�"�z{��%��<a��ХzeV��� �[�^�9c��w��g�<4S���j��]S���_A�(=lbU�б�	q=;�h�+�-���{�z��L�u���Ԍ����휊M
���־�
��(�+��:rD��Y��_;t���DQ�k��<{j.l�ɚ26��y1#�P��0�u�G�M�!w�:̩���2�C�V����
�c��[�9LS#�.��÷����2C���N���h��s���I~k�x�	[-�c��7򛙊g��=fg�D �ҭT��}�r��!OK"�L�O
��kPs��<]��^i4��~J��V����R���)�]E�E��Qq�V��>7�)�_���C���n�F�ng#Ƈ;ߕו����؇F�GE�����-�_�	/_p�|�K��n�JMj��9��S:(�,m�NJ�I���Q�I'.dGAPs-�/��OMr:��U��f�w	�-M�F��F�x˃7b�|so�댖)g�G��&!	�5c����S��� C�W�D@��灟z�m���4����C�-�>�ML,ǳҜ�=^W�(�<E���r	����!�d���]�0�wҥ���7ѹ�?���C}��^�*��(�{,�uD�N��2�H.�NU�*<D9!��e��&3�z�ԝp=�Hy��Y��U%��������B�n��E��<�RB�C��t��V�5v����G���Jzd�d��1�}X�jB#��zK���'Z�s~�@>�(�~b�y#ѱ)i(�ֽ$S�ݴ�v�W�CY5{)��������׏`<�+w�L���� � u��)t��p�7���ˬOru9�n$�ehZn�x���y���H?������'����t09�►b�Y���qM1�nz�B����|�6�E^1�A�࠷iP�n�18r���+n)' ��������#�5�Cy$%�G�$����˱�ߨt�]�`� k�m�hP�DX�C	/Jr���[X>�k�Q Ȭ�5�"r�l���C�rZx����mT\��(�9݉M�����{�ل��>���h?�0�t�v+K�7�F�t0'��
R=�YF�?���&Ǿ�ҿW�y����i"RS������),?d|o�ԟ��W,��g��+������Sxѕ�=p�D�72)8o��͜����Fq'B��v~�W]VTv��d�3~��Mנ5f(q��^1��v ��n�~��=�z�]��P�;�Ö:2�D��h�O�nz��Ts��΄��N��'`ZB���i�����{�E]��7�N������f6R� � 8o�Vn�7k������5t��z⁑G���X�'��M���l��1����oM��zrۗ�_�����]��ωU������n�b���t���G�t���S�M]\7��� �P�����(�f.u�{��w��;Q�-}/����F����EĊ��Zg(��F<��08��i��'���j	��\�$yvk�:���a�tJ��Y��]�j ��g�#�\$E�?��傋��x^���`�S��s��yka����s��6C;��J�Ӗ�sg����5ɛ<��|fHꑮq@!R���P�1^u��}�xP�����n���]�3��[�!��k������d�N�~��%�F�]�C
�%���Ot��r��&��w�O}�����+;�����k�f�_�8��ȲG�
8�"����^�E-�!�n� ��k�;v�*��k���|!ޜ��T�������-f@�����B.�֣�k �)��	���+�g�B�N;|?��|}��������NwC�$�={��:���s/j�'���}�1����
����W'y���u�j�WxGJ��A�b������/w9E�9���}�P#���R&��~>M���ڦ�ABs?�0ƒ�+�|�Mm�tB�VHJk+_��Y��e)��.Èa�I9�{���ߨ(5v�����W��-/��b�m�6����A�m��B[�3_�˟ћl�Km�\��u�������hy�=$Y2g��� J!�|M����*ЅnP���*x�܄G#�=`]s%y4�-���V1��ɿ{�����[��ʟ�5�H�_����|+�;�E-��gT���M��5�a+Rj��>�����~�l' vc���#h��/{ꭨ|�c�2�pG���%G4�QQA�ko�
����n���|����6�44�؜������El�f�͝�>�y��k<��6�kʞ�<��j8�48W�Fl��'/�(Lo�F�)w(ǊQC�@UE��~�S��ו]�7��'���N��0���R��RF�U���*�h$$���R;!1z|�Q����FW,��IƑW����-W�b�y.���p��LV~��&�{$���5GJGz!'W�&+�����*
��5�}��L����3}᳹%��ݕ k�0	%Ú�{��'�U
��q5j���e�4*s2��!*��^`��E/Ί�C�.�
���>��Ò�_Qx'`��F�>怶mJ�G���H��S�qF��+T2������v��g`q{�mK��V!��B*�$;Ա'/�s(PA���&����mU����5�
��ZT#H���.o�5�Ѷ�5v[M��GbR��i|�V�ω�,�jN���Oed# 
�ae>!d���d�Y+���Eq�~����(ٰ`����2�ӛ��dN6�_n�{�"G!T.]�� ��GwV��2��ʥ����V2�\m�f/$/��Z��G��ܜ9C��Q��'v�-��y��v�?�V#_���h%zC��h1�O��㵚�s4����^%��O<��&9Ta8a<�:����6Y����_�|���6�a�ڪ�\޷^N:�Tͳ�(@4Mׂ�k�m��s
h��i�G de$g���`F�eI�ɚ��l� ���r��^[�����R�]%�1����ux\~��td������k�ewz�zԿ|\���c^�Y�.��)�žI��!ߠ.q���_B���>称�5��9��F�F>k�Ncx�O_��lܥ������p�yFW�$P[݁h[�v'lg���S�(N�Uߺ����I���jȴ�=�&�֪��@r)��>�OF������NOS;n��M�y(��uw,v(��W�/I���KOe&Jj���T�vy��c"����q�Ҫ���<*PpH�\��<�-��L%�e��̪�w���LA���-���(���{�� �:�o[3L��X�v�Q��	;|��Wp/�\�`-������hv�E؅F�)j���������;�}�"i	=�@ ���lZn��q�x���Q�ɼ?H�9����e�b
<@Z�z:Q�~�3R�9$U��Eͭ�w�}qww	��� �4�b�X�''�Ĥ���V�>r�wco0+��&1�b����&��aN���kR�$�x���w����YZK�4S�u�2*���;��d̃��Mq���L��ń�,&I��f��/C?�ٕ$���@bo��D@Ҵ"CvԘ!ceod��n�<�<���D�wɄvr}�ڦ�BwF>"����L��ZJ���W��G����_�-�&oRu��uk5�������x�LQ�Pײ)�#��H8��ߦ���\ɋfk�デ[(W�Ov{��ő��tJ�GeuJ<�^o[@���52��o�x4|p�|U�{ץ��W8���k*�܊T��na�C�qf59T���bа����n[�A�]�H\M�s޸'�Қ_���@��y��E����y�f��V�ޚkͦh��zmV����=h��`� =��m~{To�ɩ5C���M2)�7��C
B�/�=}�D��X�@�|0@�Ȍ��;%@ʤ��w[�g,ŋ��y�l�[�I}�~�k6�����H�I[Y->홷FC��U��k.��y�t�y8[wEc��M��y>�Z ӛ���)��ׅ-͈p��Z�`��-�����Y�>n<�.��U��o�TG����Ȫ��.>�ixS޺�)qcnB#�k4�=��,���l��W��)b�t�'_�˿���LДz��"ܜu��W�>���9��δ��>V��Q�e�M�8�^G����-3詾J=j9F/�	;M���IwR���
�~T��T@��D�.�{it�z�fI��_���fcT�J�&�3QP��Dᳮ�C���O�+}�A公)#���1�K�Q�m��e\���EQRx�P�����[�_!�19W�5Dh�i%�p�m1|@�����u~O��j�~��a�*�����n9k��׊d���!(�*��-�J6ͨ,�&W�"|�MmG��/�|�O���=\c��7�
��{
�]�����zo
[u�a\.zv��;R]�����&�׈�V��#����x-��-Pд��A��bV��[֚�V�8ۊB��!�N,���ڀ���F�+��y
��E��/���'�)�J �	��!K�Ug	�i���t�����s�x8I��3Z���L����pC��4��5�'��_�D�|���60�xQÖ�S^�ד�H H鎳 "���{.K�w�[*{�R��$E��
������B2�Z�N@��^�U���8C��(��\8��A�ʠ�E��������?�/�Hj�2J(��UY�JWq,��hD(��RZ*K.?�Z� �C-�m�9�������Q�!�mB���s
!HEa����;�ۡ��֫w&}OÎ�! ���Oo(`�W}�mE��G�N��De6M�ٱ��9d��p���:*@���������,=1b���[K�����B�ǐ����_=0sj����F(7���_��79�=�(���@^���5k��$/�-=�Q�,|���e�j��L���ʽp�Pm��L`t�u��{�F-Vx7�7w�Gq�hu ���vO.�S�Ӊ|���h��I_\����1�J�,?nNj�,<�ٻ�eX)���ż1��B�uq��a4k���SnVćW�*�6��U���}M�42����$h�b�i�ӹ�cbీ��fNv3=ux�^�1�d�J1�64�mTZ�Ӵ%hjlr�0�#l�7�t~�9�G��.���n�t�]K��G���
i�Ѱz���Q��+����+�Đ ~6���U9��N�FQ�9MŅX�Ym���]�~z��_8l���%⳱A�eW�Mn�_�㒶R�>�J� !)�E��8g�_���B��O�7Lk��+�.1���NT�)Vk�$s־�T%l���	�vI�N�zQ~8�z�B�˿����g�Ĺ�2<7쿮@՛ɵß#�����24�ѯ�<=4�'����A���/"C������?ML4\�D�1S��'�l��6��U����Z��U������A>��f)�2q,��K����7��s� ����E9��ǯ�ky�	�!4�kx�E�K�7fQ���D�iR�}f��?z!�9,�����	U4��(�'�Y8mH1�7'������l'M�T_̳��+u��G�7�@:��ozBI�OMrVb���8�K��y�8��-:�sYN���nغʽ�ƹ
�7aegq��u���+dz?ˡI�����)��"z��1e}�A���\���*²��ZB=Á���I����p�����t�l��d^�B�@f�OyG�g,`_�zb�DI����!ID3��*��`�
�e�C�	B�u�3�@�����mN���Ób��;@_g`b���.���Fg�Z��8lܢ�H����Ս~��P��\U�Z��6�j��\�c1�h�
��8����b�<�-]�]��|vV�q�&iq��b�����ɡ�VCX_s����?�\�~�C�b���x:#��`�e\��\-ϲ�MA0*��Dr{2;�����M�r0M���ٞ��*eӑ"��T�y&�G��x��������U"�w��+����jCL=i��I�uU�-�0b����~���w�k����0�����C��z^��b���[!Q��]%�6�j9LTV���5Ჟ�׮�,8ԝ�O0�OS���Mz�!
Jݑ�dK5�9���eafD�������p�b���^�@����K�s�a{��K���+[���R�t� �A�+�X�,l��\V�8�(ܤ�\d����vȵ����<Z��ϧ�XE�&�<�(�ݴd����g�v�k��ЫK������s���u^������&f��7b��l1|���M܉�ĺ���}�H�%ŪH��E��h.�����I$��hmf���!��`~a^�8��@��,�(@:��+pN��:��`ar�3�ө<ţ�I��Y�����H��o%2�6CJ2Na��xɆ�>��W4I���j������a�5-�@������w���8�B��rt3A�c_@�N�$�!��Xg��������Ab��y���7����t��7��pU�ݓR�F��Nˑ�a`�<�>K}aLC�E�j���0�F����YhM� �����	��-B%�:��[���Xv�ǉqH�୫R��V��\p�`�6Cva S�9��z���.�W(�.�ϣ1޶��˱���scJ���6��F i��I쫿U���ޠ*~�p�ەo h��bq�l���i���B���c��bP�Հ0��Ll\�\�VK�-%n�j,G�v���#���w�{���ԈQ��X��Yи��a�lD���o��lmiv�y� /+q:fM�������:l����x��5�F���w>^�b;�YԬë��jz�;�nEe��M��zj�$0��Y.����g܈����Q�d���X��� �4��.^�ݙ����Լތv#�W�Lo�f]c	��vq@/X��6�M�f��лʬ�(�;W�=���fP��G)'nW^����q���h�7ԒU�����P#�0�;{�f�m���\ePv>�S�V��yl�FI%��m�0\%;��V��F3��޾R��Q��@>h��<�ԋGAL�/��P�"D�&���n���k,<	�Ƹ���(Rs�2e������O�h��9m�Lh;�z��At�pgQo[��6��K�u�EO+X�:�@'{yѸ1�wHǧH�s�v�)Bd��N;����$-���,�R���I��(a�%+��OR5;��A@�9}������c8��BiE�
d.�ƪA�����9i+D�s��䡙Y����
�H&􁧚
P��}�XV���L�}�bP"|�VU��{vէ�b89��{��V�>$�inir�]f��Nsӫ�/���}�OL��P������E�¢�V��ƞ�\erl�@_'Ҿ���K��V7���>{M��؞�A_�CP�`[��?�p�U��VKV���}�����h�m�!�1FKg	�+��$0օ�[T/Wp��R+���h�c��#r*3*p��HKI�_�����!��!���$�_�8���e⥫#V	�Q�ܘu�1ht7r�`h&����#��+]ϥ��n�*;���Kʐ�'(�j�S���8�;X�3X��6M�/hٖ�!�T9��H0�x���JI���[��^��$1Kf�/��?�f��U�vD�`�"?�'i��9�˧=�ͺ	��uS�Å鋸�p�I�s�X�[�����S+������QU��;�\+"tdEʛ/>I�k
4���4�c����~TF�8�.ٲ}f�k�7<*��B|�AΛ.^�)�c͆�pd�Ƭ�9�۪ ��YTn*ށ)oǟ�f�d����f���Cπ<�PMW�^����t���%%�^�7+�B�rU��k{˺xll�?a�� R�3"_�p�g��:�q�\����]�C�,��8� ��.s�iFm<�62��K��� >�w֎�K�JL�#�)Ivu���^;����b�1�Vn1v7Ek���*-��I�>4V6��h���b\A�4�p�����|���k3�BqX�Y�������M�H5�G�GN�I=]���ԯ˽M�˸(��磛��z2�[ϩ��2	���3���`�u��XF�5�D�٩�����G��G�7�yT�	;5á�XXπ }��r>Jm�,�`���25�����YYѹC��'��������]�`4Q���y��k��i�P�T����b����16���?�m.46�(�ۙ�S��k�s|�/�N8��`��Qp֦_�y֊u�-X4kϝ�š��*5MU��T(���t�/��!����G���A�#q^p�qB���<<7����2���� ���	<�sw�Û�o�܉�p	�/���E��U�� �Ro$�w��;N051��|C���\4ü7�H@���e�,w��u7d@����(!L��eVܮ�{=�ol��}���В���)�U�%�LGd�PY!#ؐ9���e^�Yi�³���ܷH��̷<�d�7�d�L����Bqj}B��ݍ��I�`/��xo�Բ���Ȝ�f���Ѵ��I ��A�9`B�|�0����D�l�#�T��=%��I�`2���扺��T{W�<e��^60�������辯Y���6�cW�y��fN�vL��-ef!�i�ݱ٦��aB
+�۽bv�8m$�r))CʄK�����m��O��Uп;��ǒ>DkxsC�2p1���T���Ͱo�ENl����2St�>�]0@�y)�`��9��!\uD鰟��������WϠyɁJ�x._�
U���xP��p���B�wOxץZ���u��C�W��D����{M<����~�C��U���E����*ސ^�e~�V�����ެ�`D�1��XC^����咗 P����Ϲ�� ͳ
���,y��w��t\�	te�j"�K���v#��{�T�[���z3�6��q�`W+���<���౾A��$B��6!`�Yb���͟
CE�Mč(�-�\�{�����u�b`��o�?��zo_SA(CMW�`�{��lK�ta�F�ǖ�ý���YK[��,и���q�b%^�Li��P�,VU ��z�pg�%�� 9./)jȧ���(�ft�5j?
E��ʍ��?���p,mfFs��nܦ�d�}}�Q��g�`9!�Q�?�M@G��Wq��#�!J�v'����2S�k'�@�$�`�<���oW�it�#�_9��].�?K��|��0��Bm���~/��Uͧ���g������I
��U�j�Iۣ���sf4�,�o�S��L]���������G/@n��b�⃈�k0S�����1Te٣;d��J�mI��VB�V�2�)�B֩��A!ҁ��M��P�v�:��,�G��{YK�O���rRs��1�eL:s�l�2pZ:%0�;p��XoU�g��b?���~oO-FѸ�����&4 ~٬��]��Q�䳁3[���[��%�������S���[�i� 0�TS��Y����P깏�;,/�-�I�z��)��A���Eّ�ᕮԟ���&`W�Y�e�rl<��.�Ak#����qq����e'���B�����6�C�p�0����~&=IV%Οv�I".]�<f��E�w�g||X�B����QiM�P�S��ߙE2u�,�[P�����h��}V�`��ZhOc�,:Y���8��V�ԟ�#:0\�����O�I0M��6��	dc�%��bk<��Y��?}K<������(��`�	�����9N��a�%ōeO���U��D��>�����ޜ&�!V>��l�a񬘞�J��7>7ڎ������h��AO���V��$�<pS(�w��k�� 2�H�YU(.1�i|���H�oD���芊�La)�ցLN�]���=�l����a�)���i.�,�s��j�~���3�k��
�x����,�*�a#��8�o����G��_VSm�V�����S"��<�s�'��<vm4z~��6M8�� U��qg��Vb����ҴF��rK*���A)�TjZ��3���G`j-A�l%:�j���V���e8���'6�U�$I�S}�<�b5l����P3����ۻ��T���Z��$G����%�܍i��6Z2��=�M3��c���)+j�ަF��#L?ogu�x�OB��c�\.>���'�=H���Յ]�f�6&!Tr�z�b|��T������Fv���XK+�o����T����h�Ul��N���7@�F�44
�p�2��}C2�Ę�B+Z�A/9\�7�E�%��PO��󂩁[qt�a���ׇ�s���*K���&�\4��F��/�G����G�WnS�-�.�6����N�'=�B���r�nfi��|=���?Lm�]𥳐o�ݧ�n��^���`;U�E,������~��f������UR���<#s&����kvi�m�A��zMg��k�k��z�MM��]����k�Z���*���jE�U���:rG0��zdB�\�qݫ�n_2��eԸ����(7Vlv��2St����7��	$*��7�#�ҏ�y��M����[�J��@�&g-�=�����wu~��ƧQ
v�SOJH)���	%J�3�L/IT���r�t�b&$LNo�I����������c4U�VorW䢚MCR᫕��|6̭�!��ؔ�'h,H:7���lA�l�x��?���?��{u����t���*;�h�}-릩�b��A���pO�d͑EY�Dq�]�X�٪]�b�� �(��.g��!�}�:d�����w2\lS1�ف�
�)���Xxy�b̀�~`�T �Ch[x��J�"铵�M� �c��X5�ש΍�+����i����q�Z�{.�r���7u?c"�[�'Pr��th�'��Rk=<�� �}T}.�r��0h��f5!A?Y��Ȓ_c	<C%�t����
��%���Ez[+��bX������ޠَ�wdf�}���ȫ�����H��"�b~�����{�y�Ȑ�������v}H-^�n2���FbU n
^�w�E�{�jTG[�\h���!G�)� ���4�[S�"1��"y0S����v����"6����(��Vq߇p����7vK&�e�_z�0CD�L�z�z�շ��읙+A������1h��Z��B��ot��օ�Ru�A���(I��2��~s*�Mea��,i�p���1h��]V�!MC�RI%E�kh�N��s�y��M"�~bd��w^c���9��^n�T/ݮ�s��OB6�s~�&n���LX�y/Ϻh������Ֆ+�	/v����<�2)�f���@��۱P���it�ۂ�2/��G7ifq����D+��������˧C�\ۤv���j��-�4"�E�Cv��W!�vO�����<0�f��7�+�;���v��XEF���}�{�ذ����~"���J���R����&>-Lj��ߝ��:0�5��t+�?p�Z9'����S}?�E����{E7f2ŭ����EFI�7�8epG>���G����od�	��z+7`@QB�8H���gw�H1I/�q"���а���6m���` 0=zn?.�5~_�&	�B.������47��h����w�j���������R$�y�Cp
3��j,]��˫,~��Fx�=�#�rS��v����� h[O:Fɣ:����'��y`X�%��|�8��f��?�i��;�:fk�֣�����P����>�h �jd���t�\�}����}��UMRS����H�OD����$ۼ�!x�������]8Oȧi�h�&1���962Zν���a�v�F�����Tf#&w�|3�΢�TbY`��<p��;'.����+�n�=���gN��=��(�Fk�7��"�\�(s�����vəut��F�����*�m���}2CVU��N�'���"�'��Y��Tb�o���Z�/�߂�.�[�q���'�b��"GH�%��Y����%JL�����#=�1�鉆Be��$1෗��$�_�H1��O�:Υ����;�R;��A�)5Q��<J���Mr{_2��R�oٖ��'R3^)���Iu0eM[P��
μ) ˪��!�p�J���~��;s[�
o��5(����49�b��h�2����D�Ds̄R�1���GW�H.Z�b�w��8YyW��n&�fعa]C��v)[���rK5<��XmKhW|v��}�����KB�!�?>�x@�.��BE�
B��Ǳ"��-Q��4��K�2���ؿ���rOYb����|�˺�/�n��ϖq*(��\1Dc2:7�̌���g!nT��	�Ąy�u=�o%I|o���,����J3_e6\T�[ ��Ђ�b��mǹf�c��߄T�N����U��i�z�s�U�y��5:��A�bЬ�B��o%��΂�ȈjGɭ�V;�$��	��*��Q9%G<�@g��._!JO�^v����7�$%�L+)�0)�o%�xH�"o:x�`�ѿ%i��=��[���1����� s��$�����;K�U@(׆��$��=���y��2^3��R��FŞ��Ɨ�'�n�X�1��MVBr�:��X�?�֤颃��ᶩx9�b7@*,4���:�&*g�!��:�~���	�۱,���(���Q�ڞg�9�[^�Q���_M�Q�1���?�D�{3T8������-E�����Y $��ִM��hҲ�јĶ�.�(��1�A @�8C�����X:�3#��ȅ���$W�t������o���m���>
�|K�J����U�}j����9c��P�DrВT�dyǹ �â�44ѿgR��A�w��qM'X����J���L���ɧ�]��Vyi̔��.7���ɟ�Q`���fU�~S��2]R
�Ir��ʪΎ�@��Jn6~�A�����UP��ԁ|��g?k�:����|7�<)�ָ<���U*:�Iu�Ȃ��|h�i����7��
 �����뇑8��r�	�s�G�t�*E�˯�gŤ��(2:ݖ�L\�M�.y���4����$�z��U
��I;@Z(�}�v���w��?�pK�f����T^� d�K!g�|"u����վx*?��h��-�#�	�Cm��	��5|�{�$Ռ�I����O@^w'��~Vs��(ײcZ�� �$�{�B�5�^��ح���>�s]A~��
E0K3;�C���.��SPƷ�ih�*Hp>���X�A}����r��x��x�p�i2������K9��/�g�DT��A#WQmY�o3���,�U���|$����Gt��(�� �AmT�H]�) �~��틅(�/?Ƽ��l7�`Ӭ0S�O��=n>
�`� n���y�l{��^��/.�W��%7���ݷ��m��d�3U�с��<�r��^Y��at6Ϧmwt�>�K���V����cB�S�6%����#�<U�m��#�&s�ǈ�dI�Di�-�vC
`i����+���TWc�D}��(��Z����2J-poRϏw�m����% N�8Үtp�IVߦM�����4 I7�b.w��gk~&�!;5��}-���N-N���אl������F �T�ͱ�D8��C�W�����Dze�e
5-懋�r����_r�/�	��C� ��� �."��Ϲ� 2�e�Ͷ�8��p0j����4���1�1v7MBOt��۫|����:�gűK��n媢j��9<�/��f��c�[bgnJ�M��g�|��-'7Zu�͸d��W����$^<>Y�3�R��0�1qӖ\Q�@�$�T���n�����G���a�L����{�aɼ�[�y1�B之��Rx�5������S(,�t~�fWw��N�<e��������Z*Ɲ���ĵ#��<��9́Q�3H��S�lO�ʈ�]�_����֩N��/:JE�AR�+F!r�}�EL����M�%瀾`.3��&�b8�.�3�f�8J�hA8����_�R�'�J_͙�f�{o����A�_�FI�Y��̔�)k$�TT����F��Pj��S6��m����{+g�b��\�u��V�A2Z��}䋒���0ڛ�j8]@	���La��+��S�T�J�q�Ɂv����{�X�r���~�����VD87AG��'���4�tix�,�U�2+��O�Rú�h�l��GT��3O{����q}O���sd0�5�og���+�7�����tP��&��c�7���qr׉9�2�qf��p�P�/7q��ҿT����B�"?�ٓ�_�yo;��m�e��[D������4,@���+�s I���zߣ&��z��V�"%���iz��`TQq��b����w6�!����p����&/!|�5dA9?��{��O�E�X#\��,��A!4�(��~W���f2�G��l3�w����W-)�FT��TY�5��G�@b#X)NLнPm�6�X����7�M�0jQ��_	�L�66���L��{�4��C�iS-�M�mQ�qr�<g���%A��,��\��������/魌X��v�bVĿ}'�ۯ($]IX�������Lx#��-�%��V&��˙����bY����v��S�=0�v��|V]�-F
G�W�΢�ԙb��֢�.����� �E�� V�V&���Bƀ��d�_�8���J���TT���6�$�\� ��D�ϥ��0/�&wvs������"f|�S�Y����]�/����R���]!KFPĤ����QK��LQ�=��!^Nל�z�ə��"t��R���ʺ~	}6����$��K �=��C*(>q��˱�[�|��M�o �d�_�\�SyZ��@���R�>�;#�W�0&�Y=�܉�Z��g�ge�`�3Y�]�pd����ɨs��/P��
�����Ϩ��;ۃu%)���j���M��h��Л\�p�\L!p������6��j�н�|=M��5��L����_�a�6v+���Oa����%�6��B�7�ĤPؿ��鞜����5�C��I�tE�;� �^�����S�nq��El��Q�JU&��)�̀���O�Uְ��â+ʊU��[�ǏF=��B)9�+�6w)��x$J
�Ǣ����y���s�8>ѓ=�A�s��8�eR�s�͖%wu��'�.��i�~�O�	|^�MTj�?͔ �|��.%[Z٨22��8�$ڱko����bq���/��ve[��`2�U�^�2�^ȧ��Q�	���c��L�zM@E_��rV���f���dT�c�$�}YOt�l���u>�ASu"�<�����'���,���" �j9�Om,79˕�&P���-F�Oy^�}l��_G�aV+��C���������)"kꎬ�� cߗ��ɨ�o�B�BөD�P�gcAw�E�0(���RV*������cY|��������_Wü�q����R��j�Q'����rLP@wn��/����E�ݝ-yi/t�b��u��O��G8�5 �l��O����t�I�@�y�yL|���]-�>Jf����U�^�PP7�]��+E�����sǕ���Q����,ƨ���m6k��nf�S�}�Z�^ �<n��F.5i�ZfEu�/�-�.���N�eM:OV����n���X��0&�����{n��3.	����`]+�:��h(q��@��^��akIG~S�/���c�����e�W��?R*�Nzh��9Ƙ�SǑ,�2\"��kE����-}f&y���9%�o]�Rk$���[�͌@R���٥�u��I���Ԭ�8h�X�Vp�v2�Q�T����F���̣8������8]�{<��d�%8�!||�i~p��DnԪƞ����H��h�?C��f��{Tb��,M�Z�sT9���3@�Q�G�R��k�a�Ha�j�z�L�^ /&Ld'�Ҥ��m^���mӷ]��X��}�@o�"*���������}R�N�ښ�`���� ���ٕ�dg�T�G�l<Y;JU�4cf�>ph�ܖ;��du2k�)A�����i����@���\L=�0Jt�9����
T�3����?1�^��rM�5ri3se%B}S�Ѐ6�ujս��8�Xs���1�/W��?��������q�lT�сU�Fr*�S6��e�HO�m�c��`��c�O�s��8d)��f
����:@+~���� �Q�-.����K���/a�)t*�t��^k-�ҷ %}�2���!���*�M��K6V�(>������{����Ə?6U�A����!gpJ7�1P�*�V_˚�7���qA���|�*&bhIW��vƟ�..g�C�,���Z��0b	1�������,�?/�da!sS��82=Q�*�1g-���=������=�<��=��Z��u2p��<|j5�Ũ�"sq��ʜ*n�w"zN'*pBJ�|�Ye�oU��c�������eڣ�(�<W[���z��^=�=��c̲�xw�>����"�u�Q%%�(���&LK���ZY���+F� ��}<�� N�^o���º��C�䏱G��$��W�ڄ�)J�Zu�����&��`���L���=[2�'hOI�*�>Z���(���<�R3�U��nmȯ��3��J�}�W��\~�rrzI�����^�5�g+PV���4< xME�*/���~�|"��ئ	�����G~qة,Q��E�i6?��^%���[?����>p��v�Ȟ���؃Tr�"`��Y����=��o��V-����>�.�q�`cn���eX���4A�BX���[�M����?R�5*�� �X���Z�e�.�˲��ղR�l:^	�?�Ug��G�Љ��US��s�gr��R�~xnYC���Dg��� 	�ʝ8�U(Z0
�#���^EFB]gL~���S���~HTQ7,z~A�kE��a�����gp����!t��jM��
�xP-�fm�S�5]�K��l�w��u�����k4N�Ħ�����|L/bi�`]�����4�X�B(A큕�;%�{Z��v�_���LA�s�8�1�G������b͝���㴦it�rhu�(f��T���#��������<�/s*�bƕB���`jB���k�eS(Ya)�t�I���Y��W��x?�*1��	_ʴR���2�sN�����d�5����vǰ�j=t��]�5�������.&b	I�^dꚋ��ҥ3[������:�a���f���1�XV�$0>�Z�*,�$�`E�(RǱO�v�x��=�1�;�Tiߤ�ȼ�HA^T3�7�okk]������OR=���ŵ��衂`i�|PX�/�d��m0_��]���wF��� ����;��N|�u��K�R�.�#���`���'���J�tRX#V'�3�7C�֔���'��Z��C���GLk��M�33�ר=����rIx9d��k�����z���_�ol\��)6pXV����tS\V�y"�'�>�ʳyAb��ꈪ�Tpƒ?{\/�|������#��sޞ�3R����t�}{z��1���ֆ�Z�[�Ԇ�89�Z��/\r/g��(L��f�N$U9�h�a��q`>uqӨ0·^^��}��-;\b�Qi�*��21�J}@�j�q�!a߿��)�;�4�YP
�!W�c~���Y�Xa��Y���#"��'+-gu�[L �i��.^*M���G7 �$6y�Q��w\`��#��u��2�8	W��x�E�,�\��O�d��AV�:>�9&Є��m�- l�9�!�"�*��(+��Պĥ6?��Όɏ���?y��Jp��:ŝ��vn����U�QJp� e�rn�*����| ���Pj�I���J:&��fm�=25
���ҡdǁ����,k4�hd��kLs! z��VJub"3)��6��� 0�jZ�����X��`X�?�s�*����T ����Τk��,x:�0Dl�薪�1 �d�Ó��"S���K0Z���k�z�#��7&~�P��(��+2��\G6^ח�Z4J��b	#W4@�t��F�B�h1<��U���2[�ig��Ui��J�����J\��0(��
��>7�[R�[ɯaY�����R88[��n�d�N�@�����-N������u16�&�!*	��|��z�6��k��7[z�10,=�5%��5�Tl=@�g2�k92�>�bC�כ����S<��^^��XK�|C��
������=��;��q�*�4O7�p\Qh�xÝM��A/!!���&��|��&��^`9Y%��ds�scw^^o�o�,���e�� ��Ū�@D�*������(1^b>3+x� �l��}o��[�CO`|���}��63�f�;D�* ���7D�ٿ/���CQk���4啱����`�X���D��K ��̹B{%_5s<��"XI�]DZ� %'�W���,�s>Q>R���'�Z�	�Ì#I'��T��V�����m�v]���C�hR�49zd~�{Q�8�N�L���!1a�޺��b�X¬��:3攗|q+B��,�2�D��?Q�h C�M��WCť�R�F����Ne�V�S�M���.3JCD�/W3��K�R+���`�F�R�<��,n/��؈��>2�Em�0H�6�3� w?�,�Os��֣�PT	r�ZL�#�&���G�Xf����E@B�x9��R��_�y�Q�cr_�qvP�����)�)l��J����K�����j�΀;��'$SiJ����ˉS�`k1���w�YM���MIV����*�^v!���I��AA��y ��]?�j�e�`��~~R����qC*G�焥m�(�@�b�����uA�����+�1����r�� �5�C�<�`�J/"��⾟���}"=�����u��y8 ��(��*+:(��NaK�����Y�k��R�[�g֐�y�썐晅��2��^�C�v�Ka�q8���iX�Sς�P��<�P|fi4��x��В%8f����w�ɭ/;�c��i5	�G�r���B]��@H�U��=�q���F9��P�OnV'� \ \pI��b?bK&i#�����Qk�4$|{��W��ܴ���F�D�`��7��m}�I��5�ъ�tϡ�,��m�(���lU�ou2���Rc�]�'#�z�{+�A`�[��J@ٌB��`ܵ̍��0*�*��*~1ǳ��aX�qxS������T�|"� z�j���,:�e���7[�Ҿ�h�Lt�� �A$1ȿ?A	�|���:{Z��?�_o�ii������,�ܻ�M�F��
��tO�nN�W���E;�4ڕ�4�aӼ�};|�%(7 � ���
*p�oub8���F���@��Hv/J�rkr��ֱ���t��C��!Ls�Er@�ݡ岺�4�Q#�=��Cm�j>�$n�F�^�@s��mEמV�̷l�'Q|2%���qi0��P{O|��"�	0vq������:�������+Wq��~��0�T���?��:�q��s���O=���LRBh��+�cDq�������A�/��x��	��95�fk���
 m(�DN�)%���#D�
P/���1��'H-�|X9_�����Yi��8c��F5���I�D[�Я�[[���~+��A�%���(�BM[)E+��
V��{�cz��#�����F�ܶ=�ͻ�A�����*��(��k�F`��of�s�,�A^�T���tAaq�fV���W �g�l<!F���ˮ�=��:]Ș!�>�l����F�r@�d۪�a�p�3If���+�� N�y`�u^ĉ�t~p���2G	�<���)�ݥs.��� 2C�*o^�,oZ2�8��4T�����)��:f9���o���R�}m�(����Q����65!�U�Q�E���s��oliǰM;�Ic���@لJ�:@�^����J䑪��T�g	og�- W%�"�<VC^��smx5O����nތP)��Ǻ�Hd��/��sJ��kb+`�M3
E���^e�r{Z7/�{������w�Ȭ7Y���|!(8λƐ]A�;��;G�\���RY�t���8ҿ�F%�Kf���m����)a��ٽ:�C��w�6��+T�Mt]����PyM3��IS��L����D}P��@x!`ln` ��ۍ�,n��1��ی���`�C4���;T��	��AG��a -��yC���4�����҉6O��>�7;/����I}]	�t����$dCJ�_���H>:F%�tGݔ�t��Xό��t3y���,쨳q�*S����@�b���ѣ�"�4����9��(��ܘKN����.�l�@�X'ZE̐�E'����nu�7
�~���V�	� ��V:�Ҟ����T���y¯�?o��c�u=�#Xs���aY"Z_i�%iw�y��}�r��~��v���}cCS�ZHR`�h����B����7>6��Z�ƅ-%�H��Â��q_�i!�r�u,�V엥qss�ث���s/�qm՜G��(1.|�A�SK��?�)�K�����>�q�1o�'�`&A���	�Kp��E��d&6��M�ӣ��p��J�k*�R�r���(�K�J��	Z.S+�
c�����`��ɩf���01lXB��(�X�Ɂ��B<G��i��5�sӟ6��f=I����~���߫�薙3�����S��i�p�s�?M��dړ�����N������HZ"b����F�n��`�P�i`^!� �i9^�rKؓρMGv��n�.q6��5��l/á"���3��?�&x�*v�ޭ�����[����������⑪8/�Aq,$���&ħ9WIu��Yo+���?*��Ҫ1���%ޝ_3�_��/(�J�s���/7��I��.s��xl}��T��j)y�d^\u�M�G6i��%}%R�M�z��uˎ
(ix�+��{ӕdƻj8cT�U�BXp�0M��y�dC�3��N$��W��q�!j']C����?T�������t��� �-�yS��f~�1�?L��Cl�j�
�XZ��Y)"lߐ���+3\[�|�]5�K�L鱿P��9/����d��tӾ�Ǉk��;��>�������+O�H�^'(�4�9�ОqJV���t�,��)��_�X�i�����zU$�L�<�i: `e��-���Qb$C�ʛ���V~.Lt�4�����&�cU��K���<����E쪶�~�4�4�:� ����u���}��;k��Q6�p[�g�=�|�Є`��lS�Ot;v���I��J�nT=NŪ��o��y�(-6_��߼V��c�g��M�o��`���������}�F7��/$q�إ3�U
��O�]�2$@_yn�/�4���W
��bґ�],<��vK���KM�0uv�'�M�r���l�m�Rqdh�t��֕�X�h�?}��<�+NC�@�=,��R�<\@��"��&�����E�-��ZzUަ�Ȥ��8��
�O�b���ܝ/L^�֢���Ev��>eZdݍ�����Vi�t��!��M�,է�YXCr� ?��Q0�jg�TR�SW��J؎/�M����o�� E�ŝ�@Uh��u��f�}�]U�!u?��Z9~F��X�t���S��wK�ͫ��n<��wiV����m^�X!���[���yU���|L���։�0K������-W��dP�j�v�Z�&bR{�h�V�x��<��|�j"���̋�L��7��#L	��E��qS�ctb�Vr��+�N�d�<IX�[��EDx"mA$P�t�-wyA~�k(���A4s������h�7F;Y�Jp7 ��1�� 2���.S�c�Pz�i���u�U�zt#��z��ɭ{[3

�6r�����L%���P[[�u$��<��K>�od2ELQ=�P�j�������ß�Y��'cS�A�8C���S ������J)��W��F�7`�+K�{q}���ˣ d"���,���9/`B���;綆�1���~�Q���`ьO*�tu'E^�����J/m�ү���vx<D�>�|bs�2'����J
� ��(�,������O�2��>��/�Zz��&�����o��HVs<�����z9N��/uZ��$�v[."��D�)�}/���k�c�u��XđJC���;��C����G\$A\brx�+N��7�-��2�����V�ma�Z d�E�s� u���r�Ü���0�����{P�!HQ�"����΄�^��ا>H3dB�lhB]�DɊ��=	s�)N��uڌ�.��!)S���I�����`#iy�,���u���@o��+۷*Q3��B�Oo���C�%5]P�RB�ڼʇ�iSD`����'D��UÄU���B�6�KH2�M��)Vg�9��`�)���}Ir�X��L7| ��`,���j'����*��i%��������-��4���+�˼I�J����y���������V��0���6�Jn�r��3�UZ^�4`��cƾs�����.I��ڃH�x;,;�J�ӡ'���g�`ֹt���-��$���GcyN��ヹ�qm���$(�!��N����I�y�N,BU4l� �0Mݠ:tFO.�r�ԕ��
�j}�|��M�S�v�z��>�����*��DH��s6��D{v��$g�_�1��o[r�g�X�N&TZ�e�Px�0���ӣ����?��|ׄ�`��!m!���Lϥ1)�ڔ"@��io�͌���TKF*���FG����F
0�Ϻ��%qӈv��ڄv��O�߭N�2_$DM���W�q5��6{H~�<�相�@R��U��G�*���u7����DԨ��K��^A��"�
F�˕�uݠ���W݂�8��m�x�V�ߡ<�J.�o{�P;.�U�Q�Q��e��Sd�妄��N��"7m�� fDy��"���$~���F�5��׮����cO��0k�����7-<b&
���&�Y�1O��	�V��=We���=���R�|�d��U�˖���<�kޘ�=N�)�ψ����=�n,;���b�ج�b��]`�!Է�TZE|��{T�m�kg�-
������{��M����aڎ��B��=�F�_k6ߐ�:��j�V$gt�$�m� Yi�]da[���N��;��
�<K8�n3^7it��9!��6A��E3�-�u^	�E�B�8]:m/!�eH;�~%��=T�w:'�y<��3�M�j� �֗	��{���H��(Ԅ�ʏH�#\\c��X/�<򭖲��/����W�;F��L; ��~hU^�#�8��3���^�{�g���?#�"(�]�F�]U~�H����E�E��!���񏤖E�>) F��d���:S�z�C|g!�ٛOj�W�%{F�n�����Y�x#X|c�½��ؐ�k	�qT�v,!�������MNoU��<�M[m�xL���-:'O]xY��UX&�-j��z�#�
�D���0��Z������	ϱW� �-�Ե�o���$�׭�\H[tA�����t�Yr�
F�/�Ek&�Z(s�2��v�������!�������� �W�㰚D*V�9�7��ztnv����X @���c�U�Nzy0���Mn�\�Li��
��Ni�%%�=��,O���������Z�\6��Ǔ`	/�x��oe��Y��Z����j�YB���]�ơ��g}9�n����҄�#먇��$�6��ڄ�30����QK�v(�ڶ��� )M`�v�jV�i�@ضW��P���#�O��'�KXh�؋���z3;��(����m�#�a�'G���g����[�n��h3x�Y4��3��}إu��;�x�*��|�y�kQ��.o��IT��B[�>����e[s�?S�M8��
9i!�]�][�%���� �d��<g޿��i��|����aj�l�6���#���(�?�r�g���Uh���"EE�1w���Ƹ����V�1�99��"N��I���)��3%
Q��Q���](L�]��(M,9W[y|� cz̉�b�ԅ���;)�u,� �U*�m��E��#  �e��	��A�>c����b1-a���p���R��o	���s"e����%?D���v��mI�/�[�ܑ�^�Ս5Ɉr-w[�`Nzt�F̺��3s��=��������)�ԭ���D��5IqahUq\�b�TA�;��p:���YL�ε�PU��� l-u!�3��ե�X;C���p��� �x�e|!�U�
�Ҿ&6�Vu��8@���<�6����l�:�=�&Nt��W�}�M̕ı�	
p�<*U~!�ٯ���m��Je�6l!ƫz��D�m���iU?�)�%@WHֆ�F�Ҥ0M�t��b��C3�K�Y���}�4�@����_X��r��1"	���>LlvA�F)�ߖ��IX�:�o�� #K�MaQH�GҬp����w0�U����{�'t�����'N0����},h�7�a8C���C�k?#�媸�tCm�f�A5�(�2�1)lY
��=v81bN���N�O=uԖ���5Έ��hF���-w|{ֈX�G2H�?�������1uy`��n
-��n��؆7��u"��t�g�&]D�����D��/��1FB�I$��*@F��Q:6"��V�c�����^��^��0�P�K�3VI��^Y��D57��_����Oy(�*e��恲�-K�%A=N�ղ������0k�n<y�҈(�;��/e��3Tz� ���E�|OQ8�`�Qg}���E{���.���U�����1�������)�s���p���-{Ħ?Y0F,��s�ҪPU�|�A1��t/�h80s��K	l?�}d���'�2���X�*B��R�.[�4Gy�ϭE����]�����3������(���������i[�ߦ>�ʻMI�=x��OW�����$\�8���q*'���������ĥ</7�PC @)���
_�S���Hڕw��w�n
�.�F���ă�+����a	��!�c��ZI��?���Xk��V�~��p�d�<k餀�$���<�<�J�7��*��¤�yD :	�b���dz9��b$4��x�+�X�A`� �۸�V c��}E��c��و�5�q\}#1xq�I���ڙk�9���އ(�;��1�#��P�����s�t��<t�-��˕��ƨg��ph�m�Y���8М㳦�����3�)�y�@��T�m�;�آlBFJX��*d�}���[��c*�dv$O�P�`�<h+g������ĐR�'��b��!��:_�L�7� �d�S58 ,��?�����ԩ���^ʁ�"h��]��̬�-~��P��O�B�	L`��~��[Q���z��m!�k�^���������"��r�E8�I�T����yL����YtT��Ņ��ܣ�R'�A%u�"��F��V�
�1�H��1����_��-)*:�|���4�Zo�8,�YR%|3���G�ί�=Z21����NM��/#ǻ.�Z@�ua�_�0��m�l��a�!I9�gI���n��6�
��^����1!���!m�A"t׾S��B�=ep�5_1���*e�b@��)u��d^^�TyŮ(m�4�+��4����U�b�c�$9?��pյL����H"բ�6Dȭ-?لl�=V�#��b�ŀ��p-A�� �F�Y��iF�v�)��F�h�̓���1Agf���^�9�Q^OW�q��y���;�q�O#4�.	�&l������D�THl[����0��o��|D]����Y=n�6���N�nji��g����{Sx�>}�g�0���P���-,ɪ����*���B�A�$1A�'��\��v�(9��#B&����e�?/��Fz����O�;StXЅ]С�j�����Dj4O^���/`8��b	���<X99rgބ6�iy��}��`:�����{5��v�3{kW�M�I*r��ƬhÜ)��H�����"\wv?��*�m���D4�����b��х�-�Q�
e�8�Y+M�bV�^;g Ƚ!�N�Sʈ�)��~������FO���dK�5$��z,NC4��.���@�C.˽wDS$���~~� �P� ^ŝ��2d��2�`����k��x�<�wI���Psɢl����*�x��tر��i�<ܼ4�aC�I���a�&5<��P�h'B�YrE4BS���DkS;�����3k2�Ub��'��jC�*K6>é�����"EPr�6��kƒ���	
z��o�]ճ&�I��u��9��$���<���72�*,w�k	W蕹�a���
�X̽���~����s�_�ju�ЀK@E�U���#�X���5��@�BI;�?S��k6^��fi�������<��q!�jPQP���Hz~��=�R]�[�m��C<������|�hr��[>�I�(��[[A�!&$�1ir|��S�E�f��g3�?eǻ��X b�;���V�'�D��bt�1
��M�y$�)�~�K���DON��*�̵ɍ�s�eN�;}P�~����
��(���q��^zcr����B��K*�O���㡱ߩ�ܺ��w)�R�������Ϧ� ��v��:���"�<E?�_��x�bW�s�f�~�7#r��/�WB��,�q�g�����k��ؿkQd�=d�
l	�%�9rǩr�}�M�	�r�?#|����d^t�d+"x�pQb3^�o�\کl�ݛ�K�pa�8�1:�����l����Jc
B����=�D^��x�l�U�v�YC Z���ױ)2;�c��/�6�D!��2L�����z_T )�
�ϫt�IAO��R��9ʴ��-�Ǟ�!?�>�<@���z"�8�#����8��q�A��w���0�@�����b�<&�2^W�+rr��NK�/W�D�9�`f�j\{���t�פe��n��Ga�bP{���(�A�2N@�퀔�~��Ȭ0�ğ�y��&)�"�XT^�xS��d˖��T~�8)F�����V�x:}��(�T�Z�o|� ;Gѭ��o,^�5.Ҧ[+8/M`��)���'gڭi�Z������K�#��9���?�W5��BT�6��ӌA-S�j˩;�R����G�[v������>�QQR�i.K��73��T&��u�1\~g�T�!�%*0�l�� ��z�w�����n'����E@
*#ndCro^��n@b�j�l��l�J�R�t3�� ��4f)����7_���]����"��%R�t�0��e�R�	�ĵ�������z0���������óL"�:�t������	"^��J���_~J?\[��op��_���V=�=0���-���7I.�k�7n�f�?���s-{�)g����k���Y�L�giy���Ao��7���]��o{��7�`�ͭ��p�~'�s�.�V�׵��HpQ����eW7nFɫ_A��i��U]����]���K��6cDGI� ���>�u���@����=����;�fd0���  �v_���f����g��X��=� D�G1�� Y "��71["xB�$��H����#�������S��t���J��5��r����hA���v����F4 Ŀ��*�<a/���I�)��=?���%-*�5
ɖm�쟰��b_��5]�v� ��b�!T��-+�V��[��
[�@���2o�����(�������fFl�y�W�2�ז�>��ʐ ����K��r���3����*�V�S�54F3�b�d�\�h�G����x��]�9de]�ag�W�%�J������&S�j�)�A+dI/|��e�c' ���`��B�p�5�5_X��_�O2`�O�ɣ�k.n���k�i}�IEE9+��rvjn�i�^�>�5��VK���DK�����G�6w� �P K�o_��ܫ�:��ZL��Wo�+�^�BAn�~hnp�zk��qf���!XC���V�Gej4�]7�_����kx��hȒ+�J�]h�D�l�f7���I���t��p7|�y�����I���dϊ�~�Y�ܨQt'�����B��jZ�Q�M��S�."9�t>#�����.�31�ۘx��ߐct܀|�U�G'{�\��_�	���ɂ�6��]���j����HN��vF�T\���(���>�n�K5	3�kl�g��_
$�W-��Ɋ�O����^�,ꏽ�#I@2�wo�!N(��M���ެs�h���m.��\Q����x�7�Xan*:�bo���B"˭떣���
�x9�UR�\J<���׾@缠3���Q�ǜ�̛W������}���"�x_��b���k�ߣ��|���
�M_�De$Li�	��#�^\[����8��VsJ�����~!?m��6sQ���b�C`��'ٖ���yTM��۳���#�;���i���Z!�P do[�����7�`(�3u;tef���!  ��?��~��}�l���,0�D��c�wlA�ls>%z	�J����k$+q��'���]��T�Pm�j�Ϟ����`�u�7Y���G�^Jk�Z��˰��ʢhF}�t`ړzmqS*WQa)�*`X�ڀZ�"��V�Û"I�,�5ȥް��`q��� d���5ȭ���A�}��g�Em@�p���nd��M@�f��t�Q�6��u^���Gن_�(*B?�"�藮��1�k"_q$?�9��G������r���2�&��������={'�.��m��/a����/�&
78z�~?K�L{�V�w��ƔRp��3zGuz"KN�(G��a�'�9/S�v���x�5����<�P��}��L���:�pڎ�E8	��0xEzkHTL���A���G��_=� U��	�h��X�
���ň���J�ܵ�?K?��O#r��v����b��[\k��ō˹��.q_')HՕ;n|�K�'��t���Ȩ��cm�p]�>��3�p� il=�q8�d���j�e������L$֛�\��(�]�#��������fc�V�¯(�����r�8�M�G�Vu��ע3����}�i�e�+��d�����a#��E�r/ӤFO����'�M����/%4��?7:�;) d,����0�q*��B�?4K��-������j��*H���4�M�������y��H�s�KP�u9�XjV"
i���I��@YX�z�
=�c$��
3�-3�O����"���qSI1؎����б����?�V�v�,H����к}�	�c���8&��2N��v������>o�<�U�e>r�a*������(t`.4[���Z���I%>��6�(M+k]-���8�����RD�}�1��Z#�Z��KH�K�������㘗.v��rw��"���jJ��*�X5���ؤ�{�k�������]�ǝZ��e��}���'_k �H�Gm-��g:-�g׀h��Z�$(�5:/�������Q�@���j��<q����Xz$X��ݬ���.Ԩ��S�H��;|��	#9�L@�Y��}ׅ:�2��J���{B�_V S�:2&K�IMZEe�2��/W�g��\��.M~�q�R$ ���ӎuJ�on�9�e�?]P��CNF��Z�r����7�@��I�V��������v֡�+"r>�r�k����~���cl��X�e-(��yW2]ц�.���j��(x���%����y�3�XP���ɱ1������NHWiV�c�i׸�.�&�=wv�ZkB��7,xH��L�!T=�����.�`AV���DKܥ�zQ(�S�o�1;����J�?' ��Ղ���ޭ�f���KT?Ϣ���3 �x
������d�&�쾐F����*�>]� r����z�〽.~v�� L��Р�a�����j<pk����j��^���t"�?����,�T�ϥ&&��W�ʪ\׫ɛ�<�D[�r�^�%ݑ'Yk�;��T)L�����d�,V���O�a�Va����P��|��Y
ђ��{�m��:/�99�;�����Z�|*6�p��y�Y�qƘ�5���$�}B�0E9�S�6���x��r�:I�-�[��dl�3¨{ױ��v]t%|f#k�3���k>��_�UU�G�$/o/� ��ZR;[K����0�b[�+x�'�~�_W��4���t|�D ��^W��@'�hi�����p�0eO���G��?$���"3��u�,�	���<�ҚI�jy �Lz��כ�K%Cޛ���Y�/6�����g�%�����Ǫ��M,^2��%�ёI�{�e+_zD_|a�|@Z(y<��ߔg��-	ul�m������'�o\%�z��C��X�ٳ���W�|�u�6�=G�����q7��t;��f��WXӅ=NU��@fәqd `�kG�����r������4��ㅻұy��E�~�YwC�Ng��N}�)�N>��ǐ�wV�M��F (�j��a˵��A��H.�/�ߧ�1Bc�J��� K'A�U�]H�^>T�b�i��Y�Jb���H[:�G�=}a�A՞���ٳ�GO�ab����&O���@�M���Ù��
{a~�@�f~Y��?	�U���e��8����M��< S����:in4p�bB]�=����Τ�0�z����;���/��C�敄@�0Gk�I��?���?n��3v�P�Sw�8s�� 5��Jޑߝуi3e�@��G�(B+^������pO���R)0���?d���D0х�02)�Q5: F�@����Ce�;J�Q�� �z��ȇ�=��f; ކ�s��V����lw�qt'g�LıB�)3 J��l�(��#��G�v�G�_�V?rS�h�����5��J�8;�=�.T�m<Y�ܫ	,{xט��TK��+�W<�_^��/C�0K�7�[k�`%�
Ы��$�	2�`��U �?�d��I��k��U�H�\M��bt>b5QsR��Yi{� ZN��J�����&p�0�wu�MB �B(�p��T(�s�1�b����e�&���R�%���:)�{X3�t
$�l!�,\'~�E��0�����#]~�>�(��Iq���-AUg��$Q�ȹ�눇��Nǔ׭��x#״5q��<U��v���$��U�p�l�V�y�Wߖ��'ϻ�]Ѷ
����2O��F��Jr�h�E;�}�׌ �R�&'QjY+�D09At���E�r$ƞ�+�h�Md����W%:���F�^��P�Zn"��~L0�-�/^�����n�v�Cʆ��W�hh	�Ps{\�^a9���f�Z��l�!�*v*����b���;l�0�H��G��g ���r�v
R�X[�A�t,t�+Ɗ��?D"�,�2`��n<�l�6_�������O�h�����\64���;͗-xa�?��wl��&���~��{��!5��4��{�Zޑ~�CB��Z�
H���L�=��W�7�j�]�!�5GTΓ���&s)��I��=U$���k�����_K#�R��$���b&�L����v�e#����͖C�@��,�-�B�/�M��C�)@<f��%2{�&�Ӭ����1���� �U��e���ed�Kۏ8����Ǯ����}����ОkI�OI��T�F���%+DN(��)�,��{�xA�b)ݨ5gO��+mIS큾M��Y�~�˄̳oiȗ�:{�u�	"2o�""$��ۧ�A�O^ҌlJ�5�_>KW�-���ju �����{��:�Γ��T}�a'�����JɦL��/�5H�����Gj8y�f����>ˢ7g)���X{Q�5.���q��m`.���e� ��KFg����6��@6����`TX�FU�(z)�s@�����
���D1&�e8���&]��{���O-�oE��X[r�Q��>��!؇�ѻ����b��(9���ds O�FM���U�}�ǩ���t�q�2�5�TW�0��;�ɬ>����Q��
m�k��ۀ0������C+4f`nR�[^�xj6K�]l �l�^u��4+E��B�E>���>���n$U :�=bVǃU���-=�߸��G+u^��˚�OE��"3*��f����n��#=�*�|���|�w¼ ��I�v�l��k4ad��d�fр�y�~Q
9[j�������H�����|�V1O�FAfM�ф��}�&�'�(��?Oaސ�i�I�H�3�g+��Z]��L�o��ς'7i��>;kV1�*�}-ɷ�UƔis̺���o�(q&r�o�"�X�cfj�i\M��t�VH��&wD�O��J^l������>៯e���d�p���*��[r�86|�8/G7��v[9cl�OQU�Rr������m���l�MV����	����B����c�����P�=�p�q��s�:6��J�<%{؃7}+Z� Ӫ*�!�ԕ���L��hE#Q�>�,?o\尣haB],l���Q��w�ܭ'���YQڄ��z�X��p.Ó����b�P��ݓ����ʕ�`�Y,��
�>���C� �T&1$
��A�M3V�O���I�ٖ�_	:"�Ap�H�9���y��m����8�n�a�k	��Qe�������L�Ҟ�(�ɸkخ�1�2
���B�^P���$��	�!�ϔ:�l�G���M;i������Mb�_�<(���=�6tL5(�k�|4=���7��<�7��Id�����=-���v�U p�G��bO�m(��<%��Xl]��ag���X*e��j�aR��iީ1FG�f`J�̸�u�b�?�����d�lH}���hT�%<�.0x�Ƌ�B�H5_�y=%���U�JLR�uHr��XZ��G^�j�g�u0�f��43�z�h�w:A���%����,�;�sFFӁ1��̃&�!d�@�p�hZ��gU�9f���4��Ѝ�<��s?�I�Y�t�@�g�̩I��;�E�e�跌�*Ïx��^�lFF���6GX���L�Iqe�_�0l��ሻ��©�[xöו���J�Q&����pJ{uX�=��4��: 5�ȳB$D]��XXL_P�DN�q?w�d*����Sq(�z6�ڟ E�~x�s+2>r���Ex��0��3�.|Ј��i`��a͔�eM ������gi���@��*4���$��b�["z���o\����y!éXu*yg��HI��xj�w�2�p��첡ǩpa�?-=�7TnXU��^}ЃQ˛���'+&J�|�~��4�nw�A� YsUT��E~���ϔ�N�����}s?^��2鑉��%�U>�)t���YQ�X���}��{l	+VQ�6uoM	��	l��ʙ��%D_5w��X�N����%;T�N��W�LR߻���7
�}�Lv�p�}�h�?���?�G%�%�E	��K�U��������|4�z]��)��Y�+���������x�T��B��9�y�qu�dOH���J-�zo⑵�PL�E��(yon� �p��S��-�����{pV's�x�S���/K�+���v�.���d0�����y<k�u�����4�z�f�
���:I�D	�H��G��{j0"�����$����j����r��^@6V�Z�[��F>�c@-�Y���\o1� � �Yq���g����0�^��Ynn��)~�hQrЖhm�u�b�z��h�cB�ܐ��R.���cK/��u�x��AҜ֒�Z��ΔƈDD��G�V1s�F��F�v(Оdy��P������,�L���c�=�J�x;iF ~�.�u�A�c�(Q ,щ�lWax��ZW�~������wĩ!"�@;�6E{�އM��}pb�AG�5��0�[$m�{T��T�W���� ^��r��FX-�jP��m\0��>J���x���D|�e+k�7�{Z���+c7�����NUE$>,���#�M��ɦ�i�9��K���3fW	�uҩ[#;�N��,�Z[$�@KEn;~(�܂�H7bRf�\(/L7�z)`��������K��q��D`�O%°m�P���[|��doA]?��ٌNν|	�Z�}S�V�F��!�ij
���o�h#�ݭ3*�~a􁧰�e!Z�th^?-�O���>��[�s�?h
��M����"B��_�_,���6���9�|�{4jR���\�?�I���`�B�pb������L�B�<����\|P`%Ռ���3Tr�q
��JN���]ޞ�W�����W��v�%�+}��j+U��t��c(9�&-�W��{�#A�������̃n��'�$��`�9xs߂Й����G�Y�9�G"k*�\;.7�o#g`����ظ!��DP�;�ߠ3��Z��vaI��(u��6��ΔS>�, ��VTZ����Vt �"�ا_�U#_�#ga!>���+��&�%��Z���#�^��t�N�W=�n��<޲Um|;�y����O)A);W���<��@�e�F�!�-��GR2*������:�|�\]ߖ���V�e2���pl}�6^ �U�~�{�v��sj�ڵ��N���Q$���BAe[+�ɵ�c&SF}}�pi�R�'���C�S<�.NfA9�F�w2c�oM)ZګLØ#��ԃ�U4��˾&aW,c�֖�mVr)->ɭ�@�pR�<��e\�%w�ut�8�wd��P����j�o��G�ƭ�*�[�-�<�Ҵd ��!*{�����KO����+����{���T��P���������=��ٚf�x/RV������n7믻�QD>���X|�fgi7DP��� j��h�J�b����^������!��`��Z�1�$c���� /C?X;Nj!n��M�.���*�?�$b+,n��k��A/��y���?��G7���d�m�����"LH�32L2E�q�t`;%�M�/*H�i���~g�j�-��ֶ���p�[2b��5~�F
� g�od���R"Z�i�tg�ƻpukPA/&���\���喽&BEẂ]zl�}ҩv���ډH�J�'���DaF��ˣ00�QJ?J���T�D%A���=���Ъ
5�N?�pm�-{̷�;*V�a��E�&�ꍮ�}�_2�4F@�Mָ�����
����U 䫚��FS���R���r���@�6��zGZ��o�ZH��,sI?��Q��8$�u�˗� ���7��3���ԝp�W�e�I�2~Y|���b�=�cK����V�bp�d��I�ܛul&�B�άEM��*�ï�亚��gbQao�b4�Lۑ6��;���`�h:��t�=�-�r�!�ĭ*���=/-��[+�e �m�M�f��B�_�TI%-g*�����6���O�����s��Sv�]$�	+|ۍ\�,J�1��`QSY��t��bKQx/����r���T�t�PG�TV^a�@�����n��C}g����oBZ׍t"�_[����	��!�|؞�=�[Q��C�e�dOzn��Ζ~��,�"^�Z)X.}�ʲ�28��)VaE�.pGʭg�32���V;��sui�(���WT�(�E�ij�wU۞T`z���.�� kʐqs��%MNՑ�'��� �99Wj��V��c��{�����q��t6F$��A�z�5���M��.&�I���>ؖ�q⚁�&_�基��A-�rF�f�
y�j3�b�G�E�n���>�G\�����KN��VF"�5��d|*�ֿ#r���l���� ��0��mGj�ag�(�o�1U���371��?��%��z�U���B��00��J9��L��bk��\�4�1Jd1*W�P���dk��ۜ�M�Y6�l�L��<t��m�W�"��Z�p��(T�uG�BuҀx���VD�u���t��D���.���_��O�6k3c�db�N�����
{`츠�'n[QV�G�s�}����Vp�����LK�Y���ٕ[#8��	�^�>��9}�C�%����(�ߐ��5Q	o߻@G�i)O���p�Ǧ�d��A��Ҫ���K�T���;�8燻����G���)ra	6o�Z%_���J�1����M=im�#��b�93"E�[�ܚ�*Z�,r8}��:�`��F�w5���s܀]��w��x���ka1�`����ɻ.�,��-�2@�x�5�%���=��^���[�y���  ��=��/���3,|宻You�*�������]��6�&�$�/�)������%&O����"%35e�yV��\[I�y��4��31��1\�I�Wc���33?���q)�� 񢔇����o��<��e��u���	�I�����s2	�:x��%������7�?�)g|f��w�'�ZmCS���{ri��@?���>>�ݎ��F2��,��x���p�l(W���ef}Rq�
�2�W�ޏ��(Q�e�aT���*S��馵�=(\���=�f��G��&%�~Bݜ ֗v��;��9	��������>K�>32�!�8v87� �����������ͬd��Zy��:�m�3�qv`�j7u�h�J��Z�z�`���(���z~�L&)����w�EJ)���!q=]ޡ.�x(͹Đ�-s�����\���&x���<�%u`w�-��F����1D��R*�	P-:��7x���9X�
��t�!��Hˋ�Õ]�t�dO u@Y\�Bz�7���c xQ�������,e�i&�)��%)ɵ��\Y��zHv�!4nAӴj+;{��=�Z�<a'�dw����q���C�����
Y^2�ϝ~�\����ڀ�9�j�ë9�eu:�6E�ۣ�$\��:�S�z.����W��a\��4��y5���CU�����Bw��o¥U1���2'Khy��a�,?R�qlӓO�(��>AF�S�g�N�
�R
����dB�' ��,YϤ(3GW�� �p���2?� ���vk��{Vp��B�� ����ԭHÒ,�L����@����=�e���`]�	6�8|`�P����(�0���,9=F��"BAH�S�61���q���P)��
ee�㿶B,���A|�����
;~��F�um��^�L<+�f�D��0��=�9Rr���H���<����Cg��h ��!i�Rߴ�/A�G��w��y5��~bi]�QXV�nۓ[�d�*��C��r�N��su����I�|��cΠJtV�A�����Y"����q8�*�l��Y���H��f���=�؎@����$z��������λ5�j�`|�g�OG�Җ���k�
��d��sdj*$���o<��+���S�C����
l��pyy��6���e���tݑ[���
�vr����֢8����
]v�)8��q���`�h�OL�5�<.P`�d��lfM��U���9����y$lDF��)�yDp��(�3KU���/���R�"�!KvG�^��m
aưԆ�\��c���p�Z}F8.�	3J��E����	wi�B)׈CWL�b�oQ�G�/�Fp~���-)����q��F��P��R^	�4P����Y� � ��%�i���/7]Nf7y�v���b|�gR.I�iy&g���g2(��S�>m4��h�+���h3	���	As��g>dL0|���,N �v P��k�s��d4�5#��T�}���r���*�L
�����Jث8*I8t��@sNK�PE	�Q��٣l=�-
4ܿ�{���qjUD0��p83Kc���R#���k��&��%�%�+4��L'��6���90L8�ٸu��,2���Je�g�"�^�����������Qi��K���7'o#g���Ui���t��?i���� � 51�9�1���n���@���?Q�Iv�^ٛ{�"SK�s��p/\���@dq�6�.��F2	G��Nm��u7�|�U$��]���Y[>j��7'���w�Ɣ9VˉB�c_���p�&#�Fk��A�px� }�tP�c������	�=���E���?����C@��|y2��DIIƽUN5�C����]ݺ��������ŝ�,�
T�8��Z#���0�EuEX��q��b����#���un��N:�1��N]�~�a�ɇ��5��U�fz�9$R]Hv�8��^�g���9黇
����V�}�!�A���q�`J�O�� ����,`��@���E;�Z�?⥒��Lԍ)���G5�%�k�T�e=�?IU6�:�+�J�#�����c:}��o����3�X1��:��y|��du��)#�\f<�To>Y�Eu`F�Va9Y�k�~N|z��$�$*�`��sp�"4I	��?��J�?�OҦ�vv��U���!����Wn����-��������s|@h���)�4{pfAڑ��w0��rJ�,KKZ��H�o�Z�&���@Q�����B��U�.vu"�춖�M�&����O������C�J��e������{�Ƶ��n�j�aw��6^^�%+'?ɢ�����Ul��g��eF���2�	Vw��G�0�n�[+�8r�篸�g����.�'�3q^��IQ�����(�A�4ZF��IK}�vE�#Èڴ�z�f`��+�dHS�����VXK�ӯ�Uwx;"^�'&���h�v�1J��Lŷ���#�̂+'v���rX,�-��%.l�ܯ�����ǲ�Q�`�9~]������o���!�>A�ީ镝+/3�)��&�$Z� ���	�~�/�e0�Io�����z��*��ۨC��@@�v���� �Pˌ�%v��5o�J�[�_J��߭MQ]�ڍA��n}h�p�
��W�7�ʝ���ߕ���b�qC{���� 6q$�<q��ݏ�e)�훕R~�c�������4oD�S�}t���%s��G1E
�{��Ј���s��G�Vrk�{ʶ�}OM�@~�2�q�t�g�)��pt��:�,�����9�	q� J��B��Jf��y�j�Hu���s
Q��YÁ�l&� ��E~�z�y��Ti�~�����|o�a�p��,�*��u՛H[{�E��E&v��"���$7�w"����f�=^.%x�
���*��s����4�@�F"zU�`^�!������t�S�]P��W�/0��8��P���\��҆<���(���Y�,����F4,`5�����j��|F�p*�9%�q� 1j���2�e�R��RXC�%�yX8`��](�$��(N��D}���*5��HDxX����cW�dy� �{�UBvsJ����
�>7lM*P��mܪA�u�5Lh��{⦽p�~�9c��O��"��D������6;�P8R*�X~�::��Y �y)����'K&ڴ����1��՜�����NC0u4�`wĺ� ߧu������S���1���?⌠4\�P�a���''��^}�5 z^&Ao�z�-�,WI�6$�q����:�!�ː��G�T��M�ң1�>��[E��B�:3�r݀<b��M�ղ�S�o��3w\"Y%�T��|����/�� 	���L�"��b�s�o����:���ֳ��N��s�6�k@`t��J�{E���3�X��$��o�"b�[�c��,�ʵt
��//�vǎ��~��cqh��pЯ#���O�ə���԰gBNv��Y���Tlb��:(�l4�TEƎ�� /��}�C��4!��>Tu�3;Q�b��Q�p�1���n=U�"��~Pa%k����%��,����~K7����"-H~bf�Ī
��6��q'��f�oΤP��^��5 �U��<v�ƶ�w>ۙ8����GՇe[�~��vE���Ac+%G����h�|R�&�T.��Ȍ=��%������7C�h]b�Khh��i�!v��Fw|��
)/Y0��Ξf��/I��0��TGv�l� 5�1��`�W��a��.��.���J������������Sr�F�Rǩ,����5��J���pY �QMd��͝�N�	�@�I�q�V��NK=݁�E�aGy��$v[�����D��}���J��Uf��ϴ���k[��s���(�`�����\kW�L�j��6P\;ς���Si��t�ŲpS<�x��ֲtˀW�-��ȿ��4�}V�l"��.��q��О˾�\mڷ��t�^�����9|��+�E
aZ���͟���$T"�s3h�;f�.���mb͍��G٧�qw�S��4�X�t�~�ę`�$���ƅ��CpJM����E�r���:�+�_[�&xR�:6�j�Z�ZaD��Ĉ��}@9l�L}%�F��K����"�ܕY����{!Z��}w6�Ԥ��hd�[� @�\�<n���c�pC�
���� a�e%sk �q��7ő��o����	��Ƃ˥)�v��	�#"Q��3���C�{����O:��'W��@�}�U�US�?���̕�4Z�h%���f��ٰ��X�>L�@��q��]��K�P~��ui^���Aƽbe�gUm��@��)�9��K��v�*�4�|7�ћ�cշy�M^EX��}����ݞD@����4�7��#m;�&�^�	(2�y���zQ�|�^��>���$�CN����aZ@?��Z���C���5��lQ���J�C��&Bf�c(�����γe~x�*�f����_{Ԝ"5�T���]��r��Oh^*Tѽh����VA�y�嬫�sӗ�����!�� qy.���~�7h\H�J�L��?�����qab�������+�����-�s,8�LcU+m���"VI��4#� �,�;u�dy�����fI����}Ie� �H���ޓ����U��� @k����헸���>ː~���O���6	n���:w���q/V˺ݮ+�Q�q/u�X�(�F�8HWk��\�FW�O	 9Tul7�T.%bP���Ѯ�Y9���x��Ŷ)��_�[���w��.
wi�[�bB-R{b,1��I�����D�`Z��A����SQ޾�M Z��{{�Ir�V� E��VZ�(ڠ�c�<$�;%W"e���&Ds���6-~�3���h$�zY� n�6,|�\�٪�`b�ce6s���[<&rE�d��r§�C�_�^��#����fSWU�ɀ���@L\ۆ�J��b��w���ve]���KI^6�� wЇ���c_Aﭺ����?��&��l5�{�p-[�ǔs��?9�z4�݁-TFGJ�� �H�ͦ��U:e`w�`9�9>� R7�K����K�
��=�^���<�w�cI,p�<�,9,��V���~�닔Us�3p=lR�j,}ve�іp��mFR�Q��~�":oi�����8 �a�%t�0wN��̊
��%<Wy,HLv��<�5��񿀵��ԗ���l����-�k���Ɖm9����W������ �s�����>F�˻P%\p>UI	��XKD�	YQ���?���[���c���|�\o�B����M�Q�#�B	?�����(佱���@����_�b��܎�|9 X��{J
i�d�\�=&����[)ßi�B��?X������p�A��,�D�F�c`{�����R,�@�>jC�9O��޸va��;�{A�!�n�$��C�b,��#l��������i'�X��K¬���m�Mա���%kQ�鴃&u|o�m4(C�ĭi3\:����-}�b&k��6�/d2�Pa��eB��@�����.k_��R�3G��N�Z`����[�%҂�Q�	~�뚵E�@w����E�ԫ����#�0��6bCL3�����g
�kLK �<��vōff�s�hg2`�$�RP%p��2@Q�c��9B�WFaL�p�^�|��0�4�5�A!�|�45�y�ē��0��8_�neW!�W>z�ءe�C�)7�
�MYjvǓ�a3QJ��V/���X-*Z9i�*����$z�j���J��qB�W���t���ES�*Џ��g���[�õz߀-OD�o�!' Hc��c\s�Az����u��
�@�����_��v�~�I��1֚�b���8��cU|���.~4/��6&���W��>�i������+C�s�E�m���n?�͝����œ��S<5�D��M2{y�Y%��j��`ϥ@���j֣���x� �/�^��O1��$�ߌ ������txZ�7A�h�ɯ�
��I�ָ�>V��nE� T
���X�=�R`+u��[����R� ���GK��-�2���ޭ
�aū��n�4� �Յ���0p�v�_��4�s��~m�T��I��/��jc7޳�̰y�	�CV ���j
<C�V��J��y��%����td������M� ��������۠z���쭮|@�z�YK�����X!A߳�L@ÏV����J��j�\Ď.0 .���^��@��S��l䢡��_��.����>	��ln|�Θ��#38�I'*N�S��c	Ά+��g'���6�:ggp^@6�|����1EW$"�"�G���N��'�y������<��Z���ND~���u�J�$e�j���.đ;��Ų�z/��h��?�V&QM�0�������A�œ
��ŋ(%V	9CTO�2��󓵿����Ͱ�$s���#�˝
Ct-śx�N�
�8of�����إ�е�%�="�ޗPu��X�/{�z�\������AmP���g����1L�^���7�� ��r�e�������o$s3���i�}�r^��i<���!�K�(�U�S^�����e�vZ��W�͠~\�whfbBC�+�Fb�p}J.�8��$kl���1mR���,=(}���'oJ�5����0~������3O$A���4����jn�M����R) j��i�>���X>^Yx�y�I��Pܯj�M��N�eT�*�	�^(�Ft��8�X&W
Ͼ�i�A���J���q�%It�e��.���v	~e%*�c�녬+{�j�w�ATc�9^���w��[U(촃03�~�cިw s�@�=��j��L��Ǥ�WB�et'���G;�M[W��u	6c�����%��IN���:�z�>������Olѿ 7�g��!{�	I�,K�e��"2�Vv�����b�I��7l�kl�#5�����Yj{�n��r�3ڞ�/�����#�(�э��s������.0Ǹe��y�1N�zG���4@H99 �1~'�f
{�S;�a�.��A��F��y������*�c�Ė�H������z�IXh�o�A��R-�^���,-��|�m���kbL��R\$r�����o�EI>N������#���ֆ{7�Bv��`��j/��u�oB[[��M��⶜�WY��%�,�Ma�Tb�h�*ɖ�Q�O��E��#��8������c��Ô2	����������e,?DHiC��&����R���ώ�ߡ�T���2���o�����ϲn�<㴤��[����i�+T��m�?+U�A~�`]'�dF�}5���v�6�ZR�A�3-Lh�Fߕ{�HL�D4�q�	qO�}�y/��t���q�!L7b|�i7>_��:M��|�Z��Q�Q�b\�*EꊋFP���r��Y]�3W�LAtvt��Ҵyu%q\s��Mo����h��J��L���m�Y�)�FA��[f������9�~���&q[���<�t��틢�\��)4L�|�(.�Ph ����<�N�m$n�Y�7�R|$,O�������-��'Gڡ?����9�����(�+��0�@��9�h��PE��ٸ�:��� �nP�6W3`��)c/���z�����0M���P���ZK��D�sI�R+|��^d=TOk���5h�V.[Lg�CeP6]@v�FU�D�fm0�հ`<z+v��*u|��;-��T>��b�Ҝ��D��+$tsf�A����Q��2.G�����%D"
�.}����UP+r%��f:���@�:����W
b����&��e��.ˡ��e��pG�k�
�|S=����%Q��ڳYSa�D�X�f%�BMW@c��׃��f������N���{\�����n=�"���m�$3ڢ�w��o�����HEz�t��[�
W6H%f��!���?K����y���S[V�=�R�:��.��g������<�=�CJ�7Eʋ��F��L�v�,�Ƴ��ǳ0F3�a]\��l�E���,�(,���O����n�nA�{� #7oL3zާ�o��2f:�6 Q����]:)���{���-�P,v%�c�ϏvFج�.LI�I���R#lɎ]w�D�$�
�2ܴz`V�B.�0K�#z0�8�M��j*�}����W�T._�,:d�©�hsa�����cS[��:t"�b��y��bs!+�A�T�flf��ab7��,vO_	�2��2�Ϫ�<�D��L�LQ�}*����	�a�ls���9i��lA�v�M��9�v�$�N�TR��Rwn}�V"�4n�ڟ0�m�M�#��[���a��ʸ�q۩ҾL��|�-qH|Q�גߠ�M�ɼ?�\���SBEziEnL�w���A�P�D� ��M!�=c,����.C��Pg�9��h3�c��9���}���7%���Jl�!��bT��`垤0��/ǽ2i\0�H?���2^^�8�"r	�+8����{	��K �h9we��e�W��Z�:`�CR���p���i��-�wS<sY/B nIo�w�.��r�7z�:�~��{y��9�]�D@cD����x�Vٓ�*����G���IH#�� �	iT4HT}��譁ᕷ)fn6�j�i�ٞ�)=U�6coI��Ʊr�U�<�n�H蒨е��uhkW��h���c�a�Բ��e5��M,������u��+?����P�Jn8�!�5KmN�����~T��0�4G~��3�~���`{y�JCǕj]fG�dI���eW�d���O�o
-r:�oa�Y<�z��<�/��](Fj�?W^��S��'R�P	�$��N�`V��N�����vu����؁N@��p(i�{�a{�����q9�iYSz�bn�)~4<<� >y���(qx�Ms.�R�X�@n��|�8�V�y|� {jc?�m�@H�p�<��p��Ҿ������ټ �r�N�fIw�4Dh��I���{xܑVt t���~�f5�G�*C���z"\46��h�|Z��f����J�7Q�I�MI��ԧ^�3�E�+T�@��?}��5p��ĉ�w�ل�VQZ�3�9>��9�I�dt�x���-n�(�䉦�߲^�3�&��5!@R�$Q~�/z����_����]y��dQ.�r��[��7Z/�� ���B}�[�,���M���4�ˌ-w�Hez �|{.�V~$[cUBd�xRU�(�P�Ng��L&���V�s���U(ɾ=�ܬ��.ב]rR����#l��15 |ć��,0:CR��Jw���{�����������k�a,���)Ԟ�դ3�OE_�{����X'���أ�S���q��f^�qN͛��J�M,_MJ�#'�x��Z�򏯌�h�j�t)\6y�^vf)�p~�S���Kꩼ�� ʿ��R�
V!ܒnˍ�<#t>�Z�8��v.?c�sM��?�-0	sg9�M�w,\i������J��P��a�O,c$h+'&���R׋ɥ�}w�dc5B��#`C�B�������Eۿ)1�2yͥ��j�Z�
�Đ@�ُ!��j��A�m���`u�4Z�(�g�겁+q(x9^K�u�"ڐ�4��H�R��\ݙN��p�D��H�Ru�<֑"���Z;�۟K����%����B�?�k	cyE_B(0�8��G�h٬9F�Q��I�Aby`��b�"\��,��[ƥO���,zZ���Adk5�i��ѯ��@� ���,o��HV���+���l�TVX{B!�l���6_/�l���N�����Fp$	�2aQ��f���p������`�'2�����ۣ����P&�g���}@H~�V�7�5a'e��҆�
5�4�"	!�����u��-i�4�|�A�5ؒ���t�G�������$���B@���I%����5���hb�6�u��s�:�����Q��(��{�����ٮ������}�e�;[%ah��&���+M�:Kv'!$+�ã�aMov����M"2�AEu��K?`ܒ��(��Td@" �u.Y�.L����9�'L��/�J�v�̓J��P��r\��C�XB$]mE��%||C熩�wz��={���9x�4TԺL	�!�>�.(�oWjLS���'��p�ڃ-x����n�S������#�T�jѴ��+c���ۏYn'��͖��BR�9�=��X{�gNpl=�h��Y��@�0R{+q�g]n��k�k��?`F#hcI-�ǫבݪk�w�Z_Rx�l�H�-j���t�������X��Y�=��������ab�fRZ%[�˿��obs�v���)��FݔZF�[r��0bUh�q[j.�1�f�C�����d�"�4d��	G�{)r�[�K���B���~@���N"�b����DL�k�����������.?��0� ���f�Ɣrh&�5���8��6�s�-�G���%����_�����I�;/�T�3���p�锛k2Ӹ�S���R��sz�r:���|��X����(�8����K��M\�~R�g-��י��,�U�Dn�:�6�ꭐ_�H���]���T�<����#����j5��e��	��Y(5���W�"�')�s��.П�5����r���{"N,����bIzDV�{&1���z>KW�\NV��Y���8�(���'�4nv�b%q=._����Dҝz�D�ͫ�O�(cj4�X��M�#�	
�D�9cR�^{]���l�@�.��q��r`zs��P�
r����) f�&�g�����M'hACW�����X�]�Gfz%��#kE��P��r�w�q	W�Aʽ�9�89�.�O'��=��<��tF&�9��:�a��O�5C������Lʗ,�dߑ2�"�
%1�Yd��Ty�#��NR�(8�_�B��@�R�]i{%�لm�ʺs�~	X/	.Ӡ�����<㔙���%z1����lw���창.Or�K�v�� )�>���Z�.]]��з4@X����u�~@%Gv^�y~a2CLgX��0)�C��P��͜��N��XJ��@q���̓�9�)T�vB�H΋)IwC7�����7!͏�
HY�)J��R�k�L��R��nc",���^�O���M�_��<\����}5�U)�S�w�ٚxv{��4��vB��9�R�{� M�9W!�ᅟY֝c����+IY��r����!)xo1��Ԧ���Ű+���g� �^6Bp����s�] ������ok��*��y���o;�o���ߤ|p��b<��#�H� ��?E�����9�v�s�O����f
�ZFh�RڇR�4&Oƞ<� �%��H�Z}� )�eic���A[���/��A�����K3�e���FV���������K`x��q�]-X���C��+\����g[QJ���]�AOZqEMH��lL���l��vz���G�+^���&�_Ơ�~����R8���4���M�{�g�*HD���v��k5t�1��I�}�7���4_��Cg�a��P� [6$jF�y�s��{�F����q����8�8 cL�ޞ
Mz���-*��<��|� N��U~y������w¦t�4IM��2�bľ镯}��F�]���ܹ̿���1�ڵ�3�*
���:��7C��X�T�˼�:?��ˬ�`��Ԩ>0y."��Z ��˔1X�U��L+�s���o�}�uFv�jƳd���Cg�L�<�̤�ij�����သsΚ�=4�yØ�Ɗ�GL�����i�IA�컂�˚d�37G�pQ�ӭb�WX�W��Xm�t�O��?�����E���D��m���	&��Fg�Ů�M��