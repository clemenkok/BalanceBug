��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d���麍�Ks�%$����+d7��/��������ߔ,���<�E�]��&��z>��>�X�����k�0
��F��p�J,:�D|$�'T*6��v,ֳ`�7J e$���Rv��QL���M'm�l���e��d%����U���Fh�2yRp�.}`˩HD�c
j`͎���7�5G��Ξ@��/6����=;+�Cgt�ܫ����ߥo��yqa�ĝ!�G�F#{5� �E؃��\il����A�E�sƸ��]��i��Y���i���	��'i�6�9U�x� ��n���}FA3�m޿�׹J�g�jM���&ZN�?�Y����#�v+�Pt��Z�a�
��{T��E���cz4G�r�i+���B
�l�������A(-��z%����g��я��_�O������l/�/�,}��S蝅�72~�1P��+�&�K�K�h~8�����X
�*m,NI� g����f�NHu�HBs�*�Hg0���>t�{7)`��A_�&d�P�~Ga���tJ"�6
@�N��++���@����������h��©���I˃d�ϽA��نe,F~z���^\ጒ�\��׹���GXĖ�Fʼ*���-x� I���G�"oA;HΊt�����d��� B>�*4oK��H'U�\`��,�u��'�H$��Yd^Z���r��4weM�̏sr�du>������-���U����GQT�̥����7ҪQχ����h��s(�:��T��Ԁ%:����ɪZ��P ROmJ�m�,'h�td#��d��?���/���j.�N���-J�Xlʯ�����F��3�J�"��km��_������;����1��-Ҡ���f�M�z�^<
㘯
�zOΆ={N��������I���O�o� )6-�vhI��-R�� =�K:����h��M����"�?��>Y�4�yK+,Q0tD����I�{	�L4权}�R�#V�M+|r�k@-���㦘�o`\��On�cWN2b��x�}bQ�G�����
��^H�-3���Np����٘�ceY��?ڷf
�A]��ΐO�?Ȓ`����2r�k�ی�F��!*�5���	�6����9~�CG��O���l��ks��Ȋ�|������yZW�9��wT�Y����-�K4�>�jQ��-�&葅t���u
t�	w�`�xE���-�Ü���d����c�!��.>�QZ\`��
:87I��_��P�Sx�˼ً��MV}rH'�n.~�Cz[�;��/��E�{XBI�y$g�7b
��M�7;;:��φc�/XQ����|	��1��>�G\�,Xf���>gkn��hG7��W���8VR<�����Dnn�m�V�ނ�]҃�MpL;*=YPÎ�䙙�9��P��f��<*�:���x�g;����މk�͑��1�S��{��;2tѓ�n�T9�� �8m69M]"i�A�M���2I�
8�f�w^��{^/e���Ĳ�6����'9 �um�c1V�Tuv�)u-G�S��"�|�֌?f�ݣL�W��	��4�L�B�w�6!�;���-]i�҄k ��Ʈ�V�S `ă���O-F  ���ȫW�/�߶#���k(#���`�W0-\�u��m�y� �1,tH��P.�:�`Fµ�Z�j+�-V�=�����Vr[Eƈ�&��r�C(HڙMo�PK�ƆW���G�}Y3�f����C�dCNN��W�T�� ��t��B����ګ�F���"ayr�IT�K���dd�D/��'��7l,W}9�7��qL`���9̙�&���i"g�4Q�=�~���_n��@�m2G� ���&M�̇nx,��l��[-�xۇ�v�NV=-\zb%�� �죱t�;RX��~>�*�|�Ҝ#���vӨ�q#��[k��E1�.I��Åh|�ʰ�s&��_SՂO(,-�o��5��������!+��־j�,!=�� ��U_�G�CD�b�;"����㏴cĉٚkL�3�f�PjԨ�2G��'	*c���Ab,�-����4�O�)rf"��]��j����e	!4x
dG���F�����D���Ě�_�E��a�� K�T1j��dRm��l`*!̞Y�q��L{O�����	U�� �nFJ1�e����Wx�ki\n�6Rl�=u��2((��4nhкa����z�》#�,f��z�ɥ��إR�����m2��~�(öݛ���*U����Y�>�-��ҌϜȻ}֮e)��?�r���_zt�6��W�r�,���y�h.����ʋ�LI�"&?��V�ftQ����˔ ��j�,�� m��=,���+|a���i�M�]�@���U2��1�b��thS �`��h�Lx�Fߝ�Ǌr��=Ҏ�F���]��75w��
H��/b�v��<!�K����0��(ڙ�CʶSl�c�b ��^d���$&�l3�\����c.&��X+݁�����BH$#�qd�O!Q�[��C����!�����U����`�2��wl<�?:�cB���c�؊C�"rR���=/�>UN�́����Π��%4� sq2��S����X�*��Ht;��N�(nFΐ��}�:��rЅ��]y{O�(%�1m>
�\'�%��L�[����'u���q��Q���	ͧ�P+	e\.����k��('.t�It �&̑�Zc����V��|�zԤNӘ�Y�кL�Mq{̧��N��)�l]���J���};E�:�p�z��"Go�]�ʃ�D�ZY����B�}�����-��W������e�J�"��J8�e� *�h[U��O��w� �i@��æ�\�Y)�����M���$���X�H� �q�r�7Фe��@QQ�-~�嗰�gyޥ[ �r�3�n�P�"�h��^F\����b�����do[z�ž�1���i|ԥ����a���A
���W��/Ԯ�|c�(\,S�||�+�(_��Q�q���4���c74<�T)�1A���T��V�&��RԎs3��/QV���Qױ���hB�5�1�j���R\V���r1oUd���Lv�>�b?��
�L���A����i��7��x�Γ�� +�:q�`HR.��l�� :��Z=sa��6But3���������U�������8ܬƯgc�H��A�6 �\�17w+����8ٓȞ�9fo>�|� 
;��oT�}�o���yP�y'�̀�$��=�1!���7����j��c���kz?M���s ��
�&!D�_PU����ML��U 8�&�� ��ؽ!v�����[����Ma��﨏=�� $t)�u�$�=�����V��Fʭ��0� :>��V���M�?ĵ��q�*�oе�p���W֞7��ca�5YPo�8��L��4m(���,쩩�j7�[��q%�z��6��x���h38��CW��r�)��d��e+n�)I��ޒ,ar�|�F$��j�^�;��B�#e�f�*ݥzE~�dK�n�6����� ��}�E�r�m��>С��`�!�'�@���#[	�<w��߿H�'�@��Az��T��d�s�/���c_�wb	�����H����O���ֳ)� Y�c[aS�]�Я�!x�<���i�g���i�A���F0�Ν�w������p7�:�"f)�}�p����U�F�3d8|�p8)� Tk�Y������ȡ�
� �{7-���8�;a���nV|��DPg
/�''Q��{Nh3#~��-T�]�QZ�Tƪo]�o��^��F�c�A�W��,�_AM�B�'�Z�T |�2[&]��3ǾRo.S��0D��)��v�����*��*ҷ<�vׅ�Q,s�m4"s	�au�����\�m|£$	jJ��Ѧe}:io����( ���W쁅�#h~��ī�^��ęΤ(��_��_G^T�@
=P�!��t�����i'Olp5M��=�C��)WĎ��l��=WbJ��B@���/��)�<X�ݴ8 B����s�E�����)g5��e��,i����(BF�1W�B٩L˓�T�i�+�����l�
��1�D#6���y�Jd�]���}/u�m�D���s���6�LǎM�rr��q�/��Ѳt|F���O�y4wK[�0n�A;�V!��Bu.��Ő�m]�\�Y�OG8
+8a6�I�j�wf����:02-��x��£9>^��0�=FsZ�sYon� ������%���ѥGVH"����Za�K���\�#ڬ���(S�'b����w��4VрE��՟pǢ7dF�~:������+�? dcB�����ة�f�g�����?��Ʒ�+Ǔ�*���asm�����%��RW(ɕ���׼�>DD�(���4B��>z�4���}ኆof�~Q,�K���J���x���|�g�Fݚ����󰮶��p��Xz�v)3[C��A������.��G����2��M���x���j)=�&��2*���2�_�;�6\ѝc������"͖��i���K�YZV�P)������C���:�vΪ�k��f�ݸd��W��h��!W�yr����̏�ld����V�&7�		%�7�����Vy����P��SrԮ(�L��
��1�Jy<�NZ�(��<�u�m|�A�6�پV�BH�I�ĥ=>)t�{�Y�+}b�m�LZ6�ʋF�3�
�"י���n�O��y����oX��+��.��n�4˕���M� i���(��Dv���1�����y�K�f����U��-ΤL�4S*��x5"	��J���ևo�Jj�d7mt�y��]�X���{M���1���!��͛M:P�KΫiy?�ͦ;a�g��{��q�v�n��B~��c깴��$5p��@�ŗ�?�����m��xf�.|��ط*�:k�(ݚ� ��K_�]�ʏCo���;1x����,)�,'���z`�!U�����Zl��a0Z�[S��K~,��jR��_�] ѝ��^<�3joX!дF�,Ӗo	������NL,IHQ)A-��
lb�!��Z����~}���ifR)�{x>�ut��xUe{H�:�Wǻ"(l눑��k�٫<_�vI�C�K#��(�QQ3eM|� �&� T�����kcU����Po�6DK�G�8��w�>��U�Xj툖荰}�M0Jv�>�+���#�Cf[F�!��"s��Z��`��p-Z�N7�]�ʚG{�p��p���dW�\�6�.�ӑ�5�*������+w��K�dF��L� ����`�]�]_�dQJ�h2"u����>1q߀!��Y�޲w��2I�8�g44�))�I��X��F�H	Uo�ě��jV�8I��Y���&�~�;�\T�T�h�FJw	�!����$�6��	�c����:w�uS&��ߌR*5�WB����ʍͳQ)Y�T�A�E�A�Fݥ��x�ྊ���mA�:��ϑ����qW�.OӔw��
�X���E��x���"Q����R����;f�_�2�H�}��BV��1,�,s�����x�����g!S�z&�vO�<n�{��j@��e�kRx��Ѓ"=�I �����%���*�����^.ލ�����V��=+P5Ġr��ߤt~S�"�ͱY.���g�3�N�������+�Q�������i��s����=p˘`]��TP���xӝ���.-�+6�#��9���s�g%vɻ�Fo�;x�� ������
���wqhΞ<�����b5�pP��x9��yo!А��E�|�����@���i�0�'o�o*�eׇ�1��)��!+s�k�ؼ���-���o�K<{� |�D`3��dv	��\��U1�K�ʏ ء�F�	�OO�/�o�I �K��Ǚ���.�?���I54=�:�܋���л�Ú��a�`3�;;gË䰽�f�4� �83܊�� ,f�Yԟ̝?��Q��[o�ß�x��IdXM�S�y�.���#d��&J���}#a*1b{mn� 1,�q��	(��� � ?��i�h�aB��>Dj��?��YN�uR�^�l,T�)�פ��4,�z��$Pe	 �Ğ�O��~sv��`"���GJAd��ܳW����h�`�t�:vgv�#�ޮo�6�t�� �/֐��k�w{�@ԭv�B�CjU���;O�C�_$�3������&�*{������������Ӛ���×���\!�=����v�÷ �������z#�!�#Վ����L�O�{�SB�����+`l���k�Ȍ�9�F Dk�k0b�>������v�0[�%���FU㶃�ē��V�7`�u/����b��¨���V��;	�Xr׀�1B��V�;o�J��V�U��]��9YkC"Ĕ��d�pf3P���"��)���b��WC�	U�ٚ�������0޸��B��@e�������{tm/R L�i/mjI�v0L�P�b���b�s��%@�����X��B���N��ZJ/�R�e�ߌ:����������z�+�l�f(~v�i��0V�$&���N�)���(PI'GI�2��ӟcox������b�
a�`�L��]�E)k�81!B>,�Azh�K�N5�0\�����#{�*^��U@S},|!��G�{�K������_�ۜ�g���4��.:�����1�S_�!X���Wt)�N���S�0f+ HC�AP��9C��ND5}��&���*�S�sROJ��	�;T|4\��2$�:�F��;I��W�wÌ��E�E�P�{�S��g�o
pѐ�pJ�� ?�E0�D�g�
�lę\��%��C5�9��䭉�b��ا�8��+ޑ�z�C}��� ��!U2���:uns�^��;}r�)�m�q��~),6.�!c���	"�Ib���~�!T�@7�I~waXc
fu,�b�BX9
�m#�*i�8v#�"�ҽ�:�>��#�.�V
:#W�`������;�,js�# AcH)�ޚ�
�	=k���%���!�k[���}Y�9��[�/*��!�9����ڜ黧�C%o3"캟m�O���H�#]��Z��v�I(�!��X��*�X>Fp�ނ"�A�;g���s�a����I�����;xȉX��᭷�*� 7�P�pN��p(uN݄ ��O��<
?���M��<�_��,����@�g����W䋈����Z������� <� 2߰8�KSH���g�8+)	�{Lk��=�q���������#]s��L��B�o ��kɋ0�9���T�R�1>8S�f[�r��%��}81\��^i������
������J���(Jw �˅�u��n��d��!	��k�Ⱦ˥�A�.��*���I3�� ߫��J;w�d=�5��p���1�����VĄ`�0'�A�����ߢ�I���D�3��T�3kj_�b;,�eZgc�v���g��vϗU��?v��5��V�|����E��b2���0 Y0RT�DX���w1�Hv[!�2��g�ry�l�B27r��j;����D]t��|tM�LQm�Td]n�F��9ۛ:mJ���͚�څ����ń@��@�8H�9di1��Uǀ��0`��x�a���;9R�Du<�V����
��u��?��4�S:�Ȗw2��"�N�+?�&.t�@'���dq�,�nwm?w˯�L���{sP��m�T'�\	7�˃@��&��s�����E�?<���G�0��Lq7�Ǐ.}1� 4}�qȑ�޾R�+HL3�&�'�a입N���O.�w�Jb��j���l�\ϔ�H��B���~']:�����?j���5�I��>��|~oFC��E�}�%{��d���6�cps �5V�c������d��J�z����[qJ�;��<�/�4��
  e���D�|/<�9q�Y��R4�z��4�EǬMʷ�O����M�S��n�s8tVM-c+�aq*�,����*�]�c[��]�ڛT���p3�\������\��D����T� :�2���ءP�<9�QR�_���]��Kًx�r(A���'^�Ѓ�:�EY �+�C��/�Y����	a�m	�[�}�S[��":�˳���͊z@� "烌����ȧ:o�	4� Ҡ	�V!�I| ���w��|��<O���r�H�}(?K�y!gG�E'�Sl�O�A�J���G�7r�邽���%w�7V��5⛔���Q���ѭfCoG&���JF	�ē��e�B�K�*�:蹬�1�y(3�)K;u��� re�++~���c�6��~	?���ѷ� ���%� dY�\�y�#�pY�ȃ`��N��v5�Rb�9;���D&����!/{X"�s~�	��a_�.����RK���q��Rm�`�����Z	��'>Q��tŁ���/����]��^*g�f��M=�:�u�������R�@J�&�a1�FM�=\�.���O����zS[r�1]�ܕ"��gz�m|8�_rYN�X�+e)U3�����֔~`H5K}�s+!^������aڌU�Ý_a�6��7T��I';dM�M�E��cnEؚ�!�*����"�C�{0?�ǫ���+kO\+��9/:�u���!�t[J�Ɗiq�I/�h ��#�<Ѹ2���~5�m�M�D��K����z���<l�AO\�:`d�~d��v0~��9%��O����cy�����ǵX��(X��Y@|�4D�wj�Z��G����7������x{�t�Ei@��F%����uA~IV#[u>�	Z����Ԣp=��|a���������5�PV�}u�>�Ѓ��=`�2���#�"bX��������y7��yI���g
���{Z�u�� ���؈�cH�Y�����sz�SE����:�<�P�œ>r�J#�6���J����.����l�A���-�IXx���O'� 2�=��y&G͈y��"��ދw�6�-�2h(�>�JQ���`���Ӎ!3���[�D�0�h�k0���ژ�� ��\��=�yzv�!�XL��t	�kU�sqFCM�J����"�p���q�7�Z
��]��C��F�T�����7;ůȒ��g�u���t5ES����R�6����;_������}����� p(؛b�=�]��rh� _r?H��"̈�2Q�e��P�g�Lz���d5�����r��#��s�&$����h��'�KC���Л]<O�c��O,ۥ��i��B6�v�JU�rk�v~�{�{�"H�-D�������+b)��?�t���D�� s�r1��3����!z��|̓ݞs����8ެ�?H"Ve$�\{�OJ���e�ؔ�QuT.�~� �[�˥!��O���5�������`��&�4�a�ȅ�jeT!�)��P�R���
������r��U��{�1�xOt�5�A��vu*.��ݰ��ո�7��8���<p���B�ͣ�����0����Et:���'�d*��h2�HzWzd�$$��R������k!e%T|\�ted�X)����[�iX,�>��it�|����	��O\�;=���vj�8IS^@rC�p����Kk�-���(������v-ԧ�G��#�\&���*K�ԌC}9 ��ʟ�|�p�T9�ڋGS���Y�b@l�bͱ��B��G��M �B+��	t��
����&؜OOk��>����J3"�l��0��Z%e�lb#6��S�X�ixi��F����&��®�
��+�/oq����!$=�D�����B}s�(�g�3��"��%̘s�z)J�ꈔ$��Ҫ����2s�
f�I��E��$���2�y���=�<g��m���J�"�=��i��@�	��B?�JQ�����D�UYk��y��|��#K�h)s�vJyM�
}p���!P��0$E,
������rM0�qr_%̍d��e7
C�r3ʝ���n�XΜd���
��A�`EuJ�6�9�Z�*YBx�� Sö��|�8r{�G�^�� �����ҝ˪�nБ�2Vc�+P�K�cL�U7Ig��I����M�Пatt�6\Un���/X�ƾ��*���/ӼO���Jx�Mh/�Չ�GU�x`�ត�12*,�B�`i�Ī��.{"�:r��n���)�����;�� �_o�C�w��=�6)�Ʃ�]�iA�*��G�]=��ٜ�i��y91	V��M&ϗ�O�DD�|&��%_�����O�Tw��<�ׂw�ӭLx����x��u���V٧ʽ�X�����)}��;l�t�A[��y냰	 yB�Cb�I\?`,N��C̔=���hǼ�����q��+P&�m��O���x8Q��'D\3�Q-���;�%؎ö6[H@خ���&�C��W�ݑ�{�.|w��$�sB�I�V��y�S��;x�r78
Ju�SOn�
�f�1��@iNG��]��|I�e'Ӵ`׬�u�r�S�U�v��G�-_�;��%�!��zD�P�ǚ�	��C�Y%wg�o�9����떚��ǁ���:�5\K�?O�jL���B0���%-= ���w�d�a���rN������฻S��P>0Q����Q�0}�'���l+%)�.��D�
��p�����1�bv�- X��,�>�;�W:�ݍ��{_��#x$S;��O9�^��B��򊵜Ǟd�?����-�SF� )��� V<��XO^�&�I��gc�9	W�1~P1��ј�ތ�V�dlz�;�nH��=�s�7����L��P�����=�řU��!V���+�q2/�kYֈ��m�9��1D?T����FA>j�q)N
�0E>}�+ŐAPs�xy 2;��J�����5`�ֳl%�(�(��he&���b�t��3�ڋYɣᨶ����<
i�gs�t��˳+�rFF�$��% =��nغ����-b=���Iӄs��`or�{��1�X�D���l@dO�uD����'W�7�dfiL+�,��BrH8 ��n�b
�uHBe^�\r`�;���k5u�BRo����L���G������B�{���3c�T�E���7�덐Y+
c{"0��%G x�ۗb2c����s�a�� ��!�1�&yF�����N�Аs-�w�틑�݋��f�wf���}�U�d��-�������E�U5�ؖ�u�����f��Kk�TB�����@�e��������<b�|�U�5Xz<z�c�/ϟ�d7�k�?�Ql9�5%�xàPT\kR�7ͥ���rX�~1P�y?��XP����HcȈF��L�uWmǘ|S"Z4��Ƒ��
�#�ܡ�
2�Q�۽`���H�_�xO7���N���mɆ��+�vv`RD{I�<�l��%�?Hwm9��������!S5t��ob9�P�6R@�8ĴR��4�1<�M*�ԇ�3���C���@F��A��A=i�o�{}�t��EJ0�n���m	ӻKe�����!sF��g��0Hk& ��X.7<� ��{Ϡ�	�s�N:j���U�������X��{l�=ڴ�34Ez��
0�ڐ�ߒ��I֙�I�<Ɉ[�q�	��_��I �����i��~� �)%*u���5휅Gs����X�_M���W��fE�3����R���	�óҗsi38Nw�5�^HZ��R���1i��BC}}��OOk�~y�sf���@q��lQk&�UZY�����Ț�3LZbf�J��zf
��t�c�'U���#Oe�K�1�Pd^qG��[�U���v��G�ĭC�,�u�2<6�v��o�h�4���<�nW����
�n�a��~�+�e느b�7Z���ΪF�Y��Z������*E8u�S{i��ש�͒[�YwLM.q�-���ᘰ1¼�����3�_��O�Y^�	E�m�.����K�=8�.9�����g�1C�{����q.
e�L��Q=mxi�
�DX!7'˄���>�^y$t��y<|FZ]��i�,��-B��'���6��؂V��(�*�9�ܨg�*��n_�ؚ>���ػT-���@�S��?z*�)�pݦ�U���eD�]>&������hw�W4��[�b'^=��	@%eQֲ�)N�L����2��{:��]�s���
��&Fۢ�H��O�T)���|4�k��d��iQ��� L��2��;����h)g���]+���/W��=R���ފu7[�`}U༫EG���<Z�$K���f�1F�Ͽg�f�<l�6M�cH�\�ވ����Rv�:Z�jb�Pu�aH�=���p!�cm��8.7�Gj���.�\A|d�;��m��R��@�G�x��s��@7Tx��Hl��U�+y�ߊ��3CT��z��^NhQjeM�H2���V�o�,�{��/����#'}�n����O;k4�%�����uT�@�ehV��cx��Q�3�ui�dP��V�r��ch7Z����Ԝ�r�����|�pUg���:����W��kDR�F۴�];B��#�T+V���Y��nS�^�(�t��|&���Ӗ��H)���Gfy��Nޏ�1F��{v�������BP��*ھ�1Xuߤ��rW8��o��eM����h�*�]����ƞ��_=�t�e�������p�������4]�sS �G�0ͱ�[��P��j�#���ʐI@���RǍ0�H�ʙ�{^�MZ�i�N#u��)�m"u��!�c��������dn���c�{��*}y6�-P��}���*���f�p�����q���Ʊ��*�?\Ϯ�L�����?%tmD����H�B����Jh����0��.7�������q7^ �fd��4�쩲��P�9K�z��T�ԫFfw�m�AyW�jG��h��]��K`$�I�9�#���~�T�,�E�GÄF�'�Z6���S�E $���CV"{6�ʘzNR?�[~�+��46��0�%{.LH32/@�l��v�38�Gm>�~�f�q��c��.�|Arxr�gq3m� �;�a�^�5�� �z��YW�Z��5�W#c*=
�����7t!T���"� �������x�*�2�ڪf�$\�,�O����$E�{q|�l�k+jf�yNҪE$�&���>倆�����S����)Z����;����Zg^�5���RD��,m����{�R��!�����![˵0Vh�6|m�+�C��\�[p�q��DTߔr�^��F>�{6K�#eD�q4�73�\[L5�i�w
�&�����m<!�E��V1��HT�T<���]�lVױ���ah:r+�.��,O��ZfDn|A���������;)Ϩ�`(J������/ʢ�X2����S�g��l��h�U]�Y<<:��H�m	s�t�
�*C��<�˱�S?�/y�0���$��$l�]�4W6R���v������tŻ�ݥ���E��F1S��R�K����߅/��L�r�i;�Wcv]��u$J�b�juD�1���3�1ŋ+�v�RH���F���3�j�~T�Qn����#��pr4K]��� R.�v��iF);��,m��=өG�����H�n�;r)F�d����ŸmIH��0!���ߡW�ra7�hj����	:ƽ�w"��N�\C����*�x�o��n�!����p<> ��4��~W`*$Ъ{�U�k�+P��)��WȒy5���5w|�[�Q8�d����p�M��W�l,����L^��V�^���Ϡx�C� ��o$%Pی<�`a�Ӌ�:K��T���om��ܠ�i���?�%���|�����J�[N�XC�(f��K�R[X8-܉Mc�/gK�+�,��Xf��<�,����<7-�Z�>�������S�~���
�����\U4f��DP7�����'$|�˶Mʙ�_�$��c��+�<���T�5j6�iʂoo��S���>[���j3��D+�
���+V���/M�\�+4{O��\f#�õ��A�$(6EM�]� �\�X�muf�	�+8`i�9F����]�ܕz�(,��waHq2B6��L�P�6>�-�d�Xa�:c����(v�]+,�R�n,�gf�m�xDdRP��7�'�+u���h��s�k_��Ɯ�^��^�"��0c��b��Kഽ���>E��QJ/���C����q+�Iƭ0@&`���K���XY>�%�^��=����bL�XU�p���F�Q6`��f��ޛ�V�1���'S�CFH��+6�����D�F&����rV6(rv�'�u	̜���Dd�X-rSL���?����l ����W{�z��?Κ�����tG�����N�E^�G?��^]I^٧�5��Iq�f�n�6�5�XAm�mbMe��7��X5I~��g!�������ҿ���bJ�h#Q�Ʉ�WIB��h?#�5��c�H�~]tA�,��\�Z�9�P�ǯ{S��=	�s��0$	���Rk.�z�d�S��`(Ņ)F&1O�T��a%[��џ�wZO��*4���	����sC�J]��=��VL�M}ɐ@�p�A����]j �JӘ�$�ھ{�H���k ���j���7:}&�3��� yf�����[;F��2Ƣ���o\���F
=�N-�ۢ����)D�:RW
��JJ�]p��˝=�&C �頊�ء�1�֩�ݳ� �m[�=T�om�_P�[�cլ�w������9�qr� ���<j"�/�]ah)ٱ��A\�g6ޥrm3�<��/�y|le�$ܔ���~Q
������l�� u�
���}K����H$�&Z��(���ɨ�0��)��.O-�iQ�:�͘�xY��.2G��O�}���HK2N���	+�(=���a��i�t;����	�$���x�O!�����6�rQ�0s
���ۯT�f�C�8B�i2�!p�sN�z��Fɰa�<���HO{���W����Վ������i���}�P)�ִ�aI�G��A�ʋvC������ɫ��8H_�P���[�	�7}n*f.)g�����*��o�5���4�쇮,*Br�����tv�I^W�E"j� ����.��1	9�[� <%���F��"�;����ɜRO�7�^_/�j��<�+�/���UKU�8T����o��Y!a�(9D��6Kp�	 I��>΅��C�b�u���#�<(�����!��䀗a��B\!:��M�^��}�.�W��˘��k�[]8�)d3���5�l��yF	�Ui�r�aaWN�}�m(J(��@��4%���wf���Ls�L�>�<��϶���韑�-�ܞAш�a�7��:ń� �~�σ4V��-�҂|g��e��H:��8g��I�f��h[4%灯��j����nf�L���Y�����|�N�=I��NPq�r
��tЉ;
t.�D�v���dT�}�^{y�Q:g��mr��)a�j̤�'���務3�X$� �W#��YE��lᆖ���	mQujo�;�˚go�����k�*6|�oؠ��h�y@ ���w@�j�y�q�'��^>��ә��{��Ϋ@��A�gK|Q@��4U|tC���Ț���!�Xf[,]���}��7��k��?�sm�Q�-U�ө��Bg���%�GZYf���bv��C8\Ʀ����� ��cwBj�K*|)��.8��p#�]����i�&>����!ē�4���5�^XY�櫡�#Eǥe�s�#cy��*��R���y
Er.�H���3_/j`HKg~���ݯv���UO�����]�#dUUpr�-d�kʼ	��PA҃H\�;��I�#m����U� ,"$�����i��ǮM|��UJ�w�y�(�젯q�8ИL� ��s�&� ��k��'��F�~��C�������V:�X���	��Q�7�m��ݲ���Ղ�eQ�CʜC��5 ��e��yk���a"�U�L���D��d�q9�o�k2��yCѦt����(*�I�`~tRHbBڱ��gñ�)�pqx��2�y�8�)�o�X;�
�5��Q�Kt�\/��7�s;��W�/jZ�F���~i-.��xo椞P��d���
U"�A�h-�)'�h�tD%i��ڱP�}�7kT.���<�$�m�q� w����F�l������	�1��P2CuWEi؛�E��r�����I��|�P�I�Q���
πƱ��E��Xhu��K��Z�ŝP�e�h-vg�ph��A��	"';�)�Q��#$�V�(��͉���E���5㌐�F$a��e�*F���V�*�����03���Og�s���l��p'9ҫ��C$=d���T� נ6CJ�r�2W�� \��Y	�l����c����;�| ���&<�K���O�1'�b��N�wd�"��hq�ȴ�/��y�o�'�_���Z�K�-��0����Rxg���(�����*�j�"� 6�#�H��>���	��"U���*������� 5}�.��ւ#����3�<���9�P�{�V��m��R�s�WЩ�zo�U�~�R�xP�.&C�N�-�y����~(��k���L�z3gN�%�.27#C-=oZ7�Vk��s�<�j�v.��;vs�2��Զ�ɬ��)8-�Hv�J3��{��,Wt���qԬ�[���c|E5����G.�n�F��Eg��6u'WD��埍�Pk>�Cה�[S��W��XIJu�̅U�.S�/�ͷ.ь)N�^�B��_���W��T�4d�md)�")	�7�q�(@e�Er�$bTVRGc�[*�q�.�ܗV����$iyV����kࡷm�m�r'X���v����8�jvЪĥ{��R���g#.1����!C�_>T~Ѱ�?D���<���Wd�H4�ñ�v�Z�b<:�w�e������jW�JT
�X��#$c�"�@>G����
�����)&kL+�zS��7*�6�L�l�����%�`���=]6ctM�p区�C1��J�ݙ�N�P
�f_��PU�n��y���A<�Z-8��o�J�t7�J�|�1.��`I�[b�� o� t�6�{�&5b��{�/���T����<_�\����y�QW�V�2�_����k��]Z��1��gU.��\TK����`�M���1B�c�JW��LV��Eb%�֨�`����S7I���݄%��.��p�c��/f� �DZ���E�O�zHY"�i8W:�p�\C�)��_�	p���o��#���C�G[E^U���a~���Y�sr�1 O۰�>d��$�Bnc����B�uξ|����ج&�t!�4W0?�����k����A�A��OF����-�7��ߪ�F<�7(�:��/�/	������6�gy�,��|\��ڥ�5�v)�vfD��� W�E �c�����O��0gXhC{����u$r��4�d$H���a8j���鑜K9wC�� ��[[/.������^�,|�.H�43�?@}Β��]�%=cXՒ1Yf����T�66h��5�l���dĊ�eU˸�@�N�Ƕ St��n�J��: K��P>[��'�ꪥuGEZEc`��hPo������ƾ�-� �(+�������eg`MN����8���(1J���F�L)�_�N�7��Ml^������%J�,"��h1�&�I4��F �M����(�5G�j���է�>�]��98i��68����n�p���V���w�{ɢ���A�j�a@�"�

�d����b�j�;�p����GG7����b]>���.��+K�N��OS�� &.x�-�7o���C�La��R�����u�z�'�LQP�F�d$�z��h���KUaR�~�!q�{Gy�ot�����tx`i����76DeYR����R�f��G���f�U�J8eeR9��F�?;tY���`��3���>H���Uح֫N�2c��8s�sޑ�htN�2e�5�Q�Q�9Z{��샨"�! >��XBLS}GȊ�N�-R�6�q��Gx��"OHԉ1=����~�.�w��-�7�k���է�a����=Qh��Rнoc�J�S?�M)e?�ЦFz�e��UJK����W�9q �h��kx�IOE�Tcژ6���9���>�<T�tr8λ|(��RMJ�G��d���������b`�r�m���p�Tl�i!IGO�����qd�kB�7���I�63lLx;����dJFˡ��^�����
o�Aa�/�l�l�<.T�G�V�v�ZP����ZZ٣Z6,�e�I�wElNo�.�;�� �9�)��RǅM-d��][9A��V��~�@�{\�aX��҇d0��v��'9?�pF��D7�ny�-��)k_1R�^�Z
<�����f�fޙ'Ŏ�r@��W6p��o(p�(�����]�����P�Q{���!y�c���RTݗR�tF�v�P;8Z]?[#��K.�i��}3dOC�u����
���is]�m�$@���<��ȋ[���o�C�����̩�5
Ntr�ٲ���X�uI��E��[�A":��#�33g��%�M��#�i/=�(�m�S��t\a0n39-�\�"y��b��
�g���u��ă��_��$�����I3#�I��aI�L!]�4�yuC���o]�)�A:V'�1z�����6T������
CKi�����D�B0�xIp4|�g� S��j�-�!���6!x̻��L�#�p�C!�xЌ�ҋJ��%>^��G>�}����f�?B��b7q3�)���u!U2t�4! S/����ט�MV�0�M�A���
:�dS�Tչ�X�z��H���p�7��7��T�LnW3љ��)6DD-Gm|�T_�˝���;�i"�I�R�uЇ{��bG�������uUO	5Zi���JF.��&C�Ib�z���˱ܛ**=K����h[�KԂ��k8P��M��~���&|������qP�WHóNt�|�Ѵ8oR��{�m? YE֨;�%�ٵ4K��,���n�:�"�c�^��M㐱��b�<��ȼHgm�T�������p7�s��Cڟ�b�`��f����$,��l�܄�L+����E��h/�Pa�Q�^�p���d�a��Lp��:Z��
��=Ǫ'�~Ƨ��/"�+����{tKQ(�<Q�h�W�lݙ������E�ߣ���8�C��N��&k�[=���[�����Q��Q�!�cx�x��?P�W��S��(�̇�蔫��(�0�4?�;1�?��a� =�}�،v>���jS��g�PW��o���;���foM���דڬRgqF§�m6E��` �[�)2�k�v��q�It�~� 1��>|.���p��o��#��f��q����@��i�����|P��i+���EBV9Lۛ�ۧ���`�@����}��i1��ݫ�K��*�V��RR��QR�|_��Sy"W͸���4�S�L�oyj*�Fx�2>:=��+;4rv��3��~�
�bg�+�yi��ɻ`kq���ddNI���AE��| �C�-�Ob��-Jж	܅��=O�"���%��F<[dZ�X
��}x$f�&NF��gV/���A���`rQW� S9�#e�$&�@y�Bm[}h��;!^�a����H����E
����5���G>#�YN�`��a�������	��m��w�/�:������T�D��F�cS�z�$�� ^_������0�xXg����*�jI�jǯ��έ��UGAH\x�Y�]>e٪�<�8��߄L��
w�Yx�ሰ���R!�i����`�nmK�0�@��1I�W��>�@Z�����к��b��#w��ٯ�A#��M̹='8sz���D$�O���\�@�=���)�I�,1�h�����ɘR7��U�/_2�Dy-����^^L�r�~��Yh ٚ-�9�z����1��b�#i����͜p[~3&o����k=�$�i���� �T��c�ɴ��u��X�D9��C�m�#�w4���|LT8��`x��b�T�U7�&C2�錈�fuk�D����%�$z6e)��k���$�zq���������^�=(���r��A]u��_�⿚~��O��&k�,�������D�Rb`��m�=(V�v��^��B1jP��p|Sb�R����%���t�S���o/�䵦�4�I�ja~+>�D�eM���q"Z�Z����$��ڱ�NI�" ��Y�Z�$��F��N�6�Ԝ��o2o"�������qz�jV��+����t���$->ZO��ͥ�[��UZm
+G�����R�.�#����f�.�6;Ff?��ϐ咃�w�11�ϐ�0:�tmw�%)g]�'��OJ�����:�*����2$݄J�yUA%LG�O.�I�:���:����Y
��I7m���"'���?�/��$y�Y9Ť�C�l|&����Ԝ�{�QCL]�F�x�h�V7�jȊ�dKǻ)bU[��\����e�t�V�9�Nt�Hyj t��#όP���l??����iT�RT��Z��d�������<4`� �i��X)�T�"�ڦ����Ҕ�tvi���)�$d��qs�e�ܺ#��AQ���ð��kl]FlpĔT���a�S-�U��E�>���H�2�	|9r�v�&�X�W�'���@L�ï~�و��O����L���W�R4)!��&"�T�OOj`b'Y�o���?��Vźd.E��o��]J�j�'ӊQ`�'p�	#�T�&B'�4��^�Y�g������v$�S�爠�
X�uЪ4�ߴ"�����p��t.?'��Q���a��a��6�^	�h��y#�ܼ���N<;w�jfB%�Qtjq������v�3e�������d���D)�X��U�]������w	ֲ�9��c$ޜ����������z9K����oc�_Z���)߿'�nLN���i��k_*f�3�������٧s����4IM���J�����HXڻ��/�H��;���hH���ۄ?šy�/��K��q�s!q,W*qR�4����� P���J~?����d����0������_F�pm����m����U+�[�x˒ �Kv@�7�C�谬Gc��urct��:��'�qhC�}�F��mZ�
*r�T��b����e+���R�7��h�8����N:O�
ؘ�LM馣�̘,���� ���ht�.�%��f�gl�2
)>���v̜�e�΅���fՒV�H�(]Q����&�n9��p	�;��!4�r�~Q�'m^'����x/�J�2Ȥ������ �ǩF�ϯ�_FrRF��3���&�� ��I�I,�;ޟ=�HQN��(0��C���9ϻqnujcDH�k���]/�Ӄ!�gr�H͊VVJܱ�r'ʮ%�+`�(3!��B�L�Lx�:�X� ZW~��+��>�_GO2,��Ơ���YL���6����U۝uc9N��'���&1K5$�M=�2~ Ŷz&7��heA�O���T���lF?��PU��z��H�2*���(:���-p-�Ag��P��l4��E��d5�X�L�E�������x���3�p��5�*Do�z�f�ͽ�o���:�hf5ho�#����@�����e3;6�Չ��S���z�����0^Bp��V��V��xP9�b'��/�x�]�_�.�yIRm�F"Ř�~u����d� h���cX��5�)��M2� ����9[v�Jkj�Wt$�Q(ӄ��V)[�3��o�`O}�𮋪�_��*�-����:�=���]{tF����C�a�F��p�����I��?>�k�O�����Qu۫B���.a�=����j�����N�Ώ�����c�	�`/��+�Y�3��h�ޑ�sl��5m
�Xr��� �s?��!I��M�����i�����ϓݔ��a��ީ�ta������52-� �CC8�Uj�7�"���v30��>-�]�h����H
��r! p��3�@P��W�Y/s����ҧ;8�V0k �+8:Sf���EL}-��L�X����=�e�;+��|��������Gc���z����[����l��v�^/�����M��v�xq��9�	������P���96oҞ���Dք������#��g�����Ζ�-���	ND�0�o����'��V���D&���D�:0<4%������۲@�rec�2�,sK׃u@�I���%]�P�����S����@;��E�٦� �we(���$DBa�<ۈ���ݕB�|h��G�p��A^%�g����r&!S��<�SK��׵�te�B,�;Q�GE����A8�Cp���2L�`S|;d�@�o�!U�K��E���Ź:��b|�1o�Qv��у^j�/���Ll.!I���n�K�Z����[�왇�$d(2�D�G45Y���W���xٙ9���.[��Ұ��tj�Q��I�̶�:��
�'K�uSJ�m�	�4�u�-a���h�hpb<���k"���5h�'�R�Ǐ�O_���-4酛�&��JpKc T�n���m?1/�.�D�d�2�r�@g�v�ǟ�e�T* >�^7\��&��PԬ�ˈݫ��7,���{vw��;%���!i��I��`���s��S�����c��c#��1L���<�Rl[K޵�q�ɒ�e��q�N���m�8�J��S{�k�8����D*'��s��d��J̦p\�mR��QbVH��g��iZ���d�&�oT¥Es<���/B���<�\��$�b �U�*W߶��"e��=t�
�����&��!�َ=F�E}M���C��l�#�bm��Er��R&�g ����i�"�*����@ ��m���|S�o��!�#�o뼃�v��	�0=���W�BR��d�DQ�l���+�s�y��&)ì��T��1O�e��8\F�j\��ȉVDS-|?��	5�.b�GP������VE�R��6(��)3.1vʁ���E6NgS�0%�X4����;����SQE����r��������B{?x���
"	�#�Tb�y�N|	�ukY]�z���k�^̞@���{�n������; �K���U���G^����C__k5d;zK��Ȑ�'tn��=�|�������X��2�Q��Ii�:&n�n��K8�,�
'������ֳ���`�dP�\-�R±q"����jqZڍ�j[:�P!���ar����LS��2���nƗ%�f]��u��0�p�����I�[������D�B:h�R��P�M����j'��A��w,,R�-��%1��S�q:m������ �����ƕc�6��I�'񾎵��i�E� *�d��'@2Qx�Hnߟ�}��x!�T��_����$ɇ!�`g�����h�(1!f�dL��z֨k��Ոzdhx������/~�&�ȹ^'��b@E��]���G��]MxC�B_�}�m(���)���+cB��E��U��n�aG48Y'8|�)��ۼ�mM
��(f�bt���n����s����PT��3�ʳ���k��#��1��]U �0m��i�@����p� �-�#��:�W�{����&umtr�W�Y|�����Ѭ�;oL�)�W���CE,�Ůj��yΕL������y l�B�P��K>G��_��ݫSƤ��d+ь�s�{шĳ�}��׍�A�4�U�ww�@����'(�*B0\�=��D� �jweWLC6���)�&M�*��?��B�Nۈ҄���C^��M�'�ā��ZM�>��%e(��/p]�m�0,�H��օ�ܜ�c��hyW�-�<ۼ����^���k�K�+>)���a�`.:0�rV�s��̉��^!F���S�Z�:(��|�![�T����L��t�7�X��������Mo�$te��~GL<�[q�|f.��\ぴcÒ��Z�;$FM�JQ�z�f�8�,%h@�[6�����\ȕ�24l��<G:��R*E43r��p���,�Iv6zZi�m���P� cË��{�����x#7�E{Ns!rqGԓ���R�����+�'���vhWƠ�e�N���\99ֆ'���]ש«H̤�5���l�v:xcC�.i��Caq�vH l_g�:��W�uN�H�=	��~`h"��/���qWY�����OcB�9��Ը_�R�X�~ەf�@s��Y,�2D�3�Of<���,�%d؊��@��}�m�av�ܒ�blPl�M�YPqT�;	Խ\�[ߣ,���՛���yԇ�d�$]N����UB���76�GAxċ����l�צ�M9�Td,W��z�6�M��~*!/��P���ֹ�r�� �!�vA���=N7+�Q�9~#�:X ��\�d@e�!˥��}ů�y���Ʊ��V�tTPA�8=�A& #�x�g~l���t?T��]H�����w%Q`���[���s>2Ex��K	��u���	T���^~ɦJe��¦���<����{'��j��j��BQ�`��G�7؊�@=�,�����v)'�4���O��5�H�>J<
5�A��В �	�8(lR�a���Y'���H<��X ��~�>��rgÐ&��tb�Ǟ4�+� t�7+Tn��!�vk�6��dkc�ӻ���R�b+9�4]k�t?�GʨE�����)�M?J~	~^Jo�����4�R-|Ew+�_q5����0�Ssc뿟&8�$� +��~��'�H�Ѡ5f�\FR��L�ɖ�8�=��n4"$�JI���	w�gk_YH����$[ЇT��\�(�WxH�#���6���ɚF�il���q��1ha5~j��B���������I2��������>���B�wF��R�w��D�,M&+ ���_�Ϗ�e�ظM,������P��L�,��lb��3�L�@C�<��[�\�5�z�0�?�I}q�4�[e@��'��@4�l�O��I"z���ZG�ۂ�I��U	�����	�5V���ܹ�a �`C�(J{<��
_���o�1��īe�]����1㌖��.��whO�($)��ϔ�F	�B	V�-�0<t=7���"/���c�����"��Rʓ������}��VnA�P�$����dvkR)�<�>��E�1y�:]�g+j+R��Zc�?���Ԅ���j�����5�;���b�I>��:�0P��N��~|�p�%�&4�sp����R��D"�t�8�#	$E��ʕ��T����j<d�������:i���=��,$���F#o�`&ć���XR��p����?!��t#�-	�Mu��cWL)\/,h�e�W0�i��Fو7�'�ٔ�#爵~����:�RA��%��Nw<����T�E��#8��ʙ%� !�!A�)��J:ۼDc:��-\�~�)�p4	�5�R���<!��h=uru��qw���a�ƪ�Fe���t��u(l,XH�\���,�u�YԺr�/�R�;1/ԟ��a#]�Qʻ���(�bPD���Tf�h��\*�И4yoiE���R��j�o�4��Tf��}���J1�+������p*��lR鼒2�0�P ��R���d�i�`���3iC���1�l^E���6b�YJ�S9��6��˸����%3i[�(��f��82���n�gۣU��6�vc-Qcī��g�3���	vp�1���R�X䗳6��Ȋ9�mՍ�����ho�B���@Gg��T��0=���b�_Z�Iu�<��!S8�nB��c��֤M����d�8�0$J�$I
��-�Y:�RI�Eqd�l��֙�aҕ\jOU����L3�R��VHFW�&�9TT
����b���8w��yGw�� ���N��:��9Q؞~J��OO̓�& �A�����R���@��/:�	m�l�'���!�P�$:�,�żU!��` ��)�V�k#F 3�|	EuDFO$/�Ԥ.Ђ:%Ρ�jH4����@L����ǻ��{-��dM�Z��I>��f�;`v��p�R�=���Jč�2�,�0�*�@�Y����'��6�-��;ʢZ�%fGD)�*�Y}��Mf��a���e��9���f)=)T�f� �,���k�t#[�A���G͞���� ����������B��ej��d��%�ۻZL3��r�r�ܙ�?-y�o�]R�uʿ����Z���#�.��qQ�x��)u��m��FĽ]oT*�íj���K��^��	���'� WD7�H�ĺT@�y�U�i(�FBR���iC	$�b���Ec��XedI�	o������
�K��	��*+/4�:��H�Qm��i�hKX|�n�9p�8ދ~�����J�� D̢~�h������2/N�~!�.��#��Y���'���N���(�#z/>h`u*p�m2�w��v��gB�8&��Ϛ� �g#jm��}k��bs�¬�k���&��s��c��UlջK#�Dcg_$�n��p�������E��K'G��7�0��HG&k���P�94ek���fWk�k�*��_jE��~JcT���<_���A='|�=<�6��Db�����HL"��&��.�ڗ���UQ]�S�g�΍��a��\�X<�8w�.��m��ς��Wݗ.yH�^�h�lA�^��ܩX�e���.��'͸��r]d� Xak�eq�2i�[�Ð�)���Z��l��Š�$ѝ�R�#ݕ��	X���H�V\�#�v�u/��k��O��9&ϟ.��jW��2�d�?��W��vp��a�uLӤ�_��F���$&����0>�A��p����{�B�����5i1�yi��_�Iy��C����ZLÖe�9�� ����[�a�Nn��X�nP��=����0x�Oᄃx��	��G?0Y(�e��">��w��`X��h>Ƹ6d@��ZY����k˜hmW .��;�'���6���銮��)��2�T�������.��������?�!j#��,�kHB�%and+�qW���a������5����$磏�1�SU5�������m��[�$*+����1� k��+�Z<��M_#����j��?Ë�:,��*��Z������hA���M�i��{͗^�8w��3k�:�9�1�|F�Q�o��-��2?E�q�����ݯ�\�u���L�s��'�A�T9��1q�5�{��G���"��0DK�Ӕ�!� ��S�>�7�<�-�X!����(��xvIݱ"�Z��k��a�|M�7]Il�=��ԏ���^�?����A6��(��!׵d	���k3?L(t����8�\Y��;���8���9f-��u����S\#�,���lEٗ&�#9�U8��:O� X
ܹ|vƁ��W>I�-�Z�j>% ��xX|R��HnI�RI�.�ټ����F|��&e�����&,�������O��5A�R��&�Je�V�͡奼��}�UH���|:�V���qs{49�>�+&~Y"\:���M��o���s���٠�g��T���-��)j՛�BY��c��1E���9NE�:kM]Q�J��������z1�a�t ^O�hVIvqG3D����J�	��O̴	����
1=�i��D�#�ʶ� ���)DK�>4of���~�VV��ە��H5k#mHҸe�Z�BnU-�E�h|��������:J������-bWϙ��ʏld�Z�]p��/	��T!�[Ϩ��h����<W�d�i�YŚ�|sA�O��A����l�R�o�[G�UFh;�D�- 5'�c��~{�)�,r�v���%�ѹ���u>�~�}���/H���c�֓��=c��o�4m�(��+���[�����R.������z���mEƊ��d�Q��S!����D�]��ǁe��k�TaX1���<IW�:*�h����)/�s��M�VG��z׀ώ o�`u���	a��_6����A���y�,���E��q���P	��"2�v_�	�� f&`���Ea}3�Q0��7�C�۠��k�Rh��Fc�������m#��*C���'��9�����1G��)+B�u!�K�x^>�l�����7��/	լ/SĨ��˺�S9��*��zu����1j���iM 3Ix���gny�G�l/?�!��	���so����)�0�O�dy9St�>�N���e�"�L�v�k�谌t�7�As��`��#3UKɘr�C���w�;F�`��k�tՉ��ׂ�r�o*�l��� @�d���2~`e]�z��_Ǜ��M�h��&�Y�1v}*�}�D��q��o���9�g���9��${���[ڴ�/��
ǣ[�F���d��5cI��e�@��@ ��y�\ϰ\�W������1��M�z�����Bh�}6�ᅆL�$�?��Y4ѩs�b/m8S����m���o7��� � W����
TJ��i�a�^Su8?iz�>�=@�r�(�:(�����q��JQ���܄c6�QZ��ѽ����kɅZT}#��?S���n������ql!!p��w�V\p�J�3URfA\� ���7��Q��f�U�}��tP�:�Q���0�����ò��73�L�N'C5dc.<���[��A�8���0�E�I��ue}?�I�8!8E�f��l�)���ۍ������A� d,��f�!�dS�-,�;~��9�{X|s��E]9��2G������r>K>=FҪu�^z��_�G�+6����%���'�.�g��M'�3k�����U;(�O��;��G�F��<�4��_ Bc�%�>����CJoͰur�H�U|?��WB~��,D��2c|#i~U����d)Q�L�{ͫ���TPT�Z��m��LCӾذ�;�+69�c�6"�����q���˵D�#���ԝt+
��/�,Q�
o�s_��%b�����c]ؐ¶�!AF'��_�~��`n!�M�>��F��<y�}�]�!4��mO\��uN�nT�_<%��6x[��.�KQm+?Q���	d�Ť(08�������V|��B�Gn���,pm���Z�͘�R��l3?�Pt�볼��oŝ��q��d*P�t�g��Wo�F�THf�E�M]��t��J��fc҇�J��r�(2�{@�=>�}�����t��|ԗ���Ί�B'��3i��=�7��0��С�nME�|�@�T���Ρ/?b>��N�Ҩ-���v7���;>�&)��݅��LQ�4<��ꣽl�F�rNɶ�Ѻ%����`23�Oq���gA���b�W�\a���P+��C��ƨ���<�ڠ�PU��41�P���.I\J̞����L	�s��V�r�z�QG�(�������R?���iO����/��P6�3�i������G��������u��n�s�:��ּ~#�2�, &�+`����(��p�u��)�_�7�:�O��
O �cl_����e��/QQ���|�s�K�?���l�bNƩr-rMn�KB�Q����
j���_v�^���:��{+�`�↔%U��;�h�c��`;DZ&R �@�8y��=X9���[k���h۵�]M1��,ד�����z��6<��﫭��tr7J ֢��>&���L	7�A�����5.sv`C
�ֲ,Q3���?-�Fћ�b�9W�l�!Gp=��-���7g�'�a�+w�1���1~�+^����Fx^�I�.�S��-%Я��.)��V����{"�^Z̜�Dh��4kH:C�.���>�n�E�u�[ҰY1�×��.���R�2r�����@ը�?\R.N�H:S�ަ#m�Q�ޢW
ғ����{ѥ�J9�Ȑ(�C\1�^(���\�LV;��dq��	Es��#N��DP�ӣ,��qY�9��X�E:�,���0G͹����I�Y{,��頩K����8�^Dc�p�����V̳jkgp�p����5c�"�| �g�峼�]��+�Y��R�z����C���9���7@G�f�x6�t�2�Z�0���_q��U��H���Mΐ]����)�14��k�R�lb�5�_^��Xx�m�S�f!�R��B�^Noٶm����&�~v���H{x�1�& ������Xh51��N��tz:�_�[3s�&j\X���[e���e�m�ؠ�S�9;n��Ge���>���6����z��&�߀x���
�验�RD�)Q�+~��X�<��p�9*��)��zy���/��»i5�7>�k1��@���✃|mj���B�V���@�Nm6�`m��h��X�	n攓To*�eD����(0���Zu��'"�Ȕp��8�ىpwD��59�q��G~��l�cO�ak�i��B1�����Y �;�N��kҼ�o�"��eM��l�}�U9�!��z%�)���i�1�|a�SJ�|���Ŏ��D�쀉
v��Ek[t�\ҧ�-�8���RW:�����x�۞�6y�{P3h�|f�Z�2�<�ѿ�G2~��|�^ 0�?i	zVi-���-2 �2W$�������=����)$t�����?��ǟ������0pF�l�IX.�E�����ffa]�)\���}D�H���������2GFf�;?Ʈ�K\�5:������H��K�3'�����ҫr�;�mD����^G?9�}5Ǟhޡqݰ+��!�I< �BQ�,Ov���kQ�_��%/�
R2�ӂy����R���i�O���1xuċWK�K�
=㖻�����X��l����N�vU�Dt,����ȩ�H�A������5�}>�[ef�����T�]�L����q�iK�Y�ыbw��Y�2��Y�=��1�r�{ϡ�Jhw��v���rA*� �)�h�M Zh�(�ZC�T� T� �:Y���	�(��tt[�
�W�%��#7�,���\ה�A��ۗ�_7�˄�x$��^�%
�P�q�U�qވ9�l�����J��8�X�ՂA�riZ���p"�ߐ�h�.�n�d�$�q�үr��<�W�IQ`�_6��A�{��6|��,U�1�O:B��}aY��.���AC���G|�h#h����k0��t������O�4��TQ�7;T��5�/M�����m�f��:zj�3V��c�A��H�S�+yr�G���vfV�'z!���3A�$�mz��`�U�d��%�SO���v;A��6�.t�`:��a���99��]l�N�Z���[N�r�T� ���?gg"#�������$�W�4_v��cul�}k�Q�=MR���#3��.\�*�_�-#�p/�e��4)r�bV��<��j��Cw%W�r$#�P�Z}��ڟ��
d	]t�h���#���OƱ���CY��9g�3NS�}Dof���7��6k�8uT!��j�>+�����vN���PӁҎzY�ㄟ�Ϥ�H����p&���EO�L�P!H�l�2Y=�Q�R��B��[;G��>�i.������-�B���h����.��t鴩�[�N�;�hfX6��L�����<�U&s�~�)CPoe�+�[3g�iSl�Å^����T�9��0�� ��m�B��4��lb)�����rDT���M���ͥ϶zs$���k�=�?��9O�&<q+a����/u�}�R6�	��VF��Ԇ�Vê���a��'.�=�ץ�.�������Ƚ�4�UR�m;8R��$@/?�Æ��h���QS{wu'vz�]e��}ά���#}q8�;^r�b0��&k�g�^���C�����n�EE?k�N����2l/��K�P�vl�����*�?c�+��^�s�Ӟ�����d���P�M��vM������dy+e��ٷVg�%��H�7_,MȜD��j��֣i1j<�' �E|�\�e�L�q;c3�0a��@�Sx��F�%��݈cL�tn3KD�\��ڱ{���|�k\�ͩ�m��Na�4�u~�L@m4�YP.k��/Y4e��3L���eq���ҽ�#0z9�=^~���-x��J�/F�g�3�ng��p�{�e����ҏ[G�W%k3QK����%�$��_t<����8�d��^(y�=�it��O
U����#R���������6��=m2�Z�h��VM�$7�&�-?�/K�R��l�4�&���ʈ'�j���pg/ñf2G�:?��k 4 b>�^� �&����,%��!
X,NN�N�&����Q*�>�u.2��h��e�(�y��Y��t��bLʛ��x���M��؂�Q)�7���� �x+^�X���Y@K}d����e�{}H�K��]�c���ͷe8A��S��<������f�Z���-�V_N��O.)Q�@�&谻�B���ݦ�{���Ȟ�I�a�Q'�	�*���Kb7-�;Z<g�pA�^Cv�L�}P�+�B�ʭȷ-�d𑑆0�.�-F�����m�p�A�BZ���!���!�����Ei YN%|���~��'K�L�XC����reDN,�. Z�S)�ܲ�ô�g5okw/a&];�J�X�(K��o̧�=MJ���j���`��<�v����[�/�o'�Fz��R`羺���H�<tXY�}� AD�T_�������?ϩ5��HJc�zNc�]�%M|�d�b���\m��8r���T}uH�c�-!���wp, a���x�5	�R�g���	��"�&A�����:߰��	M����Y��ʷ���q�?���>N58��M���}b�'rH���M�H}	&�(`��P�Oz��3�]��]��8��7U���x6�$ϩ"�3��z�]"D�a1���9Y�O����`���mep������l���r��x�`�{��PŰi�׾R�Զ�5F�T]"X��.k+��T����<���>5M�*�Q5���	6�[)�� c��qP�p�Q3S�͆��Jɒ#}8��}�H�J���n4��V�)	[ւ$]t�W	���c�	C�u�V�A!� ���-_n���J�"�L�`���W9,�m��"�}��p#��lC#��f:��Ƅks�������5߉�R	$����hSYX�\,���3O�[&W����E���'���.n��Q�s�Į=��J��pX>��r'��2�?`-Ѓ�BʁI���Yh^.�>�)�G�L��I�W��(�SA�b 7R<�v4�*�����^���� .6��tr[�$,`L(�^�`���嶂5�w�r8�	ɑ	�@�]L₥[D�x�S×<RР���KV���Um--� w�E>�6�Y���'������]�d��2g�H��F>q�uVStLS�w+Z��3o�!��<�m����;�?���7NKZ(�4����(��O \L'OT�g�k�eU��ک�e��T�>��B�r�!W�pթ���F�O|6���E՛|K7�<�[~�x�zf@�2�ƸQ���*U&)������Q�"�$�cQ8+��Xe��l���;-�5%a�`0���LPQ�����\Y ���C�3�Ы�n(�f��B�|
��Ϝ#>$�E��S�Ji��VbҺ��9̠�c�S�,*�q�'c���a�m.L��������/2gv��AJ�4t}S���p\G5�{r�E�_�q�%\٘��]3�ьS��j�:�	y+�R���5��HoUh���;*���%��+^���%�N_q�Ӻe�R�����*�3�,�zj;H, �$�Xܵ R��m/�B=�Y�P��<.�F���4��B��¤TW5������i�E���e��e	r���?�������l�����LtP�`�m�g-&/�7�eW�S��	|�޽����|�8嚎�隳��c��wβq�!������Sse��،�Y�1 �ڒA��I/"��af���M�Ӡ�n�	 �b���1"�K,lʁ�;��]�����2�>���3eY��@�S��3U��<�m ����@��%� D�R��q+E��}|����yG"x�(?��Tg���� ����`��"d��l��U�G��j�	Zz��l��<���������Xaއ���񉮶YYC�{%�*hl��N���$�X��� n�wr���"'$܊:{D�3��`c�y3ܞPCĵ�AE=
��&Y�"S�?<ţ��!��V|"�*c����';�p���8_����a�_�ck���[�;����#�3�m�{�ax���S#��\o�G���R�R��� �����q��T
�'��B��蛽� C[�X�jA(�~)S
��Z��Z;v������J�{���EO~=��!��--��1�`(z�:�Ep�����K����@@�tA7p:[��_��.�D��_w�Y��)9{�}cֶ\���Vx�0{���J�ub�#��iW�;��(\�k��]K}�R�H�~��� m��?:�%Tj��mj��Kh,�j�{^�Gmr�z5�=j�O�]Q�K�����-"���'����Q�݁.(}R�}
���*���'<���P�n(S���8Dk���Z������eDb�+����k��"�����\��wR8����H��(�%�p`��[]��9y�LS7��CP��al���I�����7�;��R������s8E�+�y���,�HOq}Ur�7��P���w�ҽg�8�Ac���Ԟ4>�r�USɂ3X�C�aU��)(��c�Ō٢S�p2��]����.������E���t3]P���4\��D۱cgd�8H��?���Ȭp���I�	o�,�o�3�*��o�r�%��:�w�m�9lX���*-9$靦@�7�x��b1sN��.,&'ol���� �ƒ�J��=�Û}�H2;�^�PRv>�AOy�G	0TޘR�A��͝?�tt҈x�QR"[�1(I'C��������"^�Ʋ�WcM]G�bl<HA�C�g����&gF Ⱥ��H5l9����SY嫌�g�ˑ{���TSغ3�z�������gVj����#���8Tt��$����Y��fP-3�Þ}Y��|�� �W�#�[]�x�s�Le����0,��e<FzIe|Hio
循P?�xg]�_��&�j�>c�����N��U�B������qC���>H@;��'�O�q�c=@Wmӿ:�����2��g	Z�h�iPW�z26YhEU`�^Jà.�u�86<����|��P���k��̡\LMl��;x�S �<�}g�߄:M?�\<홛� m
8���C*x��%�GN�<�~�pH$�ӹ���:뼉G�Wu|R�<�l3mSS?�H�ڗ�;R���Q��֭�����Pp:x0?Z��t������'
�,n>�9�ZQ%"��Z��k�B�7k7��<r>���Wp��k(c�Xq4X��gP�H���#$�{i�v�9�H�b����:��|��.����v}�2��zgDg���,�E�����EI� ��	oGR\���E�eG�;�	V�?���!'��l��-���$��Y���}�#P�L�J�Wt����Zy��ַd��\c.�@M�z$g�i&�UB�;o���U6��ǳAFs�1���,���97�Fq
3˧4x����k��N���_m�nT@i���M��@@k:
Z^@XP�&�����V�=$�A�	��`^h��j��+��8���n�$�P(��\�{�ir�>��N=;ո�8�����e4����)���֝Iaj=�W�\�R� �`�"+p��^�ܣJ�iA2*ج��Fĵ G���2N�a3[�¼�Ğ���4ҥmcKu8^)E1��Z{��lV+X�5m%�9J��-6��/ԵV�L_�k:X@|8�Ґa����)���{�7��a��_nJ�U�'�l�?��.^�B�~���,暊��`rN�?6#됋_��4S�S4�!O�R����5���)�[5$��Yl&�(��v�7ߖOm�.%�]�|�On< l���q�OFz�� JE�|[����kYނ�ba������H��W�`
Ҍi�t��pi{Lh�*��n���|y��0�qYb���͐}xcX�����wQ9+U?�uex��[!��R�O컴�G�&G��:e���g}�an��6r<��=��,���?�#P{\�W�lk <���X�\��B�ݒ&�$g�q(i�= Us�xp��&�s�I�������*b�ȭ���B?<�ᵡ�Z;�G�XL[
As���#{�����1�f��n$�����9x3����\`4�L�O�_��!zN帊~B钍:��uq@̧���4E{����/��@z1I�s�C����ۈ\�䮯�����Ю�b��
gKy���k4\�l��{tC(�{MW�ԡ�J�z��jNZ<�U��oX��������,�X��*�3�J0�(V�C0�A�U��$�X� о�p6��eƟ>^��,C��놊�bߒ�a���䅛LX��y����f7f�o�N�+vq��Y�-��?��!�Y[,I9�(O8fJ�zh=:��O����j�9�^��V"�L�5��'uk��%k~��0���9�"W|����n�CIp���u�ɘO��7%6��M���"1I	fny���nO����0{��E\��k��
4�.KW/���i��KWe�{��B�(b:�������<���Ƅ�����o��G����:�Vm�f.=�Araնɼr���FYjI#E�������md�U/�[K]�ô�6��z�KZT��W�j���2fY49���!3�v�V�L	�R�G]���2%��I���q7CD�:���x=n9#K.A��u6���%�	_R'
��*z��3�bUbVa��Js$	c�����H �MRm��F���k�:��\�F��#l��Z78�`�w=�f��}ݐ����tX�c��(�)�qV@��J���`���ݣ�����[^R�2B&�L�N�&�C�0�����Ҿ$Ω�6LI���Br�N�L���V%���fVJ��4�Ȝȍ�{��,B��h �^̎���ӕx��'Ѽ�h�����h�m>:��k��ύ�V��<9���r8Y��Eac;�\���z�"���2��u-�$yt��m4)����6�0����li-� �|����9՗��v�r�ry�n,]<��e���U�+�b���;�^Vm͆���������U���p�7h�i�;�:늭�9�y6:ڧr���5`f�C�l�0�q�Dn��� ɊK^�2x���5��uۑ�]�Xs��8�K�O�]�";��.�"��Ɨ����&��T=g���蠈v,Ԕ����d�|+�av�eDH��&XwtZ���W�3<)_j�eM��K	�A��������?�D6&�+Q_>�ʫ�5�F�(���DA��rehnd���]�Cm�<S�$��1E�1�4�W7�l���[eD��h�쳷�k�x=rL(�`~�ʪ;yj�J���c\�FA�#%\��1�t��}�����wK)^ny]Ɔ�O�װf�n�*D�1c�2������>��z��%��سD,�d.��Ǒ�$'��I_�J�������v�SG9;AMU}��t��"1���յ�����#�9\��W������9E���h�Q�ۻÔ���T��V(O�J��!�)k�RP�������$�|��\��e��ѼZ���ߟ�-���K$�<��i`�?���*}[\^W?���3]@}���x�]��s��gbf,�لȫ��[�#����p#��@wI.��M��=X7�2@�u�OMۅ�Z��X3L˵�/���i�%�	�̮u-�{��Ӻ;Y%C�?����_�vNs�e��BI)Ò�]�)���%��k���n��[H�n��8��ތ�o\0�IRn4N�d*2��i%���q�ݷ�x�w
2�aMU�}��;�h��Z�$�v-�o{�B��ٚ;�a�OB;�Rp���A}�*���Z�3�� M�ȉ$}���N�8���Y*�n�^�5�X
48�ٝ���M��=
����֚��i�� ���+�5dQYsd���?&;V���W�R���t��a���س�� �1��Sfy�\l�<8�u"�=K��d�=񭑂�/`�h��ı�W�v/���?L���%c:Z�k����p�ԹX�ޞU�僳��"\t,��{�a�P�!��1�Ԝ�<"�L��+^��&�D)�@���īߦ
��*2`�o���L_N�|2�Ʋ��DaOÄ4�ݼ�Z���z�;n����"}�[�T�͑��ؔ�r��袔C��U��ފ䷷�pv/�izb��y��_��}���R��M�6�'�t��$I�Ec,\\?Ǔ����~�����@��.(M��!_�˘�s�5˃�pp��E�D���ǧ����n�3�	�y���YH	�/��jG=�AAv��[���5;D@��|g�,<̄�z�x �b��?)��~u����?&�YvmV1�/v:��,a��)Cn��y�dōXP��+� t��&����v�L�+� �,��<.�����-)&�~�s��5{��X��=GJ|a8${/���}��
h���ǃ�`�%�b1Noj�t������$Gdxmy�'���ns��7���/�#�B+&J�Q=1�ڨ�QH��6�@Nn�ə��-7���&���;�v�j���~*:�+v3w��ɕ��0/��lE,8R���/�*���+"~|���Zv��tε;��r;%�3��Y��9�7��on��>-ĥWנ�R�,�K�nM�#�²�l��2/�JK���"	�B7�8}[�aưO�q7�j5�;&̛<��#��f��g�)۰f^9e���覎d��׈���'�м�>�=_)���8���Ğ���^7P|����rv,Mj��W ���g��Qr���<1��A�T�\᥾r��f�zSRs}��:fC�P}�L��E;b/	C>����Na7�!����pH�t\��r�{��c�`�z:':��Wp���g�h{�ϙ��=S4/!\�y -��x���3 Vm��SX��z�ԨH����Z�ר�&�"��3]����[p��~�#}+>�>��䜦'�U6�㖢+�`�zu�5��ߝr�.(*�J2|dm}Q�-�H�it�臆�n<��*�˾U{�����(�O��/Ʉ�oF�V���w��*�x���Pՠ�y����:S(�H���:����:�}u"�L�FN�#�:����
M�ǜ��|��[�ơ��d�bŉԭ4٬�;�x#����Rm=�� ���{��]x���a�$�97�&ԥ��L��a������-�E��3������m{�J��r_t��&'��t�$ͭU��W�g��zh9�I�?�����S^E�ʵ�`9��9��"\���P�?�{I����F�4t>v��m:U�Le��+A�m�v����Wb7j����:1����IC�>H�6% ��U��+���vGƉ<>.Fأ�6Y�������D.�g��W��PV�y���]CL<�*R�;���}T�V�n�� ,]?�8�Ԣ9r��Z�bG���1~}�g� �q�o:#s�+C���D�\������e"@��k9�!�q�s��b-(v	��c;3(٪�3��¥�/ �9&�F�Ӽ�����<yx��v&ts��6�w�۸�O���z�E'RCL�\�d�ʋN^F���k��b��m~f3���ň����+�s��D��]�j#0׀]�|@K&<��;ؘ/�[���(į�rm}cqO[���F��S?�K�Ɲxv�l�T^�!�b���	����������X2�1(oa)�"�JsU7>�
�9��f_ihi�]=Eu���'��uR���q�~2yS㥲���b�ȠM��W���r�Ҩڙ"H��.�B��8��l�7�4#����Ѿ�F�31L�� �c��ѩ0k�y��9�(��B���U_;���qS��9C���������� ���n�ҽ,�,��L��6`�����Ȟ�b	�3��ZKJ=V��!�v��J�j�+φ�zg��|Db�V�5�O�'v�1ѿf� �{��<
w��\�sVS��Ag�mb���<'�Y�}�E6-m�l�y�5K�7�ڴ�fۚa���%\}��$z���'
bZ����1��{�v���1'��$;��T@�t�����Y��{`8r�B�V$I[��	�d�����&&ᥘ�.l����(,�)�3������E��2�>[�j��`�?��/���ǂK��Y�[+�-�>c �#Foc;�x��45]��9���zk����+g�)������R?*�{����?>DǨ�lYL_[�I<���o����s�
\�-��k��w�y��Nʎ/�m��Jb���`?��!���}��Knfng>����Ƕ�A�a��:�@8'��Jj��JQ��i�+�O<�T\�zaM6MH�罩c|�P�/���r��1�YU�Y��3�NWy�NV�.ƭoؑqԕ��DG�a���x�\�w���&1��e�aHK"oZ6G&@��C:��;��P!v�$��e�F�/�g#&=S�g�r���Ǡ���]� �eѹU���H{p 
���N�Kʃ�� J<L5e�([)����7	�SPx?�:!�)*R�r�0��{�Ϗ���}�Qh|�B��-((0�~5�/qN�x4*z�gd�����ʮO�?^���W}P���1�=?֦����T�
5@F�y칙�z����0��5Oc�5YS?|%y�oO��$#��_π�w�W,`�,b�G3��N�xMj��"�;9ګy�.�T�"��)4+'�HdmG�`
��b�5�^���<�t�����k[�s��=�����9������w¤�i ��uy�,��#���	���^V��7è^IK��oF ��[�}��nn �kr���F���u��zH�7�ӭ|&gvS4L�a���n���9�hS:�xI��?^g	�_4CG� �c��4Q�����ON�>��#S8+b��sSzM|	���[W �^�U�I6M
lwP�C�rF��Os�	;�
�XhYQh${���Sy)�{��Rbo��YvU�Yp	ۗ��n|*82���G�J�g>r�_�*��i�E$$�0�ttìYZXҋ�OV%kD3r[i^m�;�t};����z��U����[y�{�������lpO��aU���^��`W�68�~^�s2?xw6��d�8z���@d�!��N\[gx�X��>��9g�٧���U��bʈ��z�Z�-�pe�ja�t���a�+T[���� �c�rM�*�ۦj��,l�������vH�twͭOl	7�awW��o�ǔ��i��u�萺�C ��~��Ֆz����Q�cN�,���C��F9��I� ��5^Vy4��K���D� �~;���^������)#�<��~{�Xx�p� �
��D��Y=�!�m΢A0�hc�u0oˎ����u��5l,���8�b�Fʂ�H���!����Z������T�R�}�?7�M��?A�aL]�K�Z�*�3�,����{����pK@��z/�XPV���ۋ��<aա]�ɋ\W<̍Vh�<EY�j �U�է�71:����Il��Bx�Ͷ]�=A�>յt�v�|� �|Gq����Z dd��C�����c}S���(ip�i�CT5[1"�F)�9���l������}�Շ@��X,جc�ZPP�/�9f����Bs©��Fv;�f���z�,_�p��LI�m��k�,c.��K��YV̳\�Bղ�Ռ ����������f�]}G��(�$!Kս3l����#Ui�P胉N��h���c�����R+���;��F}����h���Y#Dx���-p��Ld����$"��-ݩykt�v���[��* �oGP�.в����`LDč����B�u�wc��p[S$I��w�@�ś�����W\��b�����Ix<���Ú�Y7�`;��5��V^��X�g�Űc<��i,e��7���C�!�>7u]��d��%LE�]Y�7�Ů�|������u���g�Y�+�����㙖�m�Yn@�i�f�*�gV��o�p�'aIk/T�z�Zo �@D-E�>�^�[ �ת��0I��Է� ��+U�7� *�]+:3IF��I���3	E��������?�ե�ozv�):,:JT�e�1��jzt8��t����1�u�VY���+�r�p�Yܝ	��ԸiX=i�g]l֠g6.����Y���R�vB��@l]������_�"}V$l��x��d��ps��V1��c�X�?\�k�ҢT6L. �<��i�v��o�.��xb"f]l)� ,����m�&�*��*_�$,��m8�G�` 72I���֩�|(�!��Ia5����i���M���O)�%K�"�V��	cd���o3cw�mx�m�pn�IhC�֜��RkC�%݋N�!�7w��:T$(�r�֫�.S��o%�����_C��x#��E&�]�qgr�K@-�&�[�k��.�0Xg,�ꈏ�	_����=PK��;5���ǽI�����k��L��x8iG��yF���V�4��X:c��L4��)��,�*2����"���-��brX�cg��Ñ#�D[*��(M�3�H�_�Ε�4�fnh�3VחN�,�ں���}�Q�Ʉv�`��qâ!�m^a5��&��O>i�n�ӌEŘ�����{��"مe�)	���k���i���֤�e��� �f���w��q<5B��;A�9ڇj=$ܞc��>!���=�&7��w����P�g5�Z<���~v��Έ�uҕ�7RzFTШ���{��p-��Q�4�y�WH��s�Z�aBt�����s�;:�k=� ��=I���T���~�+�^���M�-�s`I�s��yyvqL?�������Q�GgA=f-�Z_}���Ԏ�:�p�>�āO�=Ѧ�qj�4vO=yAc�igY P��+!����ԯ��0	"���9�+�Q���K��7Hj�a�^#I܉�OC]B�z0\Kr\�[$Pt٢g�!�G�5G����
*�˳�|d�#�%I�x�����ϓ >W�7O$���9�T�[1\�,�-�J�MnV��c�׉���=�
�����믌���j��[�N���������=5�,r���mf��������3�=�y-9>R��W6$�<�%؞-����vI��m����퐁Ū������6hحo��L�A�b��f��������>�F>��<�UH�����r���"�!�o?�����*G��Z;) ���E�ɡ��NgX�5y[EӒ��`�śP.���e���RK�K�,p�靥��:��x�3�e�=�	�;f!��[����k�5ǆ���o�D�^9�����ߥ�%�N�{$g�-�hĚ���.��벒�9F���\��V	���5ʩ��}�a\2�-Y�x�>�+8�O��q�g��<k��D�*�y�C�>��B�?����C�a�������p���#�	ӵ�!P�j@�O&�lp��;`�	���lK�ϣ��S�a�]4�
g$78���{������u��*aa�fz =g�"��8a��R2�C�{q�C�ǲ]�����e�G>� :����xzth�q�[>gtT#���t;juP2��hj^����n2f�s�6~��
Б+U�U��\�����*Āok\GQQ�k���B�����"Cj2'��lG�0'l�P��7Z�
�ǝ4��u���e�n������)TjK��,��tmN�3%%C�R��{�S��S8Ơ?�&�e2��٣�DJ�v�x¶Ԩȯ8��*��v���X�KC�:E�J�N�8�T(�^ks�CdUQVBܫ��ŧ<�F]�)�Y��y��&%\��=��B;��XHΫ��Qe��^���~䪖�q*&������bRȈF�{
~��z�5 �4_\�`˗Y ��^ێ�M%��P/㖢�0Z�Q�j�֦i��n�ۚ�><v~�
�M��_�xsi����( j��qMF��v1�}�9ڲ%By��T	I�*�7)��8�j�ۦ!�0$��̂���n�J��e�lq�K#ރU��@�V���[�"JD�� [��ʻP��y�+�n��+-�E�+��˃NZ�h�M�4��������\�Ս���즭~)a:,x��! �q^Dߊ,�Y�B:�g�y����w#��
�"z\�V�HM�H�E���0$���|��h�71���RxD�df��Yn�&�̑Ѣ��i����b������˦����;�L��ơ[Yr%P��X�s���o��C݋!��LX2+3�0�����2u�f{c��=ݤ��:>�z�n;i(J�Q�r�fX$6���˅I�a����A���{�X��G
?Nū`F,����{a0�T(�F{dN����=8J�ar�ν���q�8������6C�i�w`��
�$5BFf��ܼ�<�R�����(M#	\�8�Ȣ�$^�+=���M�Z�*�Nx� �o�Nc������	����k�Q�X���TZ gz� DLJ�@�v�&F�is��ID��Ty�G�b){��#��|
��uT#�s�w;��/'N��(�G=
�c�u�۹Ӻ��Λ�v��v���~��w�6��BkR;�,2���;�Uolzh-\�h���h��	������)"?Y�(e,3=o�ǌzkKeg�S���JE@��ԯ<6M
��q�������0��,�'��b"��1)��U�y�6�c�D��)� 6b�]�T�?Ul��+�����D����]�d���1ף朋�N�*�W�.��qi�Xe��1�%o�|�bt>ռQf1	��4�qm���A��$�툳G=~�AP]۷	���Z��Nf�����%�v�o���B��V�Н]�4����D�J*.a_*j�AbB���/Ѭ�@�?��o-��p��-E�,��	0�Ơ�R��<��'p�&7�v/�h�Tv��J�$6*�8��3(=F��C��g�4��e!E

�kM],�{�z��{=J���R�����C3�lo�����Bn��$���$��\XQ^0���a�t!h�G9�"�+[kj]���V�� Xc�9�_�tJ��ӭ�p�а�j��Q���0���ā�aR���Hm���S'�mU�<�kK��%ԕ�T��'�X�kQ!�;S�>MWf~W���Yz'*��C���t����Û�e�N)äk�yҼ-R�u�ii�׋�+k|�V`փ'=R��k���ب$$F�~;G��z=(��]F�l�_1��zGnA9�����K�rڐȂ���͛�G�q�r9�6�}�k�����Ħ1��MԨ`Մ�z���5���k���ܠh,.�O�k�Ψ�����744U�Ӭ[�S��r*�|�o�_���4[�4�������Q�ZW�#Sm��9K1�+�D��u��r�p�o:�������UTY`�vl�����<Hԏq-K*��^�܄%�Z��C��`dD��!([�9�˦��Kukړ�W=�*L��bR$/Rg*����coYĸi��S��B��Lk:��ݹ�5~	a�l=h]dmj\4Z�Jmsk9��}9g��,�~x���giv�D=Ĩ�7}g��6���ۇ=�(ްP0���������j4u�y���-�N�]rw�+�����>�d�,�i��Ю�T�'N��r��ˌ<J��=U�9�r����B���EGÌ��+�߀Q�qnxkD+�b�[b8r=��Xzo˥�����]4��3:�^�~!}t\DPH�6$<�!/ ���њ����V���@r
�ap��$ K��%X$���!�Lx܅]D��Q���@���K�457vH��S��Ve?��?�=�T��T�Ҩ Q��H(`b�ti.�X*�m+I��F�k}���@�^������J%��4�csn6]Zɞ'�ߧ_#��<����9��'�!�zu+�O�vs�N4b5�ыƝ������.r~Na��)���R�ԡF:(����ZZR5-q�۲���7yMht��<��#6�}��s6=T:�o�_��o�7�� L�ٙ;<��wv�+��#wTU1��6IC�"D�YIC�N.4KgN�$��;���%���]e<�Jn�=�Q��'ԎC�Eq8ł��	-J�e�Y�I�ږ��M�#�;�zk��&��fC>�V3�Y���}�ϱp_r�Xn|�4Ǖ�<�������5&���dV^/m3����-Ry~�dW+ks�����l�Ǽ`Q�)�֝���Р%v�mW=c��C<t_/Bd1��w\�P1���j�8��@���n<�Ǻ�93&| �W���o|�Y�C
�^�~����Z�����5`�q��ʇ�_���z�.�}�o�P��P����j|uD!��,��0�{��#B�STԂ�R1o��I�G�ə�x�dܩ�
w��IM`[۸T`��r�Ш�^�뎬:T�=�v�܍a!�(�����5Y���XY�`n��U��N�@��P���ãp��vI�N�R�&u{�TpiĐ��Ņw��d��[U�|�@�u�vl��/��Cnf�����ˈhkz�_��ai�cХ���4r��@o1��ߟ��I����'�	��?#���L�f���~ǃE[��!6���!ڒ�<{d���@���?�b�9�op�/[M({�'����5�b�Q���ׇn���:ԯ Vq7��X�y66d�Zq�4�U6̜�<B&-���8Kl�5E!e�m#�m����1���d+L2˚FMu����vL�%%�����+���E���K?y�	��<V��뭒<#G�&�57�鮫�Y*+�n��:Yb:fo�	�a�~��x�@u��54�o�іF�T�n����u�uQ�G]4��	ג�Ͷ�%�>mih�� >?�?�sX6��������/���p¨���yo�f��a���: ��f�&�i��G��6�'u:�/�jEa��}�S##��$:H��;y�Q��K%Oj���W�c�h�ǰhG�K1쇚��R�a8ok_,Yu#��U\T��c��� ���С�hx�
=e鴰w~J��+�V�S���w��B�(1ƣ_bY¥�)��7���;���D0����e԰�����j�UĽ��Ω��?��f�(��6$�DFc�$��5��k�`�X�	Suu텓�w�W_Zz�_����m�ư�����{�' �h2�����Q6��3�r���1[���a'+�Qݗg�".f9�gZʨi�2��<< �����Y M�������Q��~%U�fZV�|�>��G���S�`��sE�E �Ͽ�����A��ȟ���2S�yqbɾz^S� XRun�n����U�J?Q��x���/�Z�a�Ș,贤ފ'w!�(���	�x��z�m��|�{���ѣLv�/���G4���m���h�
2Bu��6�ݸ:���{j������VG�	�Jۈ���X!�:��t�~���V,5JA�E�J³�B�Vu�>u�jjA������`e��+�	�~��9�t�o�ՕNzީ�ܧ�"���VV�jpDL4:���eL$g��<#���V��=�YS��RCL��H�L�j<�@�߃BA��
��Wv��R
��Ͱ�!\wh�Į=��ct]����sLI}x�|H\���~&(�����ܖv���W�Z��w!��RnhM]�Lޡ�F���@t�6|��n����,�9Gu����
5������-�j�%����>����c�6t�@��$�2�|�R�����\�~x���"�����6�))+�[��3!t)��ÿm����!�/��S��3OB�WE;�j?��b��u��w��iȊ����X��4�4^R6 n��L�X;w�	�v�)��Av�]��X�C�͇�9�SG�ߤ���K�ӗ:T��p��Օr���=%]V8C[��5N��u+�7��v�6��S��[c}�b<O�8��(�#�g>����	$B&��	����Д�s4g��<�n�F�B������Őr��§����y���5��@b�T�_���s�*B��=�\���[`j�I2.Lø����7����TvS� �#��@t�Ѹ��W���`G�w]l����U����X!�Oe;��͘�'k.l����5\����%Sg��D�2�F����}���*�N��o,\�?�� (Щ;���A4X�����HJNS[=��oёlR`T���A�PFv�ʫ��C��|VS@<
�$��W�{�݀v� �=«�����ִ�5HMǿ�|����&�T�\�l~Z�{���lyN��O��t�_<n����f�jpW��@��?�[|Q�'R0��!�D��Ɣ�w�9�D�|�+v�&i}l��A���^�"�܊'���,O��'��?����BT<�c�ľ�#r_�[��c���������	�%l��{@yϘ�e㧣V�81^�u֠Yptv�T?�f0O����}��_�
3Yv5�1VNH�&Zz�j㌨ԵIT?T#&gL�u0\��h��w낲���a�T4��sմi��*��|ՏG&����3 �@�E��(�Q�旅�aqO�yCa�gm�m� |�M�����N@ψ�����S�9�6L>c*q �F���5�sО2,|��2��,��5�SlN"X�y�fM_�.X��w�X�'��h⊺&9�wUl����^���h�x�i�z�����a'�˄{�	ȭ��]*Dy����Z~ɯ?U�� ��/�&I�r��a?ZK��#�|�h�Xޑ�E�A��(�?��̓4���V�`6�Rط��IM�xv���
�,���F�:��v;c�]�M�	H8e9a_���&s<eAȯ�K��s���ڕ�P;����N&~:���Qn]p?,��m�"bm�4=���|u,*�(qǤ��M]��˳B[���#t�n>$\q2{xبygk#sl\���\s���Q��HN̽,�-�����"b�H�����0a��yk���m6F?�(�9�w����{��Y� �3�<6:��;dr�w��}-���wOA���҂t����ʱ��a�hn���	.����q�����TP�*A3���\,�����ӥ�/���\�;�4�6�C�z���\ɵ�!<����.ҍJڰU�^y��nE�:%+�K��u�o�7�sU-Vqڲ%��ۼ#on�	����a��ِ�4�j�s��-��)ZB�x`�M�AW
`Eެuy���V�*f��8�.YH���i���,jF_y0��r��� � ��0�Y[�`�9����ԐU���@����%�&�-��L��nE�3(`�G�,�n�!���fNg`L���5T�߻!��u��ދ�?g˔�
,�鱼;rU�	(�������c��'Ҋ!@�Rs^��W%.<Z���z�ƀ�gO�������C���c5����8]^qP��9������Q6z���r0�-�Ƈ�i�R���ǈ��P����OW�e��.�R1����ջJi2Ȣ��^��F(���̔mHML�,ڻ�@��Z,�.���h
da�0h�y�(�WФ��n�ɀG4ɠ����z#��|�,H�ڈ����'
pVmYV�z��$ X�c�&6WB����S�ٟwV��5R���-��9��H�y:��ǣ���ط�׬�?0ƴ�Z�E�*qu��6�2:9ߖ�Tq�y��,g$@�#ŵxo�7�RM�]�M�e�9|,��h�3lE61���;K�/漆����HK�"L3�X]���d��g�iXGV>C� rǼ�_�6�x|נO#<�l�[����4Rv��b}+���;�zyo�V�DאH��9�Γ��9���#�y�b��u��%3`TnȨP9o;���Gc��p�"
���c�fĜa#�Z���M9w�}�̨�p�i.]�̍}�����-�oĝ+��I]7+�SQڳ��� �<���i���`tS�#��T�����bH
�^MH�Ȉ�K��$�L�� ���3��J*p���QlX�<|&l�C��b>���03����%����)W��H�|D�tj&��1;Ȋq����+�L]y��bZ� m6��Z�	�R�(9��U@=�Py��Վ�vn�>���U.G�U쳺�NAF��t<4���d�O�u׺d]�Gkr�~miXY:>@�g���*��fwq/�*U���D}�s�e-�&�5���$$ː���>�x�ւ�'E�����$�.��|mNPA����*Dߩ�8M6~[���w�SD��x��]9�c� � �C'�x��똠��;V����h�q��+:J�4%����޻!���_v�e�&͈�*k��!{��-��棎��gC0Kn�o]�{�1h]|CE�9�{����@&�gfl�n�g|�Z�N�]�%�dz�P�O͓z�-�����8CU@��$��}��u�����:k���P��3Z��p}��;0�K���9uբ,1�f��[S^ˠP6��94��K���Nv�Ѣ��M�\o2��{�"�P���&����{�E?R�'PϦ��?a�i�����_����4�W��9�vt!�k%#��H�mgl穎�`���7�W��R��d2���]}x`��ʔ�B��?q�g�Ngy��( ;ꃗ�1��:�%��2Ї�p<��Cp���ڵ�1���=Vu���:O<#A2�����M5脰�y�6����� ���E�\ł鬞�D���j�%�"{tF/,��������Y����jS%�('�'�A=n�l+
�	�5��UF��N �&�6��!&[ ]�	��Ȃ\w,g]�y|sE��.���h��b�Z�E���r�?�$�\_�m��B�s�I|�f�2u/Y�����0_e�}ԅ�G�E�n�o1"X�g?o�w�"i�_�+kH�6wc�Mߑ[� ?����s����$�2c `q��IÙ3?n�1��˝V_F�I7��c#d$s���X �Ϻpl�6@�j| ��ڕ317S�M����q��;�mh�3K
��w�n���}�L�{KϦ鈠�N�h� \p'tb�����Ha���ķ�׃��5����~���;$�{�tN�)����w����7�k0�s�jd�v�q�D�Z�yK�$D�V���M���9S���%�	D�w�@WM�/�<<���-'4n��D���Z\���i�Ǯ�,E����9�V�]����im����s -B^�v�W&�&���:�+��g��醈
ؙ$�Ӿ���4�#/ꧥ@v
����*C��`��Q��(��<��m�Ђ�=�C>�ʹ~�塷p�O!��7^��\���N��,���p�;�.�U:���!Æ�
��讨� ��Y9����e��
`U<a:�=\d�<�Ბjp"{��/��w
Qi��L������B�N���}]��K�7<�Ǡ�y��`#�Q{HľEU�+v=�%���+esUf4~��Ҫ�G�hiz'�Y_F���K�U�_��e���?,R.��;��i�u�%����noZ/I"e���矢P����SF�b}�oϡ'߼1�j��^8�p���+�vw�.�L]��o�$��o�C�,o�p�����Ah�"�}�\*H���ݚ�yޜ k�k��˲���ݖ Ӌ"a��,����V���
��F�C�[]TL9�=�d�� �4�	MC̄O��Wv~#@�;�p���x=��gf<�L���|~O������k��]��,���0^a����@�!s8(�L%ө�f��y��F�R�L���>��KE�a�Gj�ͪ��X�_N5̒W���{��e�5�S�M��L,%Ԯ3Ou���KD�<=1fǋU�8�B0F{�Nh�K���
�	��On�""��E����Bپ�X}�İt� �'�g�[ȿ��6�:s�Y��U�����'���۱jj���O�����ѽX�0<@\�!g2�d��
c���������K&%�`1�w� x��G޷��Z�a�ʽj�!���E����	2��;n�LD�X]ud�>i����ׅ4D���ĸ�J�H�o>�̑������	]i�,�@jk��f�C�ՙ�B!�&w9n���aA%�n�n�j�>C�7oO�� ���ɸ��F|P4��g�"B3��gm����EZ��jK%�7o7���]��@TW���2$���Y�^�|+x����U�HMjn�z����H�K���
i�܋k���v����_�R} ���Z��x��]��]dG��ϰ�-�ܰd�G-� y��^�ٸa	lл�<AN �Z�8���&���)ς�p���uW��@�~}&�ž�Dt��b5 !��ɸQ���P�v'�t��f��v���1U�K.�'�ڹ�*)�-����Y�@KT{T�1I&���t��U�(6X#�a��{��m-������Gc�QYH���%\6 h� ��e��ƥr�p��Q���\��𔷼
&���
a����y��� ���('�5x��sK�V80U�s]�ݲ�9(��U�%G�3�3;��t��G}\΅n��6.]�ȝ�v ҩ���^M@�F!�,�ؠ����h�=����Ћm&Q&�����j�s�����BA���n��[��x��dbDZ��>�iT���Q��e�^�@��1I|)M��h���q��l�`�qPr?d%X�Y��v9 ��yݲH$J�f�<��:{��+��>|�=�w	V��T�Iou���/!7k�_�t��L�2#�R	ۯHB�<�\�_���R �,�;<�|��-+��e��=�7r\>���D�;L;u�qTI�.��G��i'�vL�_�	��ffJ��ذ���N2�O[�z��N\��~�@U������C_�Ux{�(��֗`XU>,���gD�Y�M���F�12��*s�$9�.�a�_?�\�x�naM�y��U�"�*��A6r��]�?"N��:d�b�~����P:�z�ʍ��� �v�(�c|��կ��J��i(<ÿ�����u�sB��܇�+ l�1�!�LUa�Y�?͋��S���Nb]�Q���`Dz��}����}=��S����`g���^���v�ո�WU6�b�B|g�B��R�"૗�e����k�3"*x��%q�'T�W�"�c	Mg���uP(�%�)bF&
%�Kh	)�7>~�#J�qkQ�*�D�e>|3ɓ�����e�٤�#�>鵄��;�����������G5��l	��[�81Y�D&m-�t��P?ې8˂��1<2c��W�L\Q6�p��m	�׌����Ĭj���U�!�@%S�>�;���-N{H�E�&��B�R/�� ��^��XC�����>�5��9��y�e"�u�����Iΰ&�n6q������O��ن�Ü���f`���X'�2�h��g�:��/'���Ȝ�ݥ�moD<�w��E�t���w� P,L]A9���#�S=��Ie�	�eB����`�~�2qkfS�.{�PV�>��Jof��'0�b�r;s��l8T3�D��L&��)U?W�t9,���]��5�����)�������d)`�R^Wӓ�F�dKAݱ	NS��0
	K����-�G��L��u���m��l�X�VIj��DP�)��N+MC�����8���������KTׁ����ŵ�DYm�AI��5sWH;�֮�|	q%���@���O�n+к����>���Zu�F���Z�q�1N��Ő�k�eTѹ����������L@EB����v�����G�
�jj��R�����i�,�<��wI�@�ZNy��ʬyE�����V1��/��P��r�}�y" p*0��,��:��-��[0�s�& UL3{�m��=1뀩�`�GoJ�q%8�OH�,��=  ���b��aCU���Owa��I7!�ݠX��"Ou�-�we��y2�Ɲ�D��}�#�����U9N|)y�|4�~4����!+��C���[#�ħ�ȹ ���]g&�j�M�a��@/����$���ܐ�)����P`������mH�x��'�\`zF�Z��Mz~v���TZ��1 @T�~��p�'j�X2�(�фy�B}[�R�=��wQ[a�r��>ǔ��f%HJ�Ş�W8*��;4i���������G�KKN���$@�*[x��
H?�u�	U���q�>a�'��%Lid��qaD���xM��#/["i������j2�E;�����V�)=�4]�W�q��n��U�6�Ju/���9F�]\�MB%��D��~��4�H@o�a���7�2���x�#�uI��#B�oB��&�h�S�y���V6�N0+�W�-�<R_!0j�
�zs��6u�7� 6=c2�*,�;D�,nim;k�O�!����
��z4B��`��w���[#1� ��K�Rk�gί��Y�9��ڽ�3	�����<F]��#%���NE&"�Go6�����S��~i2/�-��d��G�!���H���qo`Z3J���)�*�!ƍ� J�������|���S����-�/������r�t�}XlX�q:㊮��b���:�����m���V����V��Ո�'Z�5`YՍ�,��z�����8v�	������cGax�ϑ�cr�
u��!��C�DLc�G8�b����RU��'�%�_�G*<�U�=��MX�@�}_~ף�kW;�_�����]��� i�j�K���\ba�~컅��XT��c���ٕ>�q�X�_2|ѝ�l�l�.^0�Ս�(��nt��@�_��:p��q	��Jj������:T�=?3�[����U{��JN���3� �mQ3T���O����ǲ�rNfKp,9�iq�Z�G��X��O4���@_=���^|F<���3�<�q���H��ێ�e<�џ�M!�`az35S(d�Xeۙ�gG0H�x95c
NXȹ΁��~(k��ķ۔���B�z�!��
��ןV������Z��y�YR`���f�Ǥ�4eYl9�_dA@�5�c��9쾐�-���a{ްE �����g�O����\��%/�nq1m�
�E���Ö6傚C�|ľ��@/��XFqh<�s?�Bp�TG����k�)��ɼ��2�=��
^����h�} NQ��Z�[���	?�����n^3%�m�H`�����̵�*�E�������CC����z/�~�ԭt���5M�FE�x�9�7�/��-�tϝ��x�m������(�>o*�����m�Y�h�|~\�>D#,�˭�Q��^h M��?�m^���w�F~F��Ly�c�.���Ƀ�9�V���&CH>졛v��#����0���%8,�����+ڦ�䰘�V�r|}�I<J�v�����m�U��)����=��&��C���1���E�X�B���'��9�}'	��D��3�%���h�d��j�j�B�-����gr����	 ��dUc���Q}��-�A&��WR_��pa�4��F�b�P<<0&!.iAa��_���:�L�,|EvGjZ�h�X�=�V��z��J�ܥ����=(mXk2\گ+�sOX�"=1#*�>rao�D ��Rv���b^4Z?t�9���	��[����1��.�ܳ�XM� �c?s=���6C�N�|�21�ʄ�iu���b4qw�mP��Yd��;?�ԃd�.��B�:_�
��_*�ȏL�E�W�t��u�K��e~���!$_�[�%�"VCr 4�Q�K6}%�C�S% �{h�ѯzť�LB陫|\��ld��E�c�R}�[S���.)@��A�."t#��A�A#�,��21��%ះta��R�.v;��<E
��S1�ܹ8ݟ�����	��sW���y�juج���<,����7�Քth�����kt=!������������5o��+f|�å'.ew���̕./,���w���k�z��	:wU븻*n!�G9G��<?S�>�p�^�u��m&H3��Y�1�8��󦮕�B�"Đ�Bs� ��G��z8���Gd=��a%kP(�Y�ʱI~e/D��|�����i|Yb�*)��â�Y2	����0��{F��q���2�����@!�mJ	�3�:zڅn�t2 ^d�y.�rqG�ے(�I!aK�,s<�E8�efrA��F��� ��{�\��R�G�[)+q1c
�D��e���n�~Gi�n�����pێgp��u]�L�;�EiRe���|I�f�$��h!�f�挺L��H���,��Km?l�I��"g`�،��|��P5�{4?�=�yg��X"!S���e#d�?�YĪ�������T����͝Q��Z!��%We��-���O]��!k�h�v҂����3Z�)kZ����W�#�*0�U����>�-D;�-�:�tC����4�.)����V��5��쉐�E-��S�i�"�.��D8��Z�K��b7u�q�;.,,�;0�SΆ��I�*��D.�T���|L��ԣ1��lV��t���^�"���x�~84!�PB:�����.�K�����!�$u�"���x��[�����F��#5�?�=K���ji����X�a�ģ��,���M��O�����s�'��T),6�U�.�'��ۍ�3m� -����b���Oq��?��-��F3}�L,��.B��`M�)Y-MV�?t�&�'� �4��*C%���sw�^�g��FР�m�j.��������6TU��(���_��g�ɱrlb���o�'��=/|p׻zI}m����\7��D0v�U�(93�$� q���0	Рd��DKV[��B�\3E�,.�*����d�bjs�����k����B��c����e�~̼�Tc�!��b�>�%�	;�0���N�fD>sg1.��9Ddɯ��Te��:M�#ڶ#��ibcX� Œ�:Z�/pٳ��b�`Ӣ�i�TG?O�P�nk�Y��M�K��b��9;����QDy8��g�m>�Q0���Ou��"��RR`!���+5Qw�;'F�Ҧ���X2֩���[�(0N���At�(��Hv�Y.��,N5��lrx��K�K��l0���	�i��*"�Td*<���A�aF�����Uy%��xNQ@A�`S��*@-�k)p5bM�G=y��N7;��(~��i-�Ӈ�Dm3�#X���'l�{;L�ɐ5��G����F�/�֏���@J�)�<=���af/�-�_>���������i�i�U8��+�� Ti@$[��?"+
�v�5��>�6�e����`	Ͳ"A��/�W3�(��6i�S�׻9���i��G-17�1D��p�aH6&	#1���}e��y��ng0Z� �H�����Mo�������3�Z�A�U�09���G� 9�g�Z��*H<���af�v z6b�ŮAkRF�5�@.C����nر)O�6sD�Sd����d~n�g̜,��q���0� Ź8��eJ6��9�Ҧ�*��N�`���BD�L�ӯQd��+��7��֭��&H�N��'�3C-K��VN�G/GVE.ޱ�*I2ֆ��i�V���Y�Ex��(����k&;+����3���j�/� o���K>6��B=�d��(�?P@3�5L'��,�n�Zȧ�b)��zzx�o^;	��'>�>��]��r��L�H��+���j��O'��aaC�]uʨ�A��W��6�zJJt�%_h� sq�V����/���l��|8V�0#=�P,����M-�}��V��a^)�q�0�K�>�j$�xA����𯒉�?U�f6�%�< ��Lޛ��R�[���X;�l�.Ù��O��,ꀹ?�8�����d�
����S���f 9v��t&I�,�
A_�i2��i�W�=��zq�! ����AӖ���eQJ]��gSm�C��/��HF��x�~ns����NE�3� �Bo�<ve��b_�������X4�j��^�պĲO�2ZΗį�qM�R��
�`]��D��ڼ�*�c�Y��P��Ɋ�/;H(���M��1��A�����c98�@�V�u_��f3o9'r7�%�ºv��K�އ&�>t�ZHɧ-���x�6=ғ
�k��]}�w]����J%?t�y벋� �T�'+Qű���3o*H�a�7���}-T� �d�!P̷�oSU1��nX�3�����S�h~���%^��"'�:%��j�M�Y}z��S��7š�� ��%?V���w��OU�H�.�^���c�v�Q�"�oo^l��ȧ�cDѿv�ANk��q��&�ցbHkp�ǽ�i���4�R��V]���3�b��$?o=�P�JSTJ�*�^Si��c���p[(Q�e0�yt�Y}>\\;�V�<����D��r����:*��?�-�V_(�]��MD�tf�9�_��csX[x34��� ��8�.*��+�GIڦ���Xg���G��(hǣ����g�f[s�ِ>1�^�*r�؅!��╡U����G����o�J�f��i"�,�MZ]�;ۘ)����a�H�IA~���1Z��� ��=TvS�����0����*57.@5ab�~��6(f����襙���%��2��Um�����EiSlǍ6���e�òÕ�b��)�j�3:so�Ø��SJj� s[���0���ρ�)dU����cEn�Q���"��#��tK�S4��M��o�N�6m��:5J�^N8z��<t�k+"�מW^i~����uOф�%�G�����A�����;O�	yr�sm���[���<�Mݑ�~����bCH|�Z�0%�=�i4�d����5F��<asH����Nc3�_�(CK��N����V��":� �������Հ�2�⏡#�6�Z��� 㕨x�7>Hx���%����Lx̾܄jr�gb�юL�1$���`��
�$?C�(�mP�����4���_n�4b��q����(9~�D��[�M͚Dd@�NLX��oG�E�a��O�cGk��@�������7x���#�H�۾��\q�^`W���##.~і�;@5pAM� W�'�������V���f�1y��p3�/�xX3)r�qi/�k�+g�[B��Ͱ06��8��r��d|d���$�
�=���X��Z�jS@��`�Me���- Ɛ�Y����AA���K��)�BE�/��@חglo�x��0�҉\��� �+i�>c�������� �W�!oF �O\�/�'�%Jk6�I�L�6�T]~��,4��q'���#����ͥy��ia̜�ɔ�e��B�[�� ��Vr����$�f��并���->��057f�_�@g�t,��O��ѭZ�XC�ٙK[���H��AzA�B{�Daە��86���q���h���oDm"��M���8������O�`�̃�ÿ\�lq�[LU�by|��L�8>���a����o�h���B�"������~��?:{'�i�4Wn�<\�@��ȥ�;�k��}e�{~����H�+���f�Pb�z�~"R��,mP�� �78�]���JI����+�v^Bn�H�"`�c��(��kZ�S�z5��M��ωK3B�����N�S�f�g�{_����vu��I�ה�Qz�'�܌����/��}3��	�u�g/5��
� ((
M�޽0+ {Z��뾝�3��6&k�J�X�k�ឥ����p�£%�x![������Om��Y�����z��2W;,��Z��	KHc/��s�[�{��>����S��A��(Ī��p�n��qܹ��	�f	�N7�(@P�x��.�H��Ϣ;��N>�`D�Eh<���)�H�g~��ڛ*�:~G�ώ� ��>Ž��E\ |�D%�`9�!SC��^jx.������*�Yt6����}��2�)��8jǈ�I�d���8���^j�����ޘ̩�&�.k�@�3$3~I�ۂ�L����$��3��u���)�	["�uQ��Юڨo��5o8	��Ὶp�FFޅj����T�8�A]N���^�\�k5��9橄mz)3RH2��M�EȖ�`���2��+7����O��1:z�
�W���2�����ڦd���ϋ>�T���?���!�}�M��~��%�y��0u̸|�e{L�:�A���֎L������߼תD?�Xk��,
�'*�*���-�1(C���ϧ�\�%)� ޟָ��Nt�Ј�kT���n����S36􌖓��ִ�>'YQ����"U�NW@�x�M���]j�����H�|4g�3h�gU�{��2==�sU铍��Cn�xi�بu��]x�@�n� 5��,�nO��� ^6�˖ك��\)�GV|�T��/!�_4èV,üi.?��-�ͭ@����
����zV���H'��E07�����̭/����ۂ��ߓa@��D�_�/|��fG~��E�
�a����Ї�����GV�C����s�4��x����Pƌ`�����|�g`wR沄�ttjM���e,��ǔ~�>�ߏ
kd���)�b.��l�~�dU�i~�<��sUgX~v4��*�׷<c�����`�M'����4jP�w�᡺��jl��y�
��zЊ@�ׄ�
�F=�������2��le.���IvkV�	�6�א�\���Z� �9��u¹�O)�k�O΍�W��w:�� ���ʲ㪞�/
 �S��3���~�PDjlx1�s���%���׶?յ���GX���c���U�J�ƪ��r�c�R�i2>�{K3���]LV��	K��_�Ͼ�S��c���0?Y�Lm�l��\�8�2e�/]�!S���1>�z%���u��K��@r̠ޥ��;ο�^�����%܉H�3<T��8A�hjF
���c*pK��p8z9�
o�N	7	�%8�#�4w����M|$��!/4Z�L��i�#���'����y�Y�ĭ��K�(1DR��@9��P���b�	��0�q4Tj3`��������(�|� i��+�������)�&�#Ú4�E�3�!T�B?3���K�8q^t�Q�ٹf�V���$�q�')fVҔ���i�j+�$ �5R�n:�j�f o��r�6�޿h�	�m��/���iU�SƯ�.����K�T�N��v�5#_�h.=g6�0���C-�hD�щM�Z��iF�x�u���+���;ϓZ�U��͕4��8�
Ny�V�����â��f[S�
B������$�������p[csD�k����/�O�Q�?��g���=J��4���"�?ZT�g�"���7��C�B`U,���`������Snr�k/�E7�QR�Y���4wN�Z�b����Oq?��{����3ە����[��G�l�jl����v��-�|U�~�%����/�_��Ѿ�/�㉛�������\� �� ���i�̸q'7Ǥ3w�P�K�CZٗ+x���\���U.���=�CE2�,NH��V+�!⪖!�<����/���_;B*(��=5۩��x{�x�;��?�Ǘ���6kDK�bU@��~^g���5o��D)6cx�_�|$�,���{F�R<���D���ڌО���������nj�l��膮�q�(�B,�wj���\ʼ8��:��,B��o#���+� n���&�U/��(�qC�Yn=��,/�}?r\LLyɨލ� B<�ӥ�y_�]/t����˺c�C��F�*�����y��{��B���'��`���O�%o�(�7���8!Ǥ�u��:���GY�����m�VE�`�����WbP-�6R�#��6[2�=� �ن m�f�ړ���������������q�H"S�K���ǿ0a�9Nc��t�E��vg|��o1����Z��q~c��G�)j����tð_���0��J���A�5��?���a��x�g���{#�Q,kgH(\v�|��Yl�&��Q�Ǐ��}��Ҟ���O��;s1�j;�%T�<�t���9�	��!�����pu�;����R*(h�8Zj(#^���[r�1������W�ָ�#|K%��K5&�+^o�,����_�d[T=qk vۊS���s�B�I�Gf{9F������0��?S��ꂭ� �d"��pg_�tn���q3>�>E�Fі�&�lRp����[��~<	�	��s���+�m�>;�?�y/p�}w�Wkj��J�7}2#ӕ�YVҶ�>�\Fxj9���01�D����L�j���A��u/�?]�YU�'g�ə�pgn�@�[�@�o9Old��|Ќ<�<�³������Է��0����Lr#S�y/�/��Qk���B������𤍧&j�$�Q^��˄<�.����G�/x�p����6���Ҏ��N�d��J�nek� ����D4 �Rg?�B!��?�s���giiMɽ�-��_��$]	U�?m4��b��C>3�}!������a�N�ъG��cdl-\��=';����w�Y��=v\
76h��١l#$�l��I��Bbe���B��b��CV���& �$z�n��l��HN_1���7�~�N�y�l �q�U.���
j:6 xh�����UTy��GD8��_�7�tI�I���r���N��]�����z�\���ZY��3�-vt��)�b���)
	��櫇�Ȇ�B����%�4d�0�t�q����"�)����c�	_Wh^d(ɮ�1q���rقk⥮���IM����W���B��6,(c��H�݊U��8���v#+Z�NC~D㎨
��.8%�~4:���֦�r߼��v��*��s������8ʈ4 cWX��UkgueV�S��%�����G��aC��I4؃��'UXaPk�G6�6�c �W*�p˜c,Q�d��K�oV�����]0+9�	_��P(�+��}*�u�4�,��c���H�;����M��{eA�|+�(]*���Ԍ�B�e
����O\$D�v���H�j	�j�M4�GF�N.�9��x�{ �I��o�گ�s���]��:����iQ��2!��kKb�F�-�����V����* xR\�u:.�kQj?q���-�>�t�ga�5���'w�^݄�W!|{i'
D���rf�V[��g� �}e�'|o�"��A|iw��$ _�������r���29�?-����ʵ�v,~RC�������a�TM����}u��sוң���r4��vq݅��'�jS�w�åHF�Z�\B�x'%�BY�eL9Bup�H�\':�7N��~���ml�z��f���j�41���*𻾴Ri!t��&>�5�/��\]>��U���<����p�V���
a�C�CYD(6#��WzY�B�>��^Zir q�L�u�*\�ޡ�뇧�قd1�H�R����w�����%�нk�7̡X�2LE��p�6���dL�?�&%��%�u�i/�C�ˣ�,*6l�	�̈��~���o���OW����5�$�l{�^<2���0�����δ�A(T�ᱜjR~E�d<u�5?�a��Hv,V�p�&R#8��Yvd��Y�4<���q�g<NT����?�&�����QI��#mqb���y6�g�:���0��%�`T-�<�{���w#Mh���n��TT�!�*sc`�F=��u�(	��DHA^�i��M�O[�q�*���}q�9�{/Ǚ_-m�0�����W���&VJ.�[s��gk��H �ڻ}�u�v$�M�{�c�o��0%�rn5��-Q�b#�G~a�IE>�}�Ys|�A�ゥ�>�2%|�˖���չD�OW��=̾J=��a�S@�"97`�����]�/)�C�Uq��b{�1[��֛s��4d2^>CA�x=�z�i���T��)��񔲏(��T�sb�C���
˪
tt�"����@���v��Ko9�WO��:����Z+��HeI���qqk�<h�F�=o��6Γk1�Gc_Qt�A8��J0D�~��G��-�2���c!�����ܣC	��|��J��,nC�m��é�J�Vs)��צ���J��	D�8~�eK}��v��̴T�Q�wgo��mR�$F.W�֬���bg��}'k�ݙa{N��:�����q�������V�;�e_zX�Q�O�[�B֝�K�!�B��&3+�9�KZ'��eGUm����΢�N.3�+�8$)�*�~�=�:�>�/��zl�sB�#[����`T�Xs�x���?��c#�.I�ve7��u��9��t/�FXV�=���6�=J�N�~	h�F-��K�cB8'r;-	�Dc�~ǍF���-W�!�Z�I��ť-��f��eJ��K���V?�=���G<lw5_c��{��0JT�C����0�%�X�%��G�|���<�n�P��-
Y	�A����N�X\Bds��^��B"�2��O*l��ޡd5��G�Ȝ�zbG��<��m��S�gq�݈��`ic���f�-��t+�7��}&����G;���7\f�H-�i),��{s�hͥ�3�9�+�?���zV?⎅r�[bΒD�>��5��t�a�@#n��1Q�ش�H��h�ɠ���u�b��t@K����O�wL�i^�4�j�9l)8�,o� A��=͸���l���#³�"ҵ{��B��rz(��� �5�{��f7�a_�4螘�1x|������[���k�� [#Q���Ku�pG/u���cX�u`&#k��I����'�@xۡ2���|W�(9ԃ0�v ���Mf���z�1U����A����!��3�C���� K����o0~��"r|�.#��Ӽ�O����$���+T4Eo?s%6���ϋ��R�S���K	����1|�/7����ƄA/cm��U�S�HBY�+ǊFC��;6�R�j�0���g8����yR/�l��Z��ۉ�ygQL?k�$���|Cm��$Y�R�H��T}�(�uU�y3N.�>�xJ��by�7�<i�.�¾u!��EI�)�I��;YdvPƐ��ײ��rf����}J]�t����.l UȮ��7�(4�~�u��<�/�8�H,��I�����𜌅�hB��f�XY__5��\
_��Hط����qǹ�6�*iT��}��oզW7�Pc���"(i�~k��X��x.?�-~�j0�f�ъ y��h=�b&���8|��]\*�K�!�u�3ˢߑ[Z,!r۠��D��z�;���[��5�:�������9
_jh��-UhV����[8�?�xi��<G�a,��8x>�o�<�3o��!Z�4ߒ�$6&�Q�o�C3��TDV���7�L���[S��5~`y������Ђ6�Ik-gX�����ۘ��u���+���U�l�+y,8�C�+v�p��lCh�(�^��)���B�^D<����;��#��&�* @兵F�לOڂ<�o�G���R�Wz�hLy�C٤��7�J��b	pT﯍�E.�xJ>'�N�H�����$�)���$O���Z�XVRP�q����  )����p����PQ ����n��'
�����"A/鹌Yʮu��i"z����I��r�J�cj������05�16�XR|dw}�_�g;볬�. (�0�p���Y7�z�wR<J��G����Z���`�~ZTn8H��Pp�dnY�ut���ߌs���Vꢆ>�ta0'ڠ��4"�U$��Cܯ�
��Y��o��N�e���F���_[SZ�=���҅�*�`��W��cԁሕ�����������_��Ɗ�y��IQ:��W�r�������6�x�� K\̍�/�~�X��˄�+�[nQ�	�Y�dv���.|��JyL�L/��w҃��i�Y�s�s�b�n�ƨ]�/�s�(B�K���j��|E��~~�Jd����Tt�vJ�,�Z���}
��n�VU�k��<�̩�v�v����l����,]̘'�<q�O}m��n��QY��<`����8�#M���.����'mj}#�� QG�?�� Hr���?�Y>����6fo�;%V���ɻ{2+<6S�$�O���� ����Y�O����اtѤ�v5�R_�gN~o�T�;�]{F���h;���Aw���X�̒��j>�u��~Gk��Z�,�_,���Fu@��[K�p���0?��XD=� <�]""�O7{�
֩U�w-�ȡ�{�+WWZ�i�HP�%��͙�����]� B�����M���	��(h���5�x�y_�7N%�4`�b���$�2��@ĢsL�*훌��[Hl���$W�H[��S�ެ�Լ��4�jjad_w�P�+��؍�&s�{�����Ew���d��1�[��GD���> ��)����Ytn��m�`�}>��;�P��)O�Թkդ +������`�_��Ϫ<�pB�Ͳң��"���%��ë�V3փ��_@֕ut�ް�b����ӑ�����V��:{�d��򬚇GI��@����gZ�:��tt_�u��0=���k��J�g����l�
qHpV�>ać%J�vrc? oEΠ���H��P�	��'�[;����oHq��Q}����t&RE�]J�
�׻��g��W�\����<%�']�'G��2?r1)�g��TiH��z䙹����2Ok	���0��j��
 w>q�!E�8�a^hd8~��gW=�R�T�k�e@-����Y�����o���7�n<wl�'�E�����>඘Lui��W\5�zDU�V%N�O  �l Z{Gѷ>�����7�R/�;͐���/z#`�8�p4M���Hv'ωu�O����|p�nh
e�!��HAs
�i����paT���u�/��h��~>;krt�b�Gb�	��qq��[�1ƸZ���w_�ם��? *e-�����dFH�r��]Bz��`��8z����Ə����ux	���c�[[D1B̪�'��a0���ϗ���&�/���Wm��c[`){�Cڏ�f����4e#�LK�j�|����x!69�Q|��g7�6=��5X�`HמE9��K'	�h6�"tL��c��E��>�2���Q��]{���IҍCƢh"�˃�B�z����Kރ2�)�G�Q�=ҦÊ�wU�m�ی"��/��	t-�ɚT%c4sdnCb4&���`�?��	�<�g0s���z?��Qε<�a�ЋY����qd8#��1�
4eSQ\�?`�5DVW�;�����T��1{�O19t˶-�Beԛ��kJ��=�7�vB��*?�d�{��x�k;����U�a�����rkbMNK/,em�[�'��K�/�{4��+u���"R�US�:	�R�w���� �t�t��p(0
AWx�zÛ.ܸ�3�<A���cE�0��S�S7/���L���z�9��̩��dEDi�k�e��������a0�<d�?� ���4��O�v�)�4o�� 9w��E�9��2��eZ��kV:���(T'��s)\ ����<�t �)��;P��������=�*��b��p-�&u�\�O~Qն�/_\�d�,��:�^̼�_?��ů�"#��kY�f�!L|D]���=�����}L��c��sq�>k��S'G��j3CSQ�4���%Z��_fC��i�f�XɩS�����	bM�ګ@���ã�9����;E��7�!������dX0�޵{�x(@���LG��{�/5�J���7] wn�12gI�!����{�'s�ՓM����
�T,5�wY�eDǨ�ݜ~�q@��kZ(�������.VGI<�cQ\=�B��������}I�����)�& �m���*�78d�1��T�Q
cb����>�O��q�1N{Z�%Ҳg9�Ƨ��U���o�=<��:8����y���Vb\�S�w�꘱�xdb����*M�1,�'=b͢�r�/b����DH�����((�����I���X��̬����]��)�KaU��@���]u����%θa���i@�D�;*���g98���CRF(b�l<TP�-�y�P��I�k�=8
(��k�R�x��J�N
��u�2ws�e��ʺ�Wh���$J7kwB�+FA�d��^�ru��N8� 7�x����9J$��hƼIc��������u�P�J��X;�"�񫄖5��C;�lB�zdR�"������XM��	�ř5'����P�]e�[ 	��$m�,���Q�ލj[�qY)�_���!��a��w�0Q�%���O�;�@X��l� �@d�����W� �r�����`2�"���Htar���q=���3l�Bu�F��4H7�N��xV<+4��jDQ
 ����l=�����Z�U��l�c�:[�E�t IP���EBm�h *�O�Q����0�GE��M�/�_�gG��-�@x��ܒ0����V���C��K�rs&Ī�O\�H)g~ I���'�Sw���۷D������Y��
I ��1A�����U�5�5$B�:�oq� �c^bs���y��}���i�JG'�߇t��%�ˁ����X\�H6s����[�i��Iv ��eT=c���Q�g�ގ4
�T����;��|���v�|S6�&�D��f�u�j�Y駠�`g&�4dڌ76C����$c��9���5�9��u��Z١�/���g�0�w���т�:�p5r\'=^CN �eJ��nt�t@�XO��u��j��[>?fВ>lS��e\	�H?�)�p{�.3��jdO����ŷq���J.(G�J���=*mQ�{�3�K�T�=y��>�jC��k�9��T�9"��Hϸ��~���zV@�
MN�E�=<xx��`��q�FrfY�cH�C$/���J���a�Y����kKXiD�$���!��Z�����I�:��X������sCF2�s��]�uz�A�`� ��g��A����!h�o��fѶ�6��H����e#����l��$�L��JoVǇR�&%E�9��2�I���U��7͡s�4����������6M�.a�G���U\+z�X��i�t��w{���d*Q�_.�k��<���B�8R�X,���(��"�Ѽ/B��u���H�%�e}bӇyĮ�n�Y_���
�Iȕj��L5������)3�IT���I9���pҰ�Xg<[�y!�s�_"k-��G�CXF��݂���V������l�eY���,~zmȅN���y��9�0h��ĵ8���7��IO2��v��wgDC�T7�1�v���h�Ӣ9�J y�,[@(֝�I],��*J�اId���O�u��dpg�D_W�Mt������zoF��a���d��d ���$�n��!��Js�U��rv�&��a30�t��9�)��ʼ�]�SF�x�Y��0�T+�|���z�Z�٠豍D����Qg�V�ڬ�J"ӹ���NO�];�*�vW�ϴ�Y�2�{��x�� �����g�ktR�l2�-��C�vI�KX1? #7K=��¸I��C�/lA|��*�%h�7�]���,��Gτ�(nC"sy�8�i?����}�)}�a55���G6�l�gV���n�lA5�/`���A�������=v�`Q��R��$-�X��[Yg�{��qv��)�P��Q0�{���ɤ8��dxX�����Ӧ}����q��u:�t�;8�QV#M�$KRG+��
�L����9O3�Q�D҇i;|STR�'i�J�)GW����'��'Y��ib�j��Ш�9#��U���9!��m6I?�j���q����G"�N�+�E���I{ b/W�`3<����[�`s�_2�M!X��DN��$"���%穒l5������X�}�{&�%�I����Ja���,ٻ�,�e�HUj6��t|0�~�k�@��9$�z�k`��묽/�Q҆!�1A�b�p��%M�b1��.��-b��E`?����G�U��p��ް�w�I|��ԡҎ���,��W���a'qi P�%�lC�G7^+��n1�3z26~��0OTP���X�9j�㰙t�bZ�A�vF�z�T�l˳3l��;�ߦ�Z�p�ՠ����W-i]��f��B>Z1W�tg��M�G�����NM�[-�V�h8��t���%�u�����xH��nG|qn��ЌL��[d�����^LH�ˠ�V������P݉O�|����������m5�� pq�=k���÷8ռ�!S����	2˓f¡0"\�[���\ mk�Y����Ĳ�Ѷߙ�b�<Ɩm���_��!�@�>a6�����6!�=��C�.�~����̸`o�Trׂ�2w��.[�Jx|l`N	4x���@$�� `Al*��-����	��y)7DD�h�Rl3��t��Jq@��b۲���u�;_�Ǌ��ޜd�J-���21U�W��.��|b=��C(�B����G�߇�[���P��	׹�'���fbc �3�K�}������F� �y��i��'�z�����Qm�_��gT?�j��|'=�Ӻ[s�5H?��wT��sIc��'n �@��Q&�o���.��:�})oq���	E�<n
�i%=u?om6Y��`��Qg��;$�Q�2���p�)@v%;������]���Z:����~�Bp��9c�xk��ؚa�ͫ�U��Խ���Q���a�_/D��
���\"ɣ��*�ʗ�Rt2�p�=���lH��K�� ��$*�8���=�^�J�b;lr�wM�_�x�O�I�5}�Y�1�Ɲ���S<2(��O�p�T�L�.�+o�-�f�!	�z��,)z���`���˅z�ܻI�
���NV1KM�q��c�0�IH �r�%�ܹZMs]��e�6�Zڼ��fc��&�&�3��C/,�5�ٙQ1J�[:*G'X���4�CϹ�}f®�z/�Yu�Y�Tܵd2��"�BݶeD�(��!��z���
�o��[�{�v�2p[��s��QN/m��"��1(�j��*�2E&�x�?����H0�ʴ���Mc����o���r�0o�K���:f��*!}�+��N��Z�4�^ZͺH��P 3U��nf��G-�m�ԡ��8X�HG�����/0C���2D *3�0���:�Mc��Ż�m�C6�1ūq��&�#h��u&�t�
��1&�b������?S��R���{(��ѥ�E�m��փmY��k��ZP�����V��|�]���<ґ�2�PagAZ�vR�%�f�d�	 "a�JԔ�]���S�,���:�=v$F�+QضZ��#n_��m��iN�S���9�4[��e�NaYdM�q]0��2@�6W_��Y��\��;�b���x8�}	�2��@F!���)5eDWw"�B,�����ߺJ�w1�d}�@�'�:�ՏZ���g�r�\�V/�:Uԟ��!u�}%/��~E-�
�N�KH�y��s��_:}�S�Wx]�韭4HFK�x�ڧp��a�;�T�`���x���,��0�9e�ZJ� ����e����2'�b��n Ǧiu@��B�Ѽ]������Lu��zl��?v9��#���np��-���Ө,�n��>������T�� ĭ��o08�̘
L�*Λe�4�;�R
S�|�'��!QN&K$qK��m�)�E?� �QP��� I+�B�b4گ�)�O$5�R䊭��a?^�t�A���w�y��\-�g��`�A[ZP�B.k~��h����>O��1g#{uB=���&�H�Ɲ����D�.�_-�ꓖ�-�^�Y�A�HS����K��թ6��{�~�V�\ml(��qc+a��f���k�</htOR�`���sn�7�#����|�M��* $�8�����e�/�*��53a�]����a��lV�𣴑4��c����FZ�Y��k���p��#p@��WU�p9�;�-Ҁ������NC� ^zNq�BU9�#�D4aa��I��	�P۞���s�N�O�\������>t��ñhj���W`�����I�ãӆ�Ӷ�"���V����09����[ʒ�ݱJ�Et��&2+�I����v��J�.����$`�� �r9�t;0�4��D�=j&j=���6����;��h�.�dc���v�������ܫ�Ң$d�4�^�d'��F��o��Y��%�F(�6�F�S��^<�']{����A$8�a�g&�&�rP�_G��EA�S�c�v�u��A*2�쫿S}�X(Ŏ[}��L��o�a�F{���N��{�5f_=B��PY�@�����b�x�T�Y�wr$A��̠>v�,��Qm!W}P��8�v���x:�L�q���A�g�̤G�گ�`��	�c�ݭ�ӟz߃�R6��ʽ��Fs����q��TZ:$���そ�+�,����\hg#/����py��_�VG=荫��H���X��Z]��X��j�Q�.!�$�����/.�v2���c�N��JO�^O�+���9�<�<4��K��2m�)���_�=o�
�v�K>\��,�AQG*�| P�����r�
 ����14��� D�iI�����I'�칂c��EZz���qﭾ�FT.1c�G ���W���Dr6Cg���o�V���.�A������ݩ���}��`��F���� =��
��Mz�ƙ`d*�B�aO�p��Gĭ�����{:��������c�g��,:*����0s�KH*)��?�����k7�~��/#8���8����oP�>�"�y���D�n?mH� gYd����w-��P��:#��o�[� ~2b�:I�v�Ң���!�l_�V�{�����[�:q>��[������t�I=���/�!(V�Q�N$/���K�y��1�;��'F�^�Pco�w�]9H%���+�5����쬞�Z���7���7cW���q��}�mm/aT�{B��FA��=�Or�+�zL�����:⎦�3���t��|+v
i��<�`N��\�*���
�6̉dxP�[�Q#�R9�[G�&z��hQ*������/ D�!k4����۳���s('.	Z�q�;���/���WÜ6~+c����cWg�hQ �k��O㰤OB�[+�f��c��e?C��h,��Y9ka�p7>��Gt~3�=D��+�5��T����<���^�F�fŚ+C+4��A��˒I��Y�5��!pϡ��(��1����g\��W~�S	��ۇ�G�ǯ���h&{jxlnXM�W'm�6���Et j�}]�KB1a4y��$��r���d��4o;Mg ���;�<���%M�FN�ڶ"��ڜx�*O'�U@m�D:�!�s�ʩv�Z�bT�j3�0��D����|@�Y�J�N	�7��Ь�4�o�̀[ŅG��?�63Rh��Ä&�2�S�h�K�;sP��k�P�>�*�KkS�;{tm�X?
�ܣ�0�M�ܞ�\���v���e#_K��'���q�A����*jOO��F_$�b�]�\�B��Պ@j���£��n���}Z�C[2�P��j��8^���;�2���ӷ�HC�����ٸ:�ƚ9\�b���.!.���G�d8X�
����� /��2�&y�on4��J�لSlA�So���r���j�;w�8�-��0^j��پvf�^Du���_Ol��,��(��*���+��n�͛��GO ��A ���ߴ+�F�F�9b ���T����<���ѯ��j�t��=>��RdW!q)6Wڻ�Sn�����_	��w�#8��>~)ڠ�S%xJ���+���1L��kj �#�D�1��3�	���qQ��σ�ʞw�[l�v"���{�	q��#��K}m���o5�t��FwR-���q9�����(e�D��ב_pM��XPxn�X�i$l�X��FN`���N;�0FΉW�l'3~�$��{&�P�rc�rc�j����x�af��J�o�8T߱������f�tR�>���gTƃITYHш���.�X�;AanI�U�t��/���9(���a�T�Y.0�H��S_�{@�E��~�.`��s���: -�0�t��X�F8�
Ņ����WZ��d�|E�R�U��FƵ�㧭��e��FL��ځb��3^$��ԨV<<̓A͊&#tM/�[�~1}t> \j׽	��>0�K����qHӍtA	X��z�	�G�DTqe��w8M=K�@��
�S�L�����~�!Ù�BP{�7�'�}�¾T�5�Ǒ�b߭�]��	Z��[1lH�P�_p��Y����nۗ9g6/DHb�� \���NNL���/�	UZٸ#��y꧌�o<q_��l��x$�=4���%���޽>�4H��A��ŋ�>�:c)�6�x�XK;+ޑ�����
��O|�N�3���?��������b�2��ؚ�:�93���#Q�Y��N��->~ti��,5cxL_�(��mr�|\84�ֽG@Mqx�2z�R�6ٕ���8MB����̇r�4�G��p�}X�[l4�h����>�w�%XR���?�Y����!��R�?[������e�cx0�H���s��^ߨ�K����;7����"V�S&�mb�	��e.�֓�<�/�Ξw��5�2��N�W9�"�N)���0-!9����N����kXxI$i������t�%�T6O��_u*^�.���jf\���Z����I���\�7�_|�M��o�T.�k��He{8}yM�,�=�R䀴���|�*%�|�jp��/t�BQ�l�%�he����z%�a�qC�A����V�ns@�ԉT�y����c����r�Hn��O4���!4%�R��q�8a�Y��X��BnK:pJ�ys�߷�������3�e��k��V�ǻ��k�z0>���>q5b��]�}w^����@���[�S9�K\C���s�ҧ�� x0p��+�na�`٨ِ�C�,���\-��s���WZ�Ƿ��	R������-�mh��������1��՗��� C0f+l��A#�ߓذ�)ߋ��yo��1��B�u:}��l<fb��5�>��f	��z��r����Y,y��v� ��oq)��ws6рb�"�dsv���c/�P����~�Ί��-F��L��	�4n�kK�7�#��F�b�u�#Mꆷj���>{|��5%N�=C36ja(�ش��(��%�`9���\���^�S�_O�3���A�<Oln0���人oH����I�.�8�u%8wH�'[�j��@[��R��8.�CR�'�����J��]�!c��w�Ԅ�B�v�T��B����E��'�1�C&��}��a�p���ajŖ��O���[@Q���|�i_ڛmT��q_c@�I���j#�5�r�� ����v�� Q4�Z/TTY2.�o��UBE
!�c9��$\�)�CA	�U���p�xJM.��G��U��t �Ƀݬ(`�zMт6D#z�_m��<�C�^�e��2�0�"�-SO����=腒ZL(��f*ׇ�5S)V�K�8UD.D
�"AC�cw�f�|���S�k�4i�����)H�6�Y�������V`�`�|j��o��x��M-���29O�'x�!:�E24c�$�
���ܘ~���
`�)�1d��i��ۆ�U/�p��@W�xX��G��0�}�� 8�؀��I���P.br#V ֵ����������F\��& ���	���x�'-�V&Ӿ4O�J�Fj��{G��A外:�v���ܿ1Pœ���Ii�G@-�����Lp/v��_k@�\evs.�K�V��v�9�?w;s��UJH���Z齟o�e����i�<DHQ��,bQU�A�nU���:�b!I�3�CQDB�s��߫md��G,���Ά��ۄ��R�V���tJ�,+3�.�K�`��!i�z߁'���=Lxb�9ǋ��R���	>K�����X.�_Q%�/�ʜ�$U��-'�f�04-�yf�l ���ת[���Ս�Z�4RHY]���NKF�<C! ��	�36ӱI+{$�����&I7��F^�m�8�u�})��ϙa��׈���/�g{(�%W�@L�Gp�e��8��l��W�D�����f�瞋.o�R�.�?1M�e/��/������TX�g�H{�gꅽ?�	5�� V���a�,P��ZA���Q�5�\�%{��?�}ˍ�� fdAy�x��w�ߊ���q$f2�C}�{T�k��c%�2D!�`���LL�����Z{X"��#�{�YA��}f@��B����*sz��sSY��.�hI��m�c$T@��|���)�~T��L�.��	��YF�M��k��8��w�C6+���G��6��d�~�����V͠V'þ��_o<��3���	%�ـ�b��0��Gî'�j�2�"���I8�e���F8��j8m�^U��?�cS鈺V/�j�~^K��n�� ��!�^+�s�=�lpu(mAb���2C�'⫗�<��W��v��-	U�t�*љ����L�&�ǝ�̔	�\C�	E��+��8�Q��-�_T|`�D��-qD�x�+��X�ք�3p�M� 
rrG:jnϷ<p"�Ŝ5e����{g$�9H����!R������b�F2}�r�9;��%B�:�ˠ�ؐr/GZ��!}�z&�P����w6Y�8���[2��gX�pې���=|���0i6���9^
�n]�DFr�P%��.�q�1+O��Bh�����WK��_��kn�������ۖ�� �YlUh�	xW����HN�A|]�j!zQ�ahJW�b�-�ɠ���J�HB'��[�X�g����c<
���k�_�`��S|;-��c�?~�&o_�=%σ�&l;,���o����U����ķ�vP�3r!�����W`�C(�C���n�5��VD]�CK���!���n�8�v�?��_i~��U�{,-_���A+cq����:�D���Q=�p�Œ����9��F[P��>c��`��z^x�ٸ�aM�F�}���b� UW����C�c�4�]\x�ߖ�� ��bie\������b\���v����9wP����	b\-�J��ָ�$4[�1Qy,�=-�o-�����-��]p�]n��/hR�6g :I��Q�ؖ%��e�QQb�]Q	���B����\>��0UO��vB�}QtW�;g$�0j�c�1�^�-�	+�œ���h%�!����,�È�y>�d�v(2�ܛ��8��m;x��[��pV���w�ؿk'"����J�؞O��x��B��$��
�V�s+�PC�Y���-�d�f� In�%HH��<Q����=]�t�=y\�)۴7*-N�Vt\�48y�ZӞ�2��n̗o���~j���'}�(ŔCDnf�+�(\�? Y�ij7�8Ql�?F��f��|mؖ�8V�ldφI�B�B��ƶ�9�C\M��m��r����F_H�@=�o����x�i���%r#�Y�g�L�0��<�X�%�S�#�y�	���1�'�U�U���@�U�H��C��`
�$x=����l��<o���z#����p̺����;h�D��P�)��R#|H�k+->�����೛���K��i��.�u޿=�B���N+�Z19%���j��1V����uƕ�u��/��}j%���G�m�v ��CJs� 1�n�j�)�9S7]��+e��7�R�������ƋI��&C�����g_o��/EI����p��gv鮨�u��2��Q��;�h '�*%���RgJz��m�r#P@�:ME��M��z�3:�ǰR޺��+L>g{��\LA+Q�G�^� ��р@��祦$sg!
:I6��j��[���eaǷ��5�e�{Ҍ�P�S=��c��&ux�b��\p��QIi��Hb���.�eꎢ]	8�kv8�Lz��>z�������u*���(�x� ��p�H)�,"��k+Z��$��<��y#�w���<�@�j��Zv�q>ݙ֞N+�w�*��(kiX�*'�����den���x�vWu�b�|�ޡ)PiK(��yխ���ʋ1i������{�+"��k8uroć���k���cKL9��"�����S��;W���G��b�!\"�
"N��ϑ�w{m3����o�i8��Kb�@�m�P�I����S�(��J{6����W�6� ��?=�"��H���UU��C��ZP:)veH��D�����)�Mi����3���ʒ�Zm�t��"���c(�F�,:����r��B�}~! ;��jxn���A(��t�t1mew��b|7�ߢuX�Hy��j�E�2噚�)��s牐c��ϯz��GؾPK5��e�0������~��x+�L�2$����3�,2�����,��|�'�Ap|�
?�>3�Rɏ��~��=�e<��k*��h�})F�8��7�A��s���/��Ϡ�'�$2Ŷ��R]����s�~ ^�N�q,�(i�(�T�ѭ\���她���@��BV^��6 }"��bD������M���4z�]�TW�����/SډX����"�����	>�[���{���G2���E�-I�j��%H`a����=Q���2B�xyjL�5�Y���4M��?՚��z!]-�����B�
U���x8̧�{�g�*SĤ��^"�0't�i��Ѣt��-U/DKi�:��oQ��K��bOe����)�� ��CzJA��vu���B�`�t/Y�b��}��@]�`�wڪ��.���d���o������:Ϙ���� &\���Pm{\8Ձ�����6-� Έ�o�`�����Y�ѡ������bLV˭ΞQ!n
��O4�
�ՠk3�6f�9a?5Ѱ*�����Rɘ���\�W�eV�Y�����Gƶ�Ӡ�z�̐� *���u�2�;qz��^�}��$q���^�!����2���]�ٸ�g�Á��#�&� D1��w�rt��E��5">T��$$�C_.R윸5�v̬&Gw���5VQ���k�5��H�Σ�,�E�}��yqv�2>��cن-%˕��d�N>wV�@�1��~e���\'���b�L$�Պ�Иa���m�����Ѽ nD��*�;0������2�qC�)�����׻�׈DEsC��N�,�h���M������l�ͥlzjЬoB��Wi��t�>_�)2�Mq�B�ݑ1���C�I��Ķ�lޮ���]�u沧�!Ö��c�Sr)K~s|,A��S���
�@��	���m��a�f���I�C@����&���Ïo��a:��)=W�S�UC�h�Z�G�D˞��-���^�`�����p�����魑U}'q��A8�!�����h%ύ��)���!^�XK��Uo�*ؑ$���   i���~!��It]��G��\v�b=
�9aS��z�@�>�&��r\A�5���O�`L6�Do��r���S��GDt��&U?4��΍*�)���~�۴x)���[���7���,�b�oRL��3����nd��nlĈ-ۀ���uA�0���-��,*e��=.xȮ0c����rX����!d��I|��4}&�_&��P<Â��|̊����mm�k��k�u����oh�a����~�E��)8+��w�!�̛C����3#��/��i�Y:i�3(�oeB��J�R[-�fa
d�!�W��rPva~�QG5��gU~#�|����[�J��N�ܗ�P�8lT���#kK�Qi�ɓ��dBW��Mcf�?RM�e���<�@=�S��	˸~�ժ G0���[������AW�"��q{��I�6�ϰ�{��bɼ8��b		9�J�ǎPr1���m��=
�A�7̽/�y/�&n�_�/<⭰S�{�en�B�����k��(B@��ݥ�:"Ǌ����1�u�U�H -c��Tr䦉�|i�d���嘓x��{ȵ��t����.g��xw�:��Ң
��_2�h0=l�F|0;fGx��V���-�ٹ���yܬ�� �؟�@�j/��aX��~*���M�#�,�
�A9�O���1�%�/J H�FJ�(�D��qT��ݚͦ���?Jr���' �Oζ��ba��~�:��a�G�i5�K�)7S�H�Ln��	���������=�w�7>+Y���R_:J':��I��8_S�#�@V��Dv|�<�C|�$;B�%�U��i[���%�o�xNG�KDQ�:ԍ:�ްda�O^Q>����NL��/4�G<�J~h���D>�P<�uebi�?��� s>oT�,�wB7�	���8�JF��NQVQ�$J�:��g`gj˫2P�>��7�4YL'L|e��v���2�����++�U��=���M�Xg��ٸ������C�n[�Dr8V{r�uv��Rgk]��8>�i�8��JrQ��>��o��#H�������ƷՕ��*��1���)B���@=$�ҙ6�O'���e�L��8�_^��&�E�:$��L�%��l>���'r��\e�t7,m�ϛ���~!9T��Oi��-����
q	 �qvg�v��:���R���g&�c�A:�N�5Ԛ�@�㗛ݿR&�̭��W��m��5�+=mې�����,m�nB��I
�aQ\�ks��'���9b����3k�y��BĔ}�u[�1k�|cm�W9������S_��B�-q��7���%?+���������fv�K%�\S'��?	�Pf�[��d؆<twj\�#���E�8H�?��L��,�/;ֳ3�v��t��X}q&�&C a?m+��1����n!��>��Ͱ+ʵ'Ei�7b��q�*;��-�:��Ɓu�C9I����X��)�)+̕j%ŦB*�"��>�����dl�"�	�m��C9�5��)�.��Bl6Q��~n�����(2/.��D�] "ܙ�j��QP�IR������>����~}�q���ܴ��bj%ȟ����p��]E�,��)4���Q!��"9}y-R�L{�ޘf�H Gç8�=���ќ��v!�^�\�^2�;L���|���[Q�+ff��us[���������<"��6Va: 0���?��@^@� �s�zH���9���L>Ҽ�L�4�\���� \el�a�|m$����$dC]]8���`]mUe��n��h�]p�Xkry�V�S�B��Nm:Ψ ��D�#?����
�;��#��s��W���u��Φ�2yQ6���.0?���_�C��P%C��']�x�26���3��7A���F8�25������Oo�:z�B�X�4Xj�s��^�N2s�q�b�E�~�9��;��S�F�D�	_z�XN��O��V���,��h��#�׊�u�
;z���a�4�}��P��U5ρ����]c��S�Pڶ^
��l+A��� :��e*{�$�N�	�elP�r'IH��"��+H%����5��S�3?9('��^Y��G�6�(�I�H�OVU�l�����<xzr��<��%���z>:a��D �Mp6�)�rM�U�q�vA(Q�KFhDN�m����eΔ9��-��Q�[��%�gA��;�"�:�)��M��%��������'�>0��t�9���W1��V��|�ŕYaWO[���@���hx�U�4��][�b,�f0����_��S]3x�X+$�nޚ�_N6�a��2e.����ܶ�_|�kkz�h��Opپ���2�@WQ"2B���Şs㡃�-��,-�CSo�"��J�j��V=Ẩ�]^��D&z��ߚ	=^N���ya'T��{�S�m�Ik\vʸw�+x����A�H���>��@���);¿(�iqq-���h��٨���7{[�����}P�%�XjH	k��!NV|�&� �>C���m��](Eq��Fie�r�VlU��Q$�!��U��Z�U����eR}|�$9�*S-�4�V�l��i9��]�j* x�Y�ah�Vǂ%�9w��{�C^<�W��,l!�vp�h�������`\��Y�_�����i��?j���v�9�xn}%�hc��UUL;MR��>.�O�~����ѫXY%�w�G�%���<�������ʋ�q`���g�#(�	��Q	�MEH�N�.�������ى/X��R=f<;���'���"�qP~w���]�D��9s�T�4�k�Z�ܐF;��C^�f�];܀DԖIN��K���|C�7u�&'[\N��"��_<Sp
�T���	�̾��{����f�Co�u�]P�!dn!/�^���Qt�E+uAR^�7��i�A��ӥ������^��s N!�<�m�0WK��imMP���4��0�f�K����'G��n�|�ښϜ��:r.B��HV1!�E��HsDQs��@�Sf %u�E�ȓ�R����D�<��?8myy���)G���	�#��P�[y���0֔q�k����El"�=�0F�i��Q9�JT"`��V�h�D�\�����k_Ό���gt#�M��PC[B�����^1aDA�7�8AT��a�&��rCA���j�r����sj��6��Æ�.�t��aK��_9�6��p�Vo����a�@����H#�'�no��\��+�Q��~5��t��J&�z��aKhz������ם#�����d!&�~������r�\X��.������%LP[�쮉��f��$7�b�ɏ��>���!�C�S).����Ni8-8�ҙ�n-$>����:ؑ}_O��g l�A&&��dm���B�"k���4�ۖ�-V�	�a����Y�.o�t��<�?r �ǹ��/5���tHX��20%9D6�^�����O�Ĉ?AA'���N��.��R�W��-Ǯ� �=��LbÇI���	e���T!DU���9�0	d%�F�f��t� a]����!���4-��IB	R~�Hr��It��VK�g{t�\8Exef&c�h��!��BщiDo!/��D	�;�I2�`h�ȇ�/c�=!�ͼÈ���T쵖�_;���4�kr��q���������d�Y��q0��Տ!��$�U�#�¢(zCl�	�x�� ���k�!I��p��]0���C�ɘ�����b�wUm:&t�O�Y�B����+��e��1�]P0������
Z�����/�a�z�䱓x0.�h���qHŠ��ϗ��/"5t}�����םw�C6f�� �7M����s���)U��+�zg��2���҇�w���D�!f#C"��EO�Y��k_��:�FE��o;N��!V��2��2c�����E��OZJ
����v<TY@��P�yw+\D��M��� �W�;>𕚐@2|e^�{����)2zj���U��ƛux��S��ݎ��g����9�v�WV\�:
�)�.Xhƶ_��ag�#GXGH��v˽9n6HЧK
.��rEW`�A5�\um@���2^x}�C���h^��	�i��������V���2$�;|E�0�/�M·κ�x��¥Cv����P3SIm�T,Y'��O�h�8q;<f"t1~tˆF��tu��xQ�$By=\��H�X��3l��ʮ0�!q�OVEʪ�V<v�K"c�5ėd�e�nJ�f���R#H]@�g�_���1�3|y���dtN&����"�:
/]A��j"�E.���>mW4�,,/�g��w��>����p�^1
�ȳ�LLa��<��`Ɣk��<���t=)���R_^�KM@2�d���A5b��n�E�jG��Ɛ}��������n]Q��n0{'�j��~��w���E���֐��"�]�w2Y7�х~(�\C��:�F ��%c$�?���K1X�o�:��>�I}�,D-��GƮ��=G=j ��,���'��+�	C�o�
���q\0��r�܊ʾ����p�;NFI2F�WJ5D��G2Y}Q��-�>�o�4�J�z�
<�e{*��'Qx�@;�2�=�įժ�����$������`-���θ�6X��*�ͅ�x[>��?w�-��/k׷���۷,���CO�5Cc�o�qE�UX�c������t +��V?�S\V9'����.���`�}U��Cy&�̜�@��
�n=���y���E�δ^�3;:��Ͻ����p閻otڝ�s������``�}$��q3���)��"	�d%0���:�v�V����TWY��Ǉ�*J~����M�e�g� ܃�55N�@�`aq1�=�O����7�|X�vNaB�h����s� ����N��ML �.0���.�&�&[���2��)x�H���f,�����2p!1�0ZH��q�|��G�i�c���
��� <7�jҐ1�����`}��V���j�@%�q/����DB�W�}l��*�W���->�om�1r%�k��mh���i���_]S��S`{�|y^�	ڼ����7Q
�E�z+j����s5��Y���|���H�^iP_��/����ps3�C���=�^�\,g��ZS�~
��\o��;��J*{���6������U>�8�����o�����D0��d�q�B���pQa!��~FQ�ط�6.em7ty-ߢ^B8�� �Mkv�[�|��(���	�� ��J��*���*E�!3��������a� 8c�-:(>��B�h1�]S{QlH:\�e��w�n�z�|��	S'Ƿ{W4D=PI�A�ԝ��M��@m��ۣ#�p�6-�"�Q�BPd�
��d��0A�8�y�$ǫI;��C����jˣ�[��
���!��[��Z�݂-Xz�������e>c���W�c��j(D�\��ed�u�/��~��k�
;��Z��������9���B`�zR�����Z�4�d�a�F�R>��pG$�t"]v���J�@��sT(������O�s\
�%�ցHi���G��(��O�w�pCC�T� [����-�T��T{���l�>���-���r|��E�:ū�CG���V5���iW�(�=êg��s&8�s��8�Q���p$a�ABY/�>7��PK�s�4v$�"O�ߞ=����s��S���iS���Z���f��
�Yh:O�}t���K8x)NKm+$z�2:��ۇ,���zVZ.�A9�A��,$^]�B��u2��w��}e��\���<�� 1ӷ��l�;���""��E �m�C~�m�B��Ґ�,�����W����)v6B�r�kug��
��{�oJ2A��o�#-��gO�GΦ����2���'�j��
\�^�]�0���*������Q&e@!~��J
��������J��"5����v^���8�_o��G�0!��
���y`ʟ���.u���,h8���P��%���i]&#��[��*$���gI���q'�I�2�`��N���$ly��a�k����h0ӆ���C��v�y˃�GHD�7�=�M����vT�w����/������Rݧ�|E�To��DW<o�:sD	гDK�0;�nD�|n�Ua0̟+!�^���l�� [���R����5|E	4�����N��J�ǻK�\��M5�ה�Â��4���E3�W�^Q��R�O�ŖH;Nq���T�zd�{|�m�f��|��]���f��Kߪ�[�b�~�����	����]��I��ؐ�=����G��r?d��h�>��U�̫8C�Q]0�,��S4g�*Ԟ�@M��t0xo(���+�6б����!�*�2��u,#^�l��[�
u=,[����t��u��i[;�`��i�Z��NK�(�?�l��H�b�Q���BJ|ѰM��i�T��#��+(�����i��'�F�r`�ޒ�̩�xI5��]Ke�x�{�" 7�!fX�f�Ik�ot�M~C���y�d�%����o��s��6�Y��y_�P;쥘��#q�l��Ǔt>��B%�k�	%��?46������1N�.J�8w�	���]�j��}Ϫ��?�)�˂�e��ᅜ�N"�QI�x����Y�5m.�?]I4��?H�O�O�
��Ҥf=�-N#��>wj٨���P,�� 죙�>I�	�����e�-��"_���ҕ~e%�#nS¥�^�N-{�ܶ��S䑄#G�P#�ye,�����F�gG5͕e�w[�<4�>��K�4,�/��p\�T���*���^t��>o��D6$n�<�z��0Eb���u9�S���rr��ݡ����X^Y��K�W��ez�����X���ID'��2g�K���ܼw ɺ��,I=Ȏ������&@%\BO;��B���a�L<�f<������ޭ�]�g�^固/�J�]�����-��v����E���:��!�&�4L�Ub�Z{GE�.���~����ߞ�[{DbL��1-X����2�>>�4���=mNa��;=V+�	(o�7{��ܢ�K�u�U(#�Xׯ��{m��ɢ����v-������2��|�U�Z����j��cä�HS4/S!�'e�+s����q�sB��o�M*����3*����B3����rN�-h��5e����6���u�ᾩ-���~������$��Ct8����~�T0��3w�*��Pt��R��*����7���
�rC�˫�=:	����ɬ%��^�}h�y�i��������d7dsV/���:��˝Pi���(ۜϓ��`/<�\����B����X��<+7�11Ü��s�\�|)���[���(�����WJ��i�E����宧�@j��A�<��:��p�"�pqUO���� Rl��S�*�u�M�z����ޕ�����e1��?M��IMr��1�X�@�C�f�t>��bMk��;q�=y�&�W���Gz0�X��|1�	o�3
 �q�}Ǿxκy���V��$��޴{'�t�OŀPj �d�6�m�5�j�;Ւ��A"����PͿW�w7��%����ڿ��K��*�= �˽����hr���`�Q�ʌ�qЛ׸Y�g.�)]%:M���8�RU�����,��?�9��MR��dYJy��NŎ�m0˶��y��W��*C�9��
�u�(~-%�%(�R�y���\)PNt&P�0-ԑ�RbA-��R-�"ʨW��m[-Y�BV�VN����d����V�ǆ%�qp8���:�M�����K�n�1���w��z���d^��ɖ}�ZY��]^ �ST�[��#`8�p�!���vPv��3��j]f�B'���J�-�X)�d�����dL��!�r����6�r��7�yk�K��L9o�)�r�����Ш6���6q'��L�r:���� �J�j�����)1�r���� Q���8��G�O�����+E3c����(H�uu,f!����P�`��H�"��nS_S�E K�80�Ġ��Cnt�q8���N�ז�N�GԣF�~�I>�vW;/'�$+�@���dҴ�f\͓����~�bY�2�>�H̒9aj��%�^�>�E��Tw;c��<�_���Z����(c��:�ݨe 9C ݵ\c\Q���E�����V֮xW��#Yp�ӵ]!���&-�.~k��D�h�߄�bD��Ǽ�(o����U�(p��<!˺�	�ˤ�. ���m�x��vV�����ͯ,koDB���R��߾�Mצ���̴��^p�_�O�	�h���Uq��3樈���<@p�.׵|�����wytY ԁj�ز`�8��5��op4�>Jp�*�C^����ΐ�����POs �4B�-C�z ���~��d9c�����Ff[����ڱ���N��k��
�zȋ$�Nʽ��;s^�J�<L>���Y����b��� ��4ЩlKw9�cDv�����uZb-M�7�7ɓQ���:�E;Rt,�Þ�U�%�����&�(�T]���ƣ7HH��n�2M�x��Y%R(�J��� ���$�n����f��mq�ir��d������<)f�.G�O���ck8�N�����i{D�S��j���|�)��s �jl����cT���q5��)�c�]���)�9B"x�LW������n���kv)�0��Pǖ��I���l��r�O�N�th�J��n��e?�)���)�`Ċ��jHr�,�/��Y�ȭQ-�1En�68�#��?p����M�I�9h�?�7-�ޞ�G(񅚵��<�&�'oS����h8	q��ԁ�G�*dE��n��|JN�ʴj�6�W�����ȃG�>ȃ�[�D2�~S��t��i/ވ��h R�1�N��yņ�K35[���Ё쮾g�9	(5C�_
��R���"�#��uZ��.�����E,-��.Gs�h_c��A��v���V����:��@[��4��$��2���f�m�����0��v6�I�b��=n���G�z�#e1ݞRc�My
K |��nzjfh�v� ��\B��������Es��W�*M�������WN�I��Z��&Þ<��������C��'���юB1
���Hk��KT��@Y�>䬾��AS�� C6ߣ"��7��$zJ/���τ�b{|��P���(dIe���Ì����2	�2�g�ۇfִ���ĀU��o%��t������S�*���U��je����)�>3V ��'����5{��`�R؞N�M�1�zѼ��m��-;u��A8�s�|�Ji#���� #{ɥ<2KL��uJ����[r���'D�.��鍖;٭�\'��i/|D!y�h���6��Uu&���]�dl��)�q+�����"k7[U>�u3[E���6l�QB�l��.�
pȀ*�yd^�:��Ϋ(�C�	�����w���c��XWe��.[�*�YS:in��r����x�����/藒%�a2x�w����  �?P%��6\�qN3��8�,���z�<d��FIM�I��N��/u�cRm�B)�����Ņ��� �Ňs!����g(3[J��h�5RPAG��|D��[��J5�$u�?��ģ��0�LO5�B"����_ɭ���
'�	y�)}䏦�^ƫ�ڲ�-Z%�<�`R�[�FJ��Im$*��%Id�͚��M�&�h��sp�MJ
ro6;'�X��h"��O���������f��"i�n�N�%��X\N�5ۙ�4��f�&����������YÚ�H�����+����k�R)���5�Y�F���� 
_���x�S�S��M���~Ϋ����(�U�-jC�1���ƻ3�J��a�U��i�ws�斎t��'�W���N���D����ZDVgW*���ۼP�~'���+��HO�YWaĵ�ő]a�LB�~xc���B���r@�2h8ȬZn��I3F���f{ $)Ii�f<��<�0�Q���ZM^�I�h�&�6�f/�"���i4o��F�N��Џ�R�.g�*���._$���y������R���H�6w�I��6���x���Dn#��3)EH�^���*�7�q3��[�O�V����IR��~��R�]Տz�L ��Ô
~!� \���#�J���-_8p�6���)���m���Ah��>(HB"��� >+���U"����/2ĝ�g�8���0c�|�!Bf|��DCo>���rR
nn�q�
�����o3$�7�w�Ѯ S�rd�b� ����IkL/1��t��U�M@>�2�e�xs9�fX���kbS�D�F���5��|�_�~���5����슚O:Q�a�[��*��D�-|�lJ�c���M�Lְ���
������Uߢ (mF�-���[��� ���פ�&�t��o�~��+�(ю(���}g����Ի(�� 26�Z�����Z1���*9o[�4�Z8~��l\C��I�k	�����a)�[3/� �6@#���m���\م�*d%ńNJk��h��k��2Yl���c�(�������4Fy��pm��?��"��pR$hO�E�fĹ��;�7�7=<!�9����h��Q�gkz��j�ǀO��tZ�x��\��.�����7AD����V�ı��{Eј�/��q�|O�&O3d2���cU��UɅ�0�Ĺ�����u)96���g�����U�/V(��DQ���X_�>ݡw���Ժ-��@$�E4�A�'���������';W���Rٰ��[� "J��n�58�!��6�@�W����q�S��z�:�_`��i$y���e�	��o��*!|�i�����zM���0����&<e
e
��@������[����ݙ<�Yvb�3�6'��|���mdQ���f�,�� AGX��s���[��P�����Lw|L�e��яEP���$o/�[/�Yo7֞��U�T'�`�R��]F�=}x������ᨽ)�Aͤ� �y�q�˙'�g����5����4���b����`[ى��`fʢ=�����
/L[~|g7jz�N�*����.\��ko%�x}gK�P�5�H5װ��d�q
�@��c=����ƛ�l��£8Q���ʼ߃��Q��ޥ\%�A!�j�%&�W��Jo�X�zwߪ8�Z�A����$s/�NEN�^��5~�$[y�_����`���1��Q���N�v��8��<���l�n�1�P�i��9J�̿w�s�% �o;�~?�f}zvayg"'��<�a�ʰ�5:�߇�'6�R�v��M��t9	�v]��N�K�D��,-�3T���3�(׼R˳��_��p�ļS�_��\<���U�:k�3�l0C�����0r�G��F�U<�!P�ik$��!�129��Q��%�ꮂ��rta��	��3j)]чj�� �߫3���_�ݏ�|9\��p��j���[�.c-Ն�	����o�ZPs�����C��݄wqs����o�����V�MX!������l̯���m_$o5`d����_��z��vI�N.�L5�y�d��83���8Yр>1���ԁJ1�J$��8A+5w+H��D�R�e1����h����N��������^r*J�#�H�K<�fזN�����Z�v�υH��n�s�A����FF�O� ����A_&0%U#}oW+���I�WN��K��~8�4���畓Zf�
�#�]��!&��V 9<se���m������<���a��bX��>��.kaQ_�x�m�$O䑦�/Bg����W���C ��7v�)�#	����7$^ΓC��`o
�a��T��G����YPw蔊���UN�Nz� �p%{w��BI+ҥɪ��1���6p�g�3b3�o�����Q�w����u�3�O�R�v
V�f���b�+��y�Mp8��z��
`��0�̫3�笚���)I"���e ݮ�B�to��]�Fp��:{cO�5p4U��wTo�h
��q֫1��]�����X��;&���4`Y����'R�K�IRp�#� v�}L0��o1d*�1��~t���q�M�2���He��@��Nl�StJ�Դ^�N�ظj���N+׭Uٷ �-�Q��dh�A/�أ5R�;PczR �/��G����:/�F''�4��b<H����ڣ�r0:i:s��B8��r�����Zy1""=>&�%:U+ѾV����'_��G��Tvz{"�����Q ��6ƭ�k��A�?�g�9{\�YuWb�G��ߛ��"G�
&D���'��D���mx��`eBej'U��(nl���:��l�
��q��_��#�=]N������������(N�*�CY��e��u�)c}������w}�P���'����̠]�˗%G��	z���>5�����x��b��������,���DΏh	d���7��Ĥ .Av@G��k���1�tn�K��m�2��Vs�Q�o&�֖��ykx\� Fs�'�E�0�E����ȱ��dJ���8��#sg�R��;5 ���LsYŽm�k���eФ�#�v��ܲ�^s�Z��\!����'Wd�}Ʉ�M���e����T�Q�"9#4�A�=���K� �'��eܮO�(i=�w�����($��`�?��R��X���(5��b
t��c����`18���
����
���N����Z����A�Q�BR��n�""�}2U�KE4Pj�qW5����n��`�%�05�K�ʔ��,X��6<���7�b�����Ų̾�*���m� ���k��^����`���`q-@V�áF�ږ��,��d,�)��$<�7�>��˖-Ys<�l|*������(_ sY�Ly���k鍓~ߎ�I��������| ���2I��3~�%�A�p�?�����+��MZ22�����b`����e�P��|{2F�"�z�"�V��?f����&#G�޲~=עEk9�4��N������b�w��GU�,�O�)h����C��{�Ϗ�I��aҧ�A	�)�m�6���s�̀D��r��jJ]���.�X��C���(���F(� {L�Ҩ��&��K%��U�&��5����wSm�
��%!˿�K���r<��}V8����%t}�r>�/:T�!9�E&��BW�m��׺�%m"Tʣ_:e�e��@}�o��ةL�?��d��uq|X�o���rKL7�,<eM8�
�v�[b�Y�K<�%�l�G���iٙ�ꏧ8�ßm�m1��0i�u�U����+�쓩�i�;I���AtxeƏ�˜�m1�@�4pq��.�6�&�m	G�;�1��.+'��Crh���l݈`�4��zg^n �. �4�X�҃騍$pWp���!8������)Rs(�ԭ��N��8�.�S E��^R��^�4��6']���C�b�%���֎��C��eU�/�@����/s�BL/�K�vH��gf�~�]�5����\���5�#�g{����u<��	�¡��޺ˌ��9�(`ɑf4$Ȯ���ͳ�o8��k��ze�=��S�v��
�s�t��3���� ����z�.��c�U���.�I���$`;�mcbc����Bިm��長���_}ˤ�:��BOY$N��<JSg�|{4@�f:b:^U���a�lZ��Q���40�-��k���1d"Ű���ai!1��d���{��oضf ��f
OqA�l�����`S����`�'O���bH��\��DH�	X��m��h�s��1|��p������(Ԡ8�}w�	W9�
�#L/{���Z.I�oj:O�����C�����@Nv/�?��5W��������t���޷���O:f��Z���S����:�����2���`F_$�!V�$� e�b躀qT���=�Vv��M�����.��T����Q��{U�<ۓC�@G��y�G�&s����sQ.6�������4��>�v;܂HDH���Ꝕ��x�l�ѡ@��*cV��%��h`����>r�HK��p�����w��b��t�̏!�f�
	?�!9���?n &'g���N�}��u����4��?��ޱ,7�����/��_ڬ��K'^ �2��q����t�XF�lSJ50$#�1�ɐPD��G܀��1l��g�-��� �.�~�4���Tw��P!�	UD��{�m��C�����#���-u�)/kUR^�M��w�`ku���v�'sE\��2u�gl��s#,�Rc�\�)��C�$���q��!��tM���S�x��R�z�:]�UH�/��$ ��{�)��f�щ-�=)�E[f\m�gRm(�0���۬��u>-�<�R�R?�!��;�0+���o��v3e顴���'J;�Vq�K���[�I3.r�-�H7[�$�;��x���A��dP3�@[{��QG�ߪbAE�+4����O�F�iZ�s��W�w��_[�b.���yXt	�Q�<lj��͈���AlY9v�7R�`�n�E��cAzF���"q1dQ=}RM����2(J�j_r���_}މt���D��X�ꕌ}�ޮ)z�V]��	VXF��m��Ob�ɳ���l��g��rg�����vg|b��=�)��G��R����/;V(��f��t6� �ݕU�I�R�_l|�xw�e�#�QeO�$&��Y�iG��a,H7XxOf�;�V�Ε�]�\�eZ�6�g^��8|�D!qџ�Z�KD��/���# ��-����GJuz��7C%{L�'�}'�Y�����0���^E�9���OMMc���і�ޱF��ZR�MN}B�����?ki�,���NH�$L$�;��/�zl���b�RX0��	�H��a;��xsSh#����ԣ=TE�|z60o�O���(@��d��O��B|���h	�fy���z�g�'H����iݒ�7\X�n�,�F���]:+�C�C�"�$Β�*A�0!ve��U�Y���b��6��P\ސP�A{��� �C�I[%�H��OV�f��t��@-	���>�%D��@�K�e�@I��2.��<̛�7�*%*�h<�7�Ȕ�	�tf��9��R�de�x���]l��%���zbg뽃_�T�m�iM6ܠt��UV�<`Y���g�n-n=�Bg@�++�[S�)�Z`p�&}nZ�!�i�D`G�}��z�5K4OY��TX��	_��D�H�BE䞲e؝5�!u*��5;u��V��~�0��γ�S�KI�w�8Vf*2sw�<����8TT���	������hz'�;�])�w���b"�w��U�Mv����[�Xd\�7%�f[j/wZ4�W�U��U#$W׶�܎��ɈV�m�v��d�Ps��罾W���>�~��[����v��gH_E�aP�\�xt�n�G�O�@?�R�;�7�X�F��4�/��<�C�}��v\5Z���x`u虩�2��}i(���<�A?�u�;ęћ��:����m-�YJF'����wb��)�8<b^~�L���̞^�q�o�l��֌��a��:�oe�ð F�g�|C�{��*��	� q�(1-~�=�~A�V����c�t�[��۾�7t�1?�ǑO��F�T�~h ��}�̞ت�ԯO�0����۰f�I��G''�=9���y�IR�P�������	�1�/�]Y�
�<V�6(uk�0�$ �ݕ�
(��3�����ͪ'�����ڦ��S�*X^�IdP=/H����ŰQ��ȥ}�i�.��_Av�du��B��T+����ك�ܥwE>���l�bL�t��Հ2�ʠ�(E>��J��L� ���b0�#���/��m�W��kc�F��;w�y xUb�J���dBv�^YxTv��s޺�Z!b��{��u��"I	9� џ��<�I��-�=����ٲ3�|�I����V�l��Z�{rh������'�M���.Y�u�sc���NgtD3�W��WrGצl\v�jE/��myr���	uY���D���b�N{t7��Z�8x_�@k]��4��"����>��n��+��ܓ��A��?:9��"TmH�c�Z��7%��7�t�}#�y�0�T��B�]e�FH�iM��"|�]F�ܙ�b�"l_��O�0�2zf���6�Ȭɤ�]0���}�$��|�܀��a�J�;�T$��e�	�P-�h��_�^�wL��O�9!�J��mG�<pW��i�K]�����|y Y��J����}�޼�R?(������t|�����S���
d��i��g|��5�W�>l�Kפ�l�[�.Wp H����H��u��"���tԅf�|���'e7ihOGĠ-�Կ����r�		o2�6��ф�!���u��O�[D�b�}j!�`����9C�/T*����v������nۓ��>��U�ZX���U5I�m.�A
�	���q��aFM�Vd�m���nX�Q��9Zn�E�O�kB�G�'g�7��	'Y�� ��z7*rݶ��^r���gb �g���@_�f}����E󬳳���?�TT�������ВQ��^�t��� y7Ug/� ��\�1����q���/�#/y��b5���+��?eI�AD�)WWeKi���ӯ�j�q7y�v�z���Ί:"^�.`	���,�U��˵"N�1�� q�9�Q�w�.%-V��X*k��]Ͻ��kw3�c�y ����ްlN�(�Y �B'`��[y?l�K��w-�j������kv|�Z1c�C�>���t��#�.���hn�<+��?�G�PXjT�y��0�����̌=��[cLY����\��������*���G`w�sJ��I_��VY��xºd�&$�)fm�H��$��K�=w�[[���k��Ổ!��Cq-��j�����{Io�#���v�E�z��5A��V�?�%����07Լ�d����`˳���[����\��e�O@߇^��q���I�V�̞���?��K��.�b����)������x���P���F�u}9l����(7�"iǾ�t���fR�(���/7Ť�4n�}���;�E8��#h3�E*�S�Y�~� �'��.���At6\�0��d.�W��X�.�L{ᰡy�[��7��Џ�������b��%l�L/��-:�1���-�X|J���t�f�U��ݱ��|��U��N�:A*�OgD/� 1��cUF�u<s�m]����`�;͈"/�P�sE�H��Մ�d���{�tb�@6[�kQ{���š��ד�zA�U��w���b,��6��W�E�T�WB�N�d����O��`>o4�`+���L~\�ƐV��3�SL���yj��W-*ScW���q���	B� ����:-�l�d�9!cI����9�2���JP1��SY�l��Ǳ՘&�b��v�C'W�[?��*�Bٟ�������F�uL �Pa�7�V304�I�h��K����Q/�-�OqV+�L��/<�V�3�wB�v��8�b���Y�23����\���PҲ�o|A�ޗU�;~+ L�㭿����'v�0|���S��B6l$�a���⳱����*%(e��;ϕ�܏{\6�y%��ժ��t�81�����k�z������&� ��;��aZ]'@�a�/I�S���J��:H]\W[�6om�CF���Q��X-�bk��E��|-�T\�s�q�)�2Tp.��B�{j�@UvWrH�|!u���Ĩ��%����KtK�ԓ��6:������<s ѩP�%?�D����|S^e:����,�l칢��ph�}��[j`f�;�H�lN���͑��[_l��v�&��q��+v�}}�A�����	6U�`��#�Ha��A���%��L�)�m^��k�t���yA5�g*�>��.1�ۅlRU�UM�������F$s��"���m�Ro�.����R�u������ϟ�<vAOe@N��?� P�sZE����	'y3;m J��aѨ �XU�����u�~��P��cm��Kz2o��#�Y>����{��厮���+�/@̵T��W]�#��*���-��'�t��:m"�KA8� x�P~E����ȩ�'R���I��Ď5U}�b��WmKM9�C���T0���ֶ�5�T��IݾT���=c׾�+Ql$�R�HuF���� �Z����>���.\�����5�"�/b���E1�+��O7�Dަo����=s�]�X�'��X�FG�%A&�q��Y�|��T�k�OV���̷�%F񹏾���|��)��B�k5��x@���N?/SI���[�`;�{�v�U�x4���n�ctHM�|�M���i)W��O�Z[2�Oz��%�Bk:���"�ƞv��P�"�����j͊��ӳ�?n��M�Q	��E-��AE��{d�2���63��{N��q���Pt}\ͣ&��,���d�E����r"���x���r�.=��Q��hN�%���W�2�zQ�`sl�E��� �ު'"�h�����c"���+�S����=���<W��Ąy�rC:>���kH�Dl#��_ƹgA��yF����#@���7v1���-��w$��f��= �ص(��Zߐ����V��̩�`�����@2�:�o��p8d�E
l^l��`�� �D����-Q�cd�+��栤S�ٷ,;"W�c$մ�`a��&�NS/U�6.�נ��
�&�*I޶�U�;<it�!L�'� ���}4��������g;�)e��xh��,�d����!M���H�o��+��/`����e�4;Q���Vt����u�E!}���|!_��h˺=h��0�Ӄ����(In��r����$��]؊x��6ѝD���pa�Jv�TWH��L}��9#j�(���Z�۽�h���d@�  �����VMhc�/s:��(���[�+��.���l�D�4|Y��S؈��GE�ﾌ;J�%�q3&�DB\j͟�^�<t����CϽ!t��:9>F$�7?b�M���+��K��j�]X�CQVX6�8��5KbgK���kV/Jk!�ܨ��(¶Ϟ��g���]�ֹ� 6�j-x����p�q�"�(�H���[�[���o��d���'vɑ�/��!ڇ����[�>��x(��*1<tǨ��bv���h�|q��g��*q�;��&�_��E��`��yvE����1ړ�+:/���y�����A���(��;���2��a_��Dro��'&H���
znk/�ˎ6�d�� �i+��ʹ�3V����k
��;�irQ�yL&f�-��K��u-�p����џh%!(��g�)�q�O��M������_�3���u�}����c�3�'��򞳗r)&�y���*�4�?&�׎�盂>�p�$�ݙ�;��)���'�(݁���tG>��,c�IM�[��!§���:�y��k��"B����:�˙�
�%�ᨇ>*��\��;��Ys�_e�(Z�,�3����;��k�"FH'�V4(��^ʜ��:���"����Dұ��ﯻ~a�?Ϥ�|���pG��/G��K�@��AH��Q���� ��pX�s�jwm����(ǡ�y��Y���vV�J3�;t�O7[u��oTw��>)�9�ܵG�u�?�����C,U��	��N��khR����S�S\��wm0H#��GM�j�όuV�OE�{9{��<���nq,y��+��L��HP��S��*��ngT�a�2�+i<�\���a���;�g1ɶeL<$N���e��P01�68槄���1�%{m�h�y��]Xw3X[��ڬ���u-�n��]ƕ Wu2�jԶ����֡=�gd�^.zɶ��_^�f�ߢl�@���cM�I�v}|�mby�'�S�ܒ;Z���fAp�;�h�|�~��Ul=�r����+�zmN��_��{����hY�orn~zp����6V��M���7�����<����{z�=ИcFst�	"��:����-e�����m�_s�5��;��/y��'�7@܌�M�]N�h�p�V��^�����'������.�Eg@P���й����E�����Sf���X�-��w����R�7ǋ?��d��˟���G�2��Xb>�y��Dڢ�f�g�U�4N�����=��IE�^��{,A�ҡJ_)�W��k�~�dfݓ�wؖ���#���I��0ތ�!���Z����!�����,��[޸ɲ�����%j�q7�Ǭh
g#XQ�̧��Pl��FI����K�:��~�3s��(+��֢;�_��?�=����\� rz�Wx<S��>��k�d�n�#<���,#���rq�����`�!;�m��3 ���\�nT�<9�P)�e�R5��@N~�.[�=�?��	�V-����"�eѸ�h#�����w�n�H�o�MJ���z���G#�������R������q����i�4�� =z�J}��Io��lw�� �4%Gz�'/��?�K"Y-浗����V��`i�U�(�"ٸ�>�bܻ�Y�w�A����[��D4��&:ƸY��b,
�iП�
:}i���w����eDݷԞ���
�hy��YTV�Ix\�F�g��3d_G�"�f:�C�n6���s	��c8��gZD%jԫ�ֽMJ�~��{h�U��ma��k\T��#���"6kh!�S�K�C������Ԓ3���l������B�-;�~5)���i�����b�O�\گt&ׅ������5B��o���[ii,�nJ�"��t��	�:����������������#'la�F�*.i�?�s�e���d;��3q�Veބ�,t� R�@!^*�.����7-M��ޭ�|�����8c��:��F5���Q��a��y"u>�G����yH�E�E l�Yl��j��Z4m�G �N�g	��B"=gr���}���������5:�4YW^�:,`�9[!7/���cp�!�ȇpG�f��Q+<x��n _��t��玊�[B� #j#�5��tz���9|w��b����X��]���B?�����c$������.�Әآ�N�l��e8�����$�����������-'��Ƃ�C@5&FQKK��7�0���(v(WAt\p���/~����0��f������� �LPA��kCx�i)[x=�"!�L�0�������	���D�E��8)��'�"�8�W8.f���.Y����%�����6?B�qPr�.������
�&�U�]����*;t����=I��OoKT� 7���u'���1
�]l��X]�¶�e�S�Y�h3D����x��[I�7:lѝ�����$c�}	������1TJ>����_>9梍�HA����[6��� a7;N��NWm~�tҷR�c��-lz�১(����7��(|�qq�fp�)��Q�L仍8�`��CsG�u^v�fstZ��F��ع�[L`����"�̤p�^��R����6���!�y�_E;+�3�y�� rA�"���&�Q,��T�&�ڸ������&?�<絜΃�p�
�)��'A�3[�Ψ�t�pHǶ_k�3�ރ����5����e�e�P�*�Z� ������z��˹�XzcK�iy��Q.����k�Я��~�F���坻�]�\�'�#�,��@�%�uひ�W,��:v�"�ؾ�hݕ�zt��@G��L�٣إ�f����2��>��(I��&�62��r���w{ ���pd�^��Ȅo���q)xS�j�2$����_X]9&�zmJ�ڨ�GC:`���^�'ZK����R҈w"jNNr�Ti����X��c�/!�,PWݭ�0\��U�N�G�7<���$��� u��F�r�d��D.]��=7��M�g{�4��w)�<O��v����\S1V�\ݾ4��a�2ù>�a��vD����ҩ+������Tf|@|h'w|����%{�����đ�Ea��������0=�r$6�YR��]��@��������HAR#���ܸ>"��l�.��v����gU`�\T��Z�!Mb9���;�I4Q�n/���0�e��s���!d79o�>��7�?7b63�%&KN��}�I`x��ݻDm�=^zż��(t��	@T�<xTI���6���	o�` ��@"���5��CZ��HY���]M��m��8��h��_~2쀗m~v@G����Ӓp���P��Lc��^#��/���c����\�Ն���s��.����&���au���"a6�
���|g��Or�S��M������c_��.X9L=,y~ ���������)���[S�a1H��$l��8�	�H��K?�/0�لF��G��k�~�>�Jf�B��e�۱�69�tP�Y$��,�U� �ܡ��-=p�.��rP��)1����so�͍�w�u�J*DhK��b] �i�L����': e�0�ԣKd�;�6Jɺ�r����w1׾�� ���C�Kۭ�BfC�
ӷ� �]��;��6I\د�i��
{K<hȥŞ��v'Wz8��������[�@�b�w�:$pf�(�Ix
�F��;�SX\N��%�iVN����8����=� ��N���C�p��raj�u�c�H�
�p����\�
c����c�Ú�u�7���,^8qnn���Fm��׿�W��ڀw���p�Z���;����8<O[�� �{̒Q �?c�C#��U��� ��l7@���Րcbk�2����)�U@����zcD���"�/�DXe�
�xY���-��Tƺn9n�)K5��VW�N;��$J"Q�.�ͯ!@C�Z�(��4���3CVK/o_B�uٷ{h^7�k)��p�ab�Ƨ$�<`�KJ��H�T�����ْE]	V��}dw�]4��R8cл^��1n�ڦ�U^nX6G
컀��t=�)���w����a2^9k��xцnTc�V�E ��r
�,!t_l�m�K��Mh�q����Q�UhJ��.��3m;W�|{eƙ�.{|�~%a7J$�fyZ&����=eb
�$��q%�k�P���>�]w��=����p��s��}N��ك="釔Z����8�\$J9*�"�M����q�Jf�`6�D�H��Y#�+,.w�dy{�ך�E���Y��~��(��}}Y�7�E���3��<�~��~��p�.z�B�ݏ�~��M1��<��;f'�#���D���v��р�q����1��L�Q��cH��7 �����U�6t\���Z*��jP�j�7��&��@%�=���8�I����k�J��0�Z���r��b)����)(��9��ڦ������ؽ�7D���Z��a@\\���J.d�i���~_�zrʄ��mJ� 2R�������6�D�*����T��u�a� ���(z*d0�"#6Po�%�#n�7��;����$��C��L!8��&8�-�e@�e���#����L���p���� � T�-�U�߶%���;i���c�S4>*fJ��_����;W���'UD��0�� L0Ç��~�O��2HV$���ó���t�f��h���/NAH�2e��7�
�Z��aOvQz��_�u��C�9���7�����P���i������.�J�5�_���ŏ�JG�@d@����]E��m�bcFS1��o���rz<Kf�D��XF2熾�:�c�K�t��/ǎ���;���E>s��r�)9����Qb~*3Y���w:Wm��'ʕM�V���:O���S���X�
_�v��Ѵ�.S��"F]B����K5�z��|I�w5��L<���a"����MK��b�~O,�l��ڑ����K��P�e�����)��(0f*��	S�]?���>Y�������o��hX���1�]�y��e�@f~��_"�ܪ���g��b%�����з�\�&Bc�����1�I��l���ދ�2y�®-)���x&b_Y9��	F�������/�l!pc:b\/L��h�(�E����I<	�^���a*��D���C �u����U��A��}��i�DOB��n����##��[R�~s)���gtk���`Ӳ �7�f7�\��	�N֋O%�ns����$9�D-���l,�b�H���A,�M��^ϊCX�[޻�T��`�Ea���4#���3<�sn	T�8@p]�,+����|�Ly,�w���K]j-�Q�4�y�}t.`gd���3���ڒR?Fr�I�.r�6nM71'mc�+�P�ΐ��^bu�^�A�%)ō �A�*B6-�?!EZ��3�>�p!�ҭE��Ro��n�G�$�G�ӹ|K��֋�R�k�fK��I���]�,
v��n*��9wA�����v��#���|������t<��tE�<�gqA�MC�#̈P��~�Kw�U4T�鮱
�����AK�7҄/���cw�:5��?8��P��'��Z/��.����������	�!���L����s��b�,t�L�K@��[�͚�`��l #S�fO!�I}��)��<qf��I�݄lZ�g?�����B�Ӧ��i�o��^)ܹ�j��XB�X�����ԙ�����+���k�e��_��C_�aC��@d��]�T�����B�h�A��80��h\,Bv������$��hEj ���0���w��ȮF����L���6-��n��'\E46wC���Qy��3Z�&q��0���U�&if�'�JR+"z��am.�){p�B�aR7�@&cհg1�e�R���}��?�#���@�V�)܈u��^�L� '��H��d�!���iԀ���x�.��!GMUR"AZ���>�Ƅ�G�f<���ao�bN��[���_?.^
�9];�{�q�;M�� �H)�X����~��(c�Q������2�h����LI�<j�#���-~}�v'1�PN���_3��D�g~��8�ػ��,������)Xlz��X����iL���;���ͅ�:v���̠��W�9�m�i9NO3��.8+TE���H�A pu�*���ZA�����lQ��{�)�@σ���>�Kݧ�%g,�D�~��ф������RO��n����P�y�SQ��Ͱ�?�{H;OR��,2-!jFb&7����a C�w ����?�5�Y��p|�o(�џ����LB>p�Hu{�'-��͏�hk��!�x��­\��� oZ=���p�0��N�5���,��c��Ѡ�+}������wnQ}��U7o�;���t��<�f�7w�?��J�!���l��|�97=P����!$���גuqd0Q�?`�V�DŖs��%���0�~���<����i�Ɛ$�ҍ9���+c�� ����� ���`pBZs)j ����y��:O_�;��f�&�H@9gq�5�K���%A͘"�߹r���ǰ���7�}}K�	�`����D�y�+?��3��?�$qQ�уƱ|��9�?n��Lu�,9H�M�#[�iG|xS�O�,2oUP1��<�=�g-�ZE�VaBb�9e���R�NI�(�o~9;y*Ⱥ�ꦤ�$�^�h�BO�<Ų�I��X:�m*=�N���&I*ݔ�ӣ�|1���E��1F�J^^���I��19�=��oZ�ʗ6h}b�Y��xn��>�þ�Gx��Ϛ2�.���h���3@-8"C����8�K��l:DB]��ј4�i�q�5i�n�S�Īt�qڑ3���C�l�Ա�n�������8c1�(D�KR�ا���V���0>�OrQ���&����+���'  ��������x�����"J�bE��Iht�
j2�&i�8H���|l���=��6�����+J�GV'��}�a�j��9�#�a
1l���E�;������&!��baz�O~�k.L��=�qD�˧�a���ѓ�
�I$�y=E�l��;_{�-�gX�Ѩͺ,Ş�$@��ko���^���X##���:G����a�F,��˫��C�D��
��[�8�;$j��j�G��	މ͞S�������@����90oRj������+[�x��H�)rs?���B��`�� �L���d�<_;')SHf&n?aqћQ�F1S+���Iֲ���5��2�}C~��v�JX;�f�$r�h�7��F/D9w�ˁ^-N���������Jk�YR"���&z7��7�����]��-�D����o�䊓��������eF|�c�0��خoK���J|;�|'c�rfDw�6#j�":��~\\\:~ۯ{C[�l�N�3�8�9%]�K�[�0'~!���!;��؉���_T-+�q�Up�C�s'��tQ��	�� lb��Dn��g[��auOV��w��-�Zތ
�{4�������v_�ʎ(k<�.W����JK���Ǥt�W  ��0q@��@��
�77f(�UIb��B���ka�X[I�W�1�M�m��i ;V����U�p�gm�j�R�>HW�uKI��=Y]P8��RH�X��E&H\���PܩQ[�H?�Մ&ל&����ë��)���j��t�t�a.P�t�ڙ��^E]o�����B&%`!�,\��D��n��ty�DmWa �"��"�!Gx��$��)�*�s�9��_�S�̪̿pr�Q4|A�q�Z������I�G��i8
��J� �-6Y��)�)��[�h,^��N7�"���*�؝m{�M"U�-ԡW �C�+����M^@��O%ީʾ�g���:\�>��4(c���p|�e�����,q�FtU]��j��`�QА����SGg��.�M����c�\A�S� �=Փ�=����jV���� [h�Azy&o'J��Pj��3=B��*����{%��(���"����V౲V����Vg�n�v�G�Y��HI`?J �H���S��g��N��a�'�lх���~��E/T�0��R:$榓��	}J ��U������x�t���� �ǝ��n�8քx��3:m)TXٯ���mND�:9I�~(G�4\\-e}�\�.c=�m��h �C�kT>�
��'�=�E�;��y]8��#)"��Kc�4H�z��6��x�0���"��<��6�V(qcO8���m��pg�J�&�#��L��)���7~D��
$+xjW�2N�U�"�K+xAL�nL��N�nJ�F!<��c�@4����B��;b�4���89^��g��l�d�;O��ۦO��� �Q���^rf��`�b`��Τu;�:K�jU�^T^�� ������8��YU�T�8��+��{=%J;�8�9��7���CI�EB�Q�q⩈L��i�)l8>E�~a=h��2�L\�n*�@��%����ӪЌpI�ۿ|��a%N$���/Ĝ�Ǩ)�J5����Лz(�|�hՐ,�m�Ww�Ȳg&�+
��i$�k��m0Ե������
Q��e=���?�Z��O�zP
���פ��a"�����I��nDK�Wd#�!Cˠ>����~^Q��ʺ6���շ$:ԩ,�C��A$���"O+�H�Ɉ���Uq1g\��a

s���~�H|��P��1�wjXE��]J�B������F���d�4�p��hu�p7�<G*%T�I�-`����B�'���Ԃl�c�#��㟉Kzh�y��+p�qWv�\��;p�6�����O��.�o\r� `.q��s�`/�˖ȹh�@���Ig�X��6��\xH�/q�cK��F+�~�K�{y�
��''
k|A��H7�����Xa��������ų�6h�狌A�ɵ�����.���,9X$��-���&��=�6�����D�'���v͞W/3��g���u�"s/�K���O�*�
:6�>:і'h��ѡ��}�*���kiq�N�ϭ��Y�V�����P,�ҎB���bW������=��)x��\&�����>���k�M[���,�t�b�s],Y���c�� "�i쫔�<�}�R�Wc�LN�qRU]9�a�Oc������8��c6�}���׀��\��
*�S����dL����o.�u�����A����5�π��ԫ�.E2���k�}ypF����ܐ�����,iΠ���@��H}����/�����b4*�������-�i�h�N�� t�rή�����`=�F�Rb��~��I��*tՋ�&y;�r#@yX\��i����̳:,6YU�B�nX`Zd2�3m��^�9����<W� _�R8 ����Փ�����Y��]HΗ��m�����a���	���+��IU>�� �7L�=]����d��������`�^�;�~�a9���p�af1��>��3����MZNtTȏDc�1�s���o
��6����'��-��o�w��x�{щ�����<��_�)�����P;�+Q�c��1$�氫�Tq��J�\6�`䌍g_rG����i� � �¢l���gp�J=��l�:e�ǚD^�Tv�,��I�kB*Nl��t�~e���%μ�[��
\B�����Ä\	i5�Sjp�o�����ji}�dbM��~j�]�Jx�"
�b��w��g[3����u�*x��k٘*�A)yj�����(��/T�b C.�2P��!4�R��b���}�=�`/#�O@=vy0�`(ּv���N@8�8�d����[}��s���
�����g��_@���6T�D X�y�t�f�e�M��+o1�Pb|�zb	��P��7����E��v(�$��9o���w�g��AH�R4�@� ����|YqϷz�7s�a�n��Պ{�ͭF~����DrT-��[�wQ�����ϰ�%`���bd�Y����4����-�'��uw����ͱ��aT�z�j-��: #���gdUY��Hڽ���F!qf��ދD}e�y�c�^T�8\�H��3�u��X&���}�1��lD�A�[2���}�*aZ�X*���%4�yÜ`g�����`��LH6�B~� �������I!�"U���Q��Z��:�:��� ���`̾�4������Y����4��Xט.�p����ܓ^WeR�P���1�o�pF����[}} 7�w����-q�<��r:�n֑�56��w&`�A�)��84�e�r�5>���o�>���mx�u�0u.u�?�-V�j
�8�'����?z�"�WFO���0�P2i�����O�E����fW`	*��@c{F��T|>^���;H��\��oP�h�t�a�De"k�xj�'}$��4��@B�N�|D�u��){l��x6c!��#��V ����y��X�{o���?C��.]�VƮ]���5a��֥JY�^��[tF#1��dN�a^��B����"�tG�a>������=@H8O����M��P��qVf�P:�ɬ��'���}�W]�͆dx2��Q{s5r���z�chK��~���f���,�V���wn�7��P��`�e�iH{�U,n3�X��m���6���fd]�#���i&�o�`�� �M��������4�6E�_������T2�0H������=�=>Hx}�2ᰵr����dC#/]X����t$.!+��k;���\���+�y�q�n����2� ��3��c��n�>&6�8�]Y��~L&��/=�'����yQ�=�ZX�ND��tffҺ��K0[8J6���;4I�?ܼj0�ܡ1B:���H�3��*B���x�~bs�K�Jϙ���8Y|��h쒉Į���C�/O�B�Wj�Q�D���C��CJ>��a纐VK�)��1������KՁ.'g=����9W�Uw�!� ]!�ݨ����^�|��͵ r�R�M^E\���b&����>��?z"l�4�ߴ���k�x+j������A��z^�)��I�32�ބ��s����,��#�a��[Kk=*��p�(����K�pT P�LZ������3���LR�!*�;p.]���'*G~y!ú�c�-)��4:hK4�QXd���������~�]��J���-綩<�E����ǆd��Cw�C)5y����M�ݹm~�����S�.#mzɳs���8A`���0 i\�cϞL�����_����55��lN�ҁ��0�� 8j���B�ʩ��Gڐ��L/Z<=�-D0uq�8]*Ml�����+ؗ�j�/��z^tqF��� ��Hʻ��Q��W�E>�k9.D�#r����ȳ��?��K�'�Aol�+���t/ʩ���&���	���x�}�TtS}���( �/����,ړ�z"so;�1���S �jf��)���k�)��7
�H4̥>F/}];	����
�$*�u�oi8���� 9�m�@�y^O�9�LDۡ�%�!x��$����~e�m6�A1	����I}�z*�9ay����D�77�V��ݬ\Яt���n�.%�M�,�
8!(�7�\0��X�l컥�&�!$?-�9_�Nڵ@��*-�޼��pԻ��k��~�q�"���:�h&�����2�T�Vp����P}��E�ߪ�ؤ�ŅN2�P���ߏ���@/���[��WU[�v�����rE� ��fG��7E���<^Ǔց+����r�KAï�9kA���򷕔��"��Ķ���u��x�+ߝ����"ZJ���\G���ha�ȸ����5�*�1uF��u'���'/pd�ש�v�j�_B{�@�	`x߷_�u�{�;y�f����F ;��=��\l=�jl�㘋s?����8�B`�9���b��~�s�:=T�F��]hHqw{������Cq���ʰ�	�S-Xy��PN��f0���%:-)��7�I��*`ڴ�|d�]1K��L��di\KLj��/`vsfQ1M5��[ܶ�r��f"��߀e��
����n�X�W�O'����Gg@J��#uҫ��F'�hz�M3�A�����
�0��P��*򮀝���@��?E�5+�K����FLb1�zw�+5ƣ납Fj���^�B�����~��j[s�M�Ȁ��(��4N�L�4�B�>�Q;����U�f����P ()pj�94�.g����ZX	�h��a�(�P+�y{Q����	9E��_�;���i�`�K"�|ǥP��g}�D+{�6bH~gL�D֣��g��ݱ��JD�=�u{3�e�ֶ����x�t�<�)J��HA��Z����y�?:��aNlA{�G��q������+�#"B���&������ �C6\rPCe�5P���}�^f��MKrg��5fI�eL���`��e���X�(H��-Sؼ��JG�B^&_3u�:E�����c����)h���^x�jͳ��K�U��B���J>�$���pi��[�-Ɣǫ&�b�Q����9�s$Ñ.������5��?e���@dE?��v��X)���x������{���p�B=�g�.�Be��*�%p����������6����ɿ�*�orL�7���Uکe�O_
��(h �e������	%)��,/Z���89�]���U����$�O�u�)�n��m1�(f����c��dZ�����3)y`B
P�h�`�f�oo)�J��١/��n�M	G9�q�����	�B�J���|����W륛��l?ە%��B���,"Vl�D��y�B$�:�.@\��xT3SG�����$�y"x<�������_�dR�D�s�ϗ`�~�9��K>Q�6VM	ˬ0��Px	N׸O���h��sK�;�K�B�m�B��TN�r{�h��IT[:ūu�vj��Q#O��s��{z{��X�x�V^��}t�=+C�_��}�c�Ƃ٬|i�:-6���0i��S�*���U�C邶���?_�r�#s��g+�9t�*�<��vz�e�d��]���a {}tE�����h�E��͙�o�վ%�����J&GS{���?ew �>k�az6-q>Dd�E�v2B�`�_�Qu�#�]��0���=Ӈ�D��fknG8 6[�*�\U����0�⢻��S�P؁\���O����x1)�G�ra�kϔ�������޷��~�2/���Z�0��A�4�>J��DP��b�sRr~��������Nm)� (:�YF�b+���!{(gS�� �GS���N$Z؏
o��{��A��ڷ��N��k|Qr3"\��r�^�}�:�\h�LV��/v�Ӹ�`���8LK��!�O���7y�A��?j����-!�&�cb��}h"92>������E�m���ȇ��<G�Ș\=���neumtQz���l�mk�Ns=c�t�)Ӄ�3�
x��A�wP����� 10���ykk�c/�/��Ӕ��j����H��� 9���I�S�����{ڹ���[E����_{|q?���7����cp�l��X��H�\��g!�I,��慾'!��'���ډi���3�x�}�v'4�	��@{�B�g��r=�S _�.���X��әp a�[<4t��t<.��F|	����j�X��oi���<��0�V솹q�'��m�O�B=�-;�U��F��ɉ;�}��KrΑ:U~	|� ��8T~�u�ͻ�q�D���_+ L��tC:��f�k(5J=��6�0�u<����W?�/w:#sR��Ul�kX;Z�Q��D�w+�"�� �a�t�m�h�,���]
�b��o}U�'��=�!��M¶�+�. �_�� }��i7s��;�6q���8c�'L�N�F�W�H�?h�sI��l:]ա]�0��ܱ Sȋk�+tf</�:��[��ښ���|�Y�Pڶ���S=���Sm$
6�'p��fOU�;�gd2ݥ�lk�A����x'D�R6���
�"/4-���=&��,� � �S�Dp��>� q.�R��t%M�G�"�!Wݸv0�����xP��H�`<���1Я�Zx�>��.R��I$���Ϟ�	<D�j��br��$�i�����U�+l�#g���)h������Dj|d����F�XB=�b򱄍QItAf���.�`��ҫ����v���Y�>����M���Ӕ��R c>Z'�i�g�؋.�+�=��1UX'�д:�E�Q�ܛ�Ö́�x�{�/L��t8��.�3��������"U9�	�s�?�4u���\k��+��7�;�j<�d%� ��LP���rw�;��	1꓈O�5����
e�����_�mas:��dЖ�W	�@�.ao��p��t#���f)�`��^�Y,�ɠC����*Z�Q�"����D��vm3�ϿNq���R�[�F_T�ˡY��"{�ڷ� ��e�D+IMI��HU��)Ԁ�����v�(P{mf<����~*Ƣ['Xn���2{'�D%�:5ԏ1�R����P���qH�ͯ��_Z�+.c�҉�����oH��͝�`��4��U|�@�-$�y�����Pơ�ڱp\z�Z�<��|��oP�T��]B�U�����p�9?����|�y]j��35��� *P�p���v-�ք�
=l]�o�`�dT�{JO���s�0���;�<U_^�����{#/'���2�\���7}/�f�*��M�b:�U�"�\Έ��]��p(��Iޣ��nI�l�����z"C��)0]xw3g���;S���%C�*�'�k8J�%�Ip
��F����m=�x!�ʬ�rN?��֊���u�sTm����j�~hq��=��@AY��I0?�S�\i��>w�ݘ��Wh/Y)��1�S����e�C�j���o��+/N�'�eI���w ��^.�I^o����eڵ7� ���[��!�u%7D'd�:|`O1	�)<%?��g_�Z5r4�6�ބ��_85y>����Y��S.�R��i�����x�������m�I�BY]S�0l/W_�H�L�d2B'`�(H��d"�i�1�~e��%f}~�-��+3���zJHW��(��C��g�,��� �|Y�.�v�h@h� ��$�c_�h�ۇ�	�^�_���_������U ��9u��^~h���ت��E���t�S�\�`y:&����`���<�k��`'Ұ�nf��񟓂���*����=ñ,"4�\�\��;�u&����@����7� =�5�♈p�/.�ʎ�%Q�~�G3����xp� ;�"�����XU��1|_��T�}yǔ;�G�[�0�!��}S��|�/.���;
�+p�\%j'J�|6<���\�%��t���k�m�g8�kˎ�e�]��-�-����;���e�d�
Oˈ�c����nn�!�?��	�L�:���E�:j ~^�tsݞg��o�#�O�\t���u���H��!{!�p0����}ʩU�R����3]�
�4o�l��XI􋆖2t�!���O~m�[�/��s���5r�2��i�*�V������i�b�6�{��{��m̻�̓��w�n��=T�����SQ7��kd�6�������S��<��K�Z�̓f�@@*8
+���m3����v��,7�+��q��qX���"S
c�ܟ�� �̇�FZrux/���]�2)�
���)M�~��U�c������8��g���	tbizPW��B���N��A&<��� �R�i���Z���2�z��I"���8�B����Z��.�zq�؍�C�iƐW�b������*_,(���)Y|�,�@�8��r垞�z�x�#Ӡ5� ո��m��x�㦷7�����y{G+YC^��)E0E�Ӄ�cxA�=���H�{p3��~j��Ϡ�i��B�Ȁ��
f�71@'�$�.Z�L�?�y/�qY��oz�qF��Y���^�L����6��� �<�����ż@�%�κ���J�.X,&����s���I�+�
���Iѣ���n �ik�{r��o#�u���O�❿�|*oOi������8�{P���!��:pǒ�����}3��ۯ��3>ٙ��T���p���Z�h-Sf,�g����ґ����$�v�u⹗ ҋ����W����]�=ja£Cc��r�]�?�t�@�V�
�ͿU��60�w������6?���iYw�Q����O��j�?ޒ���BӨ=�G<&�9��Ҿ������.��&�_Z�mm�#]Y����|�n�0����N۟�@���ۢ���;��?屹��"T�dFfK��=_�D�� ���q�F��6Ǌ��`x�KIj����K0�3���ug�	"}�A�k���9TrNz����]��5��r���Oz/g�(w�p_��U�uZŶ=u)�/��cVJ}k�	U�����é���Jk�a��'�(����jm}D����*�~�_��9=���6�k�w��o,ũ{D�i�Ϫ��6'�[H�y�c,�>�'���g�(�=�g��ζ��== @)�c͎�S�3����Fo�T�O���TH�t�5�)'��������L ��|�bG��T�5�9���5��s�*��X#�gx�fVy�\8������C�0�"�@���/�:�l3���ܤa�'^�fq��J��]A����V�Q۹o��8x.�z��z��7��'� ��7����*  �%�U&���+z�����q�&����
}@yy2�[.��[��ӛ�%z�i�S�ɯZ*9�f-T�'��ď��7t�!r�ri#�2��F��?����Ap݌*�6��v�yk=�{n��2ʳ��dʂ���/����9,0�9��D)CL�u�W��q������u��L�`�~�{%��(c�`ns]�C�ꔯht���Z�E�����39����m��f98�}j���2����M�<:�H3��e�A�4�G��I�ֳR�gO%m�51��g͚ձ+����K�Vhm�b*��0�s��&��n�(��ewQ�vt��.����$���V��A������.2������x�t2ZR�1�T���r�����pO5�f�$�<�PRp�_�8dl���Y(��M�W�[�B�â=���sU7U A�l�I"�����҄,�<�	$����'�mB�X~K�gb��,�\,�k�3Ɏ���S�	�Z�w�ѭ�h)5ݔ�~�^�br�Kh���x�����&%{���.������R��mT4YQo#\���������0SV(>r���ǺJ�M��O��ډ	_�VK5�$����]�3ƻ:ئN�^���F��F�:�N{��lg�J����[���o�<�S����H�u���I�.ć�c}٣�B>bn ��3�؆�FM}�����ￊw6�n�v���?!E�E�!$�]����8��v�Ef��nm̆v��m�%��i��L��������k]z3�n^��_����#�*�y���l�\�r�<��s�'� ��d&pTG���A	�1ԸP s �"g>�[:Ȼ��zJn�a�t�>@|Ɛ��P{��ic��H.�Y�6��}n`��"]e���v�B)F�g:�;?	V �6�N8���RM-<�T� o�uR"G��o� �5�貈j<�ƕq����9W�`'�$&S���T���gf��Eɉ(�R�G�~������N�h�-�W��O%�����<�&v�0A���J�Օ<�1s��96J.1��o�خ K�ġJ�io$~������+���͡�������u5]�d��������˨1��DB�k�비##W��������wT���Ff"P�Yn���^��L�kۓ�[j�+�6�b�5�̀����p�<p�ř��b��1.���k%�d��Ѥ�a��GDCi8=�,����������x/㑧��X^�	��2J�S�ךl��v��\$�)��ת�>|y�Z&��mN���{Mze��B�b�Ǳ�>�?"��� :1L�ư�]u��@:L�@�j[�x�q	F�<K�M��t3\�Z9�g� }�3|��ǔF�'�I\o�Ll4�b�+��5;��˘�2��1L�4�M�uɵ_e�"��]+�:D�~]���v��8*#�&-�C�$m{�Bk1*�>]e�)+/x9���>�`0��P�[Fn�ے�$C�c�͍s��G�Kz��,o��$���K����;�����ܝk4}x,>{Ŗ�@]�%���I&+O�sv�����h��6��S��@�
������8z-�ǟ�l���yO��{��8f��/�)���F��~k:ʨ�@���^�_lZ���aX����L�[7�wrq�63��a3XE��g��6�lߒ�2/�9֮j�w���WOUY�������0��w��� 4f��̠8����o1q2�sG�
vV����>[oD�N�`���0��$@��q(�y�/N�X7�:�4^ŕond�f�-�A�(�Y�������mz=����Ɗ�&�H8qI!�����ϭ׾3g�s�0Ae�L��$�!�|3�Ew�%$b��SB��r-H!�c�i��h�u����D;)��qi�B䛫-g��X"=��y�E�NQ	��g�A�?g���^�,-ϕ�&c��B{���Ծ��/|>�CVS�t�-BaO��fU]��g��&����F�?,�T��w����{މD���EŞ ^�:[�»x�kAaa'���p��/%�.l�]��F�E�Õ�9���%��ȟ'���U���hg�/�ǱVpN�ml��#���,�`L�V�ij�7�ޒ���/Jz̺~𛶎�W,�rB�3�'�+�]�T�Geg�b8hD֙��5��2�$
d�a?0��u�q^p^�=k3��?d� �6���Z���@����MI"�Ҧ��p����yoT�2|������VJ���Ǎ�f�܀>�\5t�Mjr��{O-
Jgq�y�CY������Ks�`�kE�pBrn4'�Иt>�6���ri����r؊ڭFK�V�\�ߜ�|�@�zT�2�4�ei^���v�œh7r�? ��nr۩N�_M��h�p.{�\F	Q��뱂O��L�&ŋp���l�#]<ɴ'���L�W��:���(��?����|G�	����n��l���N���^���SC�X��^�a_����� �8�m�S�l��'��FGF3}����T5��c�^D���K0|e�@��
;̵?S!$�C7a�X}`s�cr\�Z�p�c�i^&uꍠٶx�@��p��g��A�=�C�^�m��u��ȝ���I"�_�Cp�����S N���6��P֍��3r��<&�����㑠w0,�'YS��:�D¶�&��M!BT��6wUĥE3 BH�o��!+�2�Ϲ��N�Y�k:Q:zm���RNӧc���(V��ħ��z�1҈�9��/��Ꭿ�x;:-_C�&�FЭ��_�t-d�Dy��$�YZ�h(�b�jL��>��t]�n}x��, ��Nsٮ��R�)�1���Ɖ�!�_�9�ŵ$ژ 9���N�b	b���X��D>A��w��A���R9�~�c�Ŝ�ۄr~�����X�e��?��T"p@�����&x�v���2�c%��!uP^x�J,|��R� Ә���R�)�s��+��!r��%Y�]��&�fѝ�.���l�7���+�3+r*�$���N�>D#Zv5;�3~���cg&)p';t�y�)��e�iJ�V����&��W�"����l��P%�J���mͯ��!�1l`+���̈́3]Y����a�OYa��;�m "y��gIXm�gHZ��5q
1Ǆ/�o�[���b�b��~�2ZAi�	,�UU� ض�a*zA/E�~j'�IFС]�Ðͮ`)���}��Gw�J��?T�5�K�k�W���s�o�KL���m��CF��յe��RЎ+0Z?H6���W��QcJ�g�b�_�*��6�>*ɰ�������A���xe8��f	��<5���+ǂ	kTX5��
6#��w�_\�0'��M�{0U{�X�V�C���
��a��V�<{9̀���Z���=��ID����n�$O�gSX�@?lP��,nw�N;����N�{�g�Sg>�IO�/���|D+[6��oEw�[I���A���l���eJI���-�w6��ah��+�m���t�<������dW����4��}��ɹ ̞8r79�m�]85�����2���b�nJ��Ώ��P8��Xޡ�YC�;��_&�z4��v+�HEq_X���һq� ��=��bQ�����/��w�^2M�������>�3���O�������k���Ap��.b؋�-����Yjt_H��x��?Wڴ�j^*,p?�Cq ��M��P�U�B��	�e�`�9��m|���)����p��l���#Q���!��G�2Q�|�?<	� ���YA͈կ^@[������S_&YVg�tB���T�;���p�`��<`^�a|��D�]�/��I��ˇ �J�cb�&��D'v�(����b�;P���(��í�Y���sά�2ҟ#SK�/�Ni����mT ���C(<��e$�|r^$4�ń��W\:q_�2f�70���뙮��f<M�=)������u?���}��!rν�����NS��Ԗ:��5n��W�j�`�}�}��gLUO�T��<A54S�Ҕ�qF`xR	P�bZW���q�ɧg�gR� o9KiB��-�T&�I�uN6й����q���;%<'�n��B-V>)�m���l�Q��P�;P��S����� �MPW��T�s�a�E����a�{�0�'[q"��N���T��ϲ�@7q�l�;����{y�xJ+�u��sw�C���	t���g3&���Z������/_0��s�ڇ35����Q�!��_�P�[i�Ϋ�P�<���V�S��ܖ���z���x�P��nD�anא�E��yX���>-�r��*��\�C�%
��.��O.����Tj}˵p΀jRM/W�	����g�E K�Iuڊ�ͪ��,C���!�x=+���ҫ)�e�6Bѓ�@����ul��ಎ)��䌗��&�WT�,��y�&'29�f�CV��e}`��ۤM!C֮��c�D��SwC�@�U>O��Xf<��P�.�W���V\�B/ �f�t)/�a� �U_~��J�}^bd�Z���1��GyJ3z�#U�M�SJ��;�
.�>��e���N�G����+Np�n}��ԝ0�5��ˈBD�-��9��_����p���Æ��M�źK�D��Kԛ�t��H���chޕ��UBGF��E[4�Z/,�e�j����M�ʺ�� ��DW�U
:�)��$��]�T,�ʎ.���MH��]
�*J�Eup��购���r��Z�XX�Qqvg=��177.���Q�lΟ�猝�3� G�J�� ���|���z�FTe~��܋x4�4���`23���%*� /Y��q�[az��hx��l��gC��&Zn?�l�$X��Pc"a�b��gp��������qځz�jB�,����������L��V�)��8��P�ɕM͙��7	�WKQJs���$��
%5��|��Ln��H�M5:�e�����[K�"�3�C����W�}QBH!&l����%�g�z�����|8��(�v��}�����s�\��Agoi�x�
�l��?;]FM:-5�4�N�����̀ھ��Q�<-3>:�z�w�NR�l��'\��e
���-i���rJ��X�E�s��yJQc=���c=@�P��0�:��xW@�XC�J�e������x�����\-j����,X��)dG;A�\H�����y�b��	������/V�J�>+����^Kn���������]������I���N#��-{�!C=O���i�"�
�q�t[6xQv�<uS��6Hn^[�T<?=ž�[~���z�n�j�e#��x�����>�/8	(8�fۨL_����z�I�?�2T
7qJ3�#
��Ϟ�C��t��c˯�k��C��Aq2�u�rv�0=YUf�
e�O~nKl���|	�MQ�1�'�B���1R8<>���6���^����e�Df�^�cE�Jm\��Ҭ��bm>�oW�p�Ol�7g�(�c�QS�jT�}dsJ�h�N�Oy��,���]|O&W���&�3��"�j �+_��}ÞZ?��2�!������/��)O�9[�N���S��:��2�[���7(��pG�&W�K2uHx�i�2��my�o6h1��B��m�a�����@Ū%ɸu���fà3~Pr�Q��ˈ�a��݇�����h8����ח�2�
���wǨ���4G���H+t�
3�;n}PW�Aq�7z�G @zW���7���	�Խ/�H|f'�t��|�r�������ս	5p�Hl��u6��"��n�
 ��p=ߛ�����C.�A�o6�o鲺_pM	�B���9Bi��ϸ�r�_��!oe�jW෦��	�\���}G"�ӺU������e��L��LV�Xh86�ׂ�4�ч�{���f�Fs���/���n�fZ.ZC'� �G�댁�d[��:�۟�����R<d�79��I.h�~	OtAX�f	?�L\�r3�z!���d�����	�%����i�a�l��[���4�tctH�'8wk;}��������j��*��� ���'!o�U�K��S����+��u�٬�����z~	���E[U��k���ծ��xBƓ�֨�{�"���a��05�����>遾.V�o�SH���%q _?�A�+�ݕ�¯`�2[V�.��H��Te���e�ޛ�����(S+@�����Ec0�VGJ�qD��]���V}yIO|@�М1t0�����*w��V�+bhOp��[��j G�6�1���� j�Q�G;��?�-/�"I��.���9A�3��&���N�H���4���<�T7H��+��V�tO�ϐ�g�1+zRԦ�����JC)R�+���4�A6T'�z���ʻf�F=�VîpIp
�3�?�����f?�
�J_��xY(|��C����rIPK��(�"Nf������X�:��9V.�� 8���OI���|o�&=y���dɖ���fF��Ȁ��
+y�]����E��f/��ح�}L;�s�kt��"���wT�Z4�2Xc��Pb�)�?�Z�ƛ-���`�s�ʽ�D���ѝ���Q�&.į�Y�T���6 �x����ώ��4�GVi\����?g�w���j�� ,�/~��X��>G7�S*N{�7,�������zx`�����x2��M��s*�z���Y7����ֱz�?�ZC�M[��	�m�/�()�M�y�!+)���sh��.���ظ}[yk�L�n��pU��9��#`e���83�t��C*VY�h�Y�5�NC��ٳI�����b�m��Y~�އz��P�_�5C����<G�L܃��w��U��AfC�W*�]���,����+����71L��A�#���<������!���~Ç\��i�>/�,Vc��*���Hs��^^>�P�B�B���"h�w1�<���w��bE�Z�'�3^ț�����~� HcHj-�&f*Z��Ow7&A�����8�-�IO�bҡ9�ۛ�r����-�Y� ��m��J��(���_��ǌ-Ę$�eCs�3��8^*�[���3��=��xWi�f�����[Bs���Ֆ�����l�YEh�&474�Kn7��#h����p�᱘�$2��
覾 1ٕ��E��I��0FKTa��
YPֺ�6��q�Ѕ�2� WiB��~�\��w���wa�03K�񳘙A���Jɭ���	�ʗq��>aP������v��
��~VDN'�T�����z���é�X���*5���]%H�HS����r�&�\��u˿�3�V�GQm'����o�	vϮ�f�6|́H]CZ��k��17%�&[��@%;˦�!���`��Q>0J��/ۧ�b���}e�\ǜ4yoY6=�Bb_��R�)>V��獶�Ma��UUL����6o�Bc⍏��X�糉��͟1��?4�ĭ���K3����Q9�e�*�'"�:���R���=4`y0�;ܖ�����H?`-��+��"N
�f!�]��Kj�T��dgIՃy����y�N�ԘO�Eg���N ��g���r���]��Ƙ��.�s�Z�$R���"R	;�_�,���1o3ָ|/p��,�پ?���n"�hjlDW�<��ڤwp��"��d\�Oe����M��\/�嘬g�5�	�k�j� �Y����3N�!C֖=������s?F�>����oL��53�8H�0�~�����ܥK	�Hq*��P�2���9�p>�R���xVۯo�)Гf�D��}7+]u�w�~˯�h�JBo�/O���le���i0	������u�-t-��Z=��:��~}�bs 
(C>�A	f�`�vܥ�{�{�vlS3z�R�&H�3��IND$9���ލvG�s�.���D[�]��.@SnJ�Iqjf��29"R����Eڷ���c�fp����w1�i@�����d䡳�}�2>.�@�?�"�x�F��j������$�q����Sec���v�<}��tqe;d}1� �b�/S;1(CKʞ�>p���rL��7*2L�����W�5=!���.�����ɲkH��w_����� D��$��T\ʢ��#r%~��2%��,�y�KV^��
�[/��{�x�*���*��+͠��M�!���� 2r��H�8�6������Tf�L��!9��1H2�sy:%I$������P-�Y��gV��6<�P���M�ƶ�:��R�'8�=���"@�a���i����f(]�|0��@/^W�9�K���Q(��q$�.���<�O<4RX���/��z��캐�����<G�������aJ7�چ��(��:?�vp���M�&�,j��Q�P/��l^:�pǘ�$;zP�N��}+>�UD)����?��]���7M5��23z�G��:�KHUb�o�y����ȩاv狫�ju�Λ+���qU���l<6�	��sR!��tUQK�w}��
��	R����� �d
K�<��.��l7Y��2��Y�Ӭp%�r��fC]�w*�Wj�O�ȧ�J�^`�)$r3��I�Z��Ҿ��iկ��O�`��ُ��s�i�Cv��z;���+# ��?\m5j� �p�h'=��U_�p-��~G�� ~�|�$��9W��W5l<1�+wt.s2D�7�x�=c�p�v�1](�tGI�=�"BS�r��>��r3��j�R���"�$��˚�r��Xcɲ��|<NoDH��w��t�D76�FIN��.��F=m��-��lR�&�pG���C#^�Y4 ���&ؒԙAU|8O��S3��?�x�*�E;C$v�0BF�<������i����TF*l�J>F�D�<`k��I%u�$/�$흳��v�+ͣd�n�ge����������r�[rˎJz�D��r�{����Ӟ����%C�r����-��3X���{�ӿ� )?_�6��F��b�t"^�ޥ!XP��6ʱ�<08O�դw�̒?!y$���u�_� 9�EYv�u]������+�%�(T�Va�z��}��n]$6����_��:���)՝N����{�h�.�i��Bq�D��\ꇸ}�O��*�%��"���a�o�g�#zw�Е�W��	���S��˖�?�����z��A���7�8LS�Tf�ers;��	���&4D�s��x��!�8���E�/aQG�g��)��Jqk��u���9R%��m�hpR`�'�9��9��7��B���Tf����I�3 �F,[}�ڐ!�[��[�M�d�\�ꇘ����Mn@S� ��u��"��]�U����M}��Wv���_���$�,�I�#ڐ ��*B���J�'�5��I6*Ӵ�8��Mi7�#�k���JUf��sj\�*1����ȐJS �n#�f�Պ��HC��c��xو~��x���&��^��<ꢚ����9�)�W.���	���>��]���"H�ڂ� '�c^~`S���p�~2�0� Ѽ+���n����l���%���G�|U�p{!�̟��`���a���Q�ی��
�aWx�X��EAw��$����RI�Q��Q�l����N�XN>���K�^{����?ʖTd�� �fR�fv_�j�۫�}�V[����y��}]������.e��,P3<�	��}FH���̤�p�(�]�L�W��8.��|G_�[Yn���<��F��O���d�Z������d�!�GL�k�L�m�#Y�c��=;kz���Hn6���Ҡ��=��ʁh�b@Ĥ�ޠp�-�me�rǺ�;�=~-0'V(���~��#���Ef{��� ��/ǦJ��(]Ѓ�Ί�r�a�9S���(���W;�ę��+��T�����Ѳ9,���ҩ9g��!2%���SN/ES9�M�^�����Kr�:*&g�$ F����R�W~$X$X�����?��CA�
��&魚?��!`�e�I�[�=�_��僻C��;�����J{u��𿞢��ea���\�zqNJ��;�����A[�6�Ht>�3B��ǉ���?X����p���9�����UޞxkTb�d����'�}lg0:�0'!�;�ӳ�-�S��h�"70�k�,�KO��� x�9���7�~�lvC Zd�n+����� ؈
���'DQ<��;���SU�]G�td3K�� yR�n���SNՂ�q���kL���XZ3�|�<��R���!w���� ��Ll��	N�z>�_��r#0�9(L'�A!��ޞ'� M7ɘ�l�ŕE�F	Jrк�-�y��t�u���?�45�V7��{��S=��Я ����,Av�VT�hR'��f4�L��iG����Q�MX{�=1�!��iFn0d��F3�if�Y��+���/�}�-��0 ���Vp���t����#�Pe�~��_��BdZ��®�a�:"�w�	!b�|h��mdiPe5hCh�KF����dy*=���p/[y���
��-ֺs��v���>П&�&ʺ���K3�\3'@E2�r����"]�Fh\��N@����<�D�^�װ��q�%JT�Qqa�Z���}!7���aǤ�o�Ռ� �+g�G��Gn��d��8jm��#�������~*��U��]4�-9��]�I�B*
�|d�����؆?�$�E�_�u�-`���	񖧆�m �����3����T�m������I:�%�h���<l�y�d��a�{�[���r)#�~ A��R=�-�"i��n�eJV�jm;��*�q�Ҡ��4۹Oъ
�%Hg:p���IJ�>�cb�ԥ��	�EG���**�C�L����S��d�0 L`�1!��s�nǏ{���@}��.�ǫ\=�6�\A&�tUQ%�u��#�[	���˞����S{ [�0�(�wܛ=���5�&vm��#���o�����5�����"�l��^6��0��	��a��ϓ�Тҭ��,��l7ID]�3���lUUTk�z��VSpt����i�xI,a�g�*�A6)��	���%a�ʩ�l�w�	�{nEbx�����{�ZV��G�$IlL�K�ƼJ�t7c��4�d��ڊm�>j�-S��h%�Z��Y���,���XU3s*N=���KL��λ��NL��C�:��6��b%��cc*�����(��D�R�m������ukJ�ʋ[�+�O�G%��r����N�2��8.q�z�4��&�Jq��2GHw&u-��թ���qW��mQ�e��v�}�����)�{���9���}�Ϙ$H�wsX�$���:x���C¯|d]K�M7� < �Gep��%J i���ZWF���XeCɪ�/�XǏ�R��Ma���-�o��fl�n�S:Sz�oPv%O`'�a���D/(���U�+X���N�i�ߨ�,��X=��� ]���E��]��@�,s��-Ny�c�>M{��s#j*W�[�k�'+5Ĵ��G�)�	J: ѯ�����Pk��Ȱ"�ZTu{��n@l'��̀��n���*l�Q�.N��3��]���u�����N������/U�L����E����1�%N�Q�
�ꚜ7��������?G�O��/��۵��~�w� I���bBD�����8�z*�[? Kx�{v��6�9�>��o'�P�������F<�T��+Ti>�Z^@�Oj�Q�ptז（u�Ɉ�| ��UkC���N7M K�*����iZ���_Q��RI?�?���:�دw�b��z`r���ޯXTeu%�#p%���0�3x��Й�N��%�lc�hŌ��B(��ѯ	q�(fzkK�'d��!2ď,��Ӳ 	�!��l0�*H���b<�t�Lq^�����_��on���՛��S�Ӧ�.��o��e�_g��<S��3<Ln�Jg�#�)�`��S��ؕ��?�^M��R�z:^�Gs�O��UL���c��r_p����}qj�a��ƀ�T�Z��I��3�y+ƒkF���r���oh�
�ϸӻU�3�3���Ѽx��~yB����AjZhV��Jd�9t�әZ�(a�0�U�v��<�Oa�V8qH$�P-Z��zV�[X3�l�9pU�A�\�ܝ=���-�ӧ��c'�2�uH樳��\�x����Śf�9'hE3�Q4�l���{Nu�X:�ަ�GpԞlҽfp�u�k�q�T�Uh>�{9n�-tR�f?��!�i���`����'��"+�0����%�[�d�c�9}����fP�O��	����,�{k(k|�wV�VD>E��-nPa:o�+�z���$ľe��37�:2Ƕ'�	�N=��J������s�I�o� ��@Vx�d��f)v�����{��sSg��Fl\?p� ��@'��S��ݽ�YY��|�b��^=E�d͡|�]��xfm���o�.�@l`5����G$�	��X� 
K_%�#F���>0ٹi	!��he˂���l�pV+ǅz��2�����H&y��4�w�'�_�/��M��K�[q�G/���@[�(]t�W���980�
�ʠ�%���K.t�̄���>N_l�����k����y`1�t��@RU;Z~��.[���m���Jh�a�X� ��O��=�����V g.�������Z�:ޟ!=��H^"�1=j�k�+6m�4�Q�Γ�2����v)cC&������aV�0np$C� �D�Z��alb�.4`E��p}=(�6��߿���]�q(��斴�p�I'*m��:l��lў��M��I"z���o��B��Y�K[��1eQ���i��o��cO[[븚�Û�4������䴰t�L��/�c�j¯e'��r��'����-��vL栘��n����t����6��m��&)�?��ǟ<L:Np{�" X?�"5E�{��C^M/���B�J�v7+
�@�r��f�1��ƣ��Zl����z�6�� |�q:��5a�� �'|�tcU72F"�(lS�|Eʜ�6
�0����9&? >�7 #�M����8Ȫ6�T��Yb^��<��%�n����1U_Ģ��
ן|5"0��s����AP���m}�G��
4���8ބft�@4�j+��h�2T�����>� ���������O�'���0�"0,����U3@i���B�"~KW;��#1��T�/?A.N��8'Nj����F=�Ϫfm��{"LV�	<�fQǺ(8	{ 	�\�Q�}b����8���]�sU�ɤGP��pY�ך�r��V|,q!)�U+�gc I�
�.��s��h� �fx����-���3���l�CG��땭��4�׺I��8��o��\�y�6�9P\6�*����Q�Mpl&��N���P�q	 �}Iҭ3�u�~l��{ze��k�I�����#��T=o�~�^U��J7�iT.�%�[hs�����Ǘ�>������rw7�B���lE���P��q,7nY��{_αC��������q�+�2GqM�S�f����Ў�lb��/��+���t�K�.EE�q}�?a����fo��<m��l���5m9B+���+\w&�4�O��-��5�����`f��Z�����e)ܭ���\+��~�������20*$��|#,�<���؆.��r���dÊi��m�'��S��װ�r�yMV/�	���$1�� ���l�&���� ��﫬b�+0z�:A�ۘJ�������V���L����4k���~خ�B���-��u��KA�c\�qf�Q�n^c�A7�FON�*�1`C,�2�0��1]������Γ��k(IG^<%�좝��ש�,���L���F2d��B��)cp�PP�b�Cm�B�ޓ�?Eځ�u�{��eDd�{�2�G�v똩{?o@Hr�S�4=�/�ű -����h������~H�Y
��K���D���������w=�I1 ØPs�Nǋ`Y$m��������=�)����!6��@�`�Z6���g�(����+�ds��V��J9��et�fH屻Ő&̅e��P����>ǚ�����i_nZ	�Bh��<�T�4�Up�kۭ�6L�R��e����ƅWs��[�w���2�[�
UF�}zH`�#ź��uML�H��땪��.�.�T�L�B13'2T��S�
���
����G�)�n��Ga׫R�:�a�a9k ��;�S!j���^l�Roa��4�:^�E^V<��>T�?�#4ib�z�4}���Lg���I��h� ߗ��y��[؈g^�]a����2��@t�&{��o��m��pi�������<��5�3�K�e�0Y',8�yQ\`Q��IrX-r�0FVH��)����+�lI
�5������������[���e���V�W��ύH�_���o��.�x����OupG�#|�cO�S��/�٤T��{����a�L�4�ɻJ��Vg�e�
0[� HN]��%�,W�PORRL��M����ku�q��Si�FwњIO�gL���\�X�d�ux�F�몖h�AF�&��O0���i�w�
q���c0�D��Ou����:/�>2����@�f�uJ��e���a���`h�e��w���?��pT,��03g������>�6��ؑ8l��C����1/\])�B~�+�x���~IhV/`"̼ h�5?�]W ��+&��ra�NW�%{�ws@ ��}ΌoO8��9�(ݏ�)<��{��v�&K-�D�Uż�!�ʃƞ�ij� 
`�`�Z�W@Ի�ƛw��TH��B�k+ !��>�l�Qw�#�;_C�:{�;�T�*#ɉA��ǣD"�5��l,k�Vj�)��R�B"���}+85項��a��8����n�I�g�9ܧ�#�Ր���v_l�[Q���� ?%���'B�F?�����xh�j<k��aP��Y�\�i|�W�t_��3���i�=QY���X��Ӝ��솵�r����iʶ�� �X<�_h%U`kLY�� �M��

�Ģ��V�-�N&�#Iz���۾����d��6���l�m���g�2*T��� A��<�uDٿmX>�JIm��� >�	{2�x ��:��t�]8�N�$���u�Χv]�2�62���8R^�҉�$�]�H��Y�<��<xz�)]vO��[�ԯA=��%X���ʓqRdo9fYoEJ�	B,�?�W���E0l�t���g�G{�>�K���T�4����h۩��V@Kn��5)�b��l����ɸ}%~�2�`,��e	з/�k��������1�mc��L������n~�))�2�笚�>Ho��B%�<�;���$t�b��b��unH�	��WL,)����6��g*-"}?x�LpеY��Y^��?5�
�A�0���|r�f�� �+�J���(fj�����q�c]��[�ٻ�������\��g�2��VHD�,��]�{agfƾw�	mUP<5q�by��$v�u̡���CNe$W����E�"N�C`Oq�.L�_�gO��$$Tͅ�.�$��t��j��H�N�Q4�cn}�F�`�t�w(H�^;�r�9�f�[N,Z�tq'�~�dT��Aʱ�D��4c�RX|D�0z��bƬ������[�9�� B<E�������g�1,�㈒���"�5|h(U�ؠhŗ���B޴�]�v��6���Lc{�s�d��2����"�[ם-k �<Cn�\�SV@�j>q��Q�����-�Cc�(gJޔ�+USOi��~A�9�"��Bx��4����Ѧ,U�:��N���͹�� %��������6��!3wj��3X��!|���y��`�*��:�J��k�*܎���)F� �A�
�e~	x��Cp����щ�z�F�@*�x��\�!yi~���8��(�-31yr�c��,Mj�e��=��_�A|q-+@PSY���M-��������0����S&Si�VZ��4E�Z�y��m�D5/����m���e����M��M���G2��Г�!�\z8r�����*�m�.�?HS��R�"�w(��f�l���G��K�M�U��}h�ܗ�:�5!��L�vJ�#o;7A9RM�d�	��7"]���V�?~���yQC�F	y~}�ub��ϒ�"��Bi�flfS9n0^��/2V�*7s`��[ʑ�{}�5�L�k�<8ڶ����e"Ѹ��p(;dTv-Ľ�[Գ�IҚOSr���i$��b0U�%T*�4� ��42p��ӀM���Lb��y~�^rR�����3T_��
��K�o�bi�Q�h��m�!o�Jo�O�M�C�%�Q9P��aX_9
GU���M��_
����������QT�e�DnW��5>�����.��f��G(�)��\�G�+R���<�@+������=<J�8�-j�|�oM �V�1m�\3����_��gaH�~�5��u����κM��%!��S� �*%���;���q�ō%�y~� ���UYX�s&��[o;["��j}p�� �K�mz��z���Cy����;�/���Q�1T(��!�;��M�ih���a��RiAMc��Y���^��bu�b�6�&�}��1ݶ�^���06�0\l�����f��U~�)v'���6�zrb�xW@J��>�d���ڊ���r���;�Ġ�5����F�
�t2C[3�v�d�W��ǳ�A.�6������z8����]چ�N�!=�Gk�^��
Q�2�N#\�������R�d@��@�taq�����-��O�U߻�=�⋹?������c�����E/���-��ΐ�]T-(�Q��E� ]�p�ɡ�;�[�3�}Zs�9�uD/�+e�]�O����c{�l$ 	��JVG�XS�zځ��׳�ø��Ig�EUj��B@8,R������I���Tw_B�o�t�`�#�SH�Gڄ'%�7��$���S&�-���f"l{d�/B�Z�"�b@D��){3_��Pm6�(j}=cD��f��	�q���?�*��4N����|*��W�ؒ�*-��Kk@W�s(�l2�'6@�@��z�����'ߟP�g����o��R2� 'v�v�Z^{��u������U\ϲ���Is�������.yI�N[�P%�GH&�p�"^~ ���-t�0/����g%�	}m�*���^���F!=9�����=�K��;�����⎋����8zp@`W�\9Ge����8ڼ<�Y0,>0HeZ�`Ze�Ϋ����A,�jl<@���W�Q���_-�_~�֛/����Z�nmP�]eu�,s��)^M3(R�����a�7�w0)
��==n���Ȇ���C׀���_�e��=�V1��21u8�=�r����b6��aC\~�1[��1�C��j��rЪJ����ؙ𰶼����3�2%���Bh3�v\*6�Њ������\�=�Up�h��j/�T�S1��lW�@#
�B�<�B��̰�%g��z��)H�e���q�w4 ^6�t�!	���!?�_�0)��0��ö�vJ�AJ�J�)˯�2�B�1RU<��&{,���b�v������)9�����G��ޠ�]*`r�ˉ�,ދ������t0�-�b"�������(�'yg+ԋ��`��^�ۓ�s:��2mL�B�XI@	���k��
��p�U��.e�3#�&n�Q|�k#s�eX@s��ӆ�X��&����j��6�7�2��vz�Q�|Q�_�L��9��| QuY�?'��ZZ�z`����F<�ͷ�z���"�J7�$�Ԋ��O�|��ޘS��P��ce-޻D�ih,5��^/�aɛ�+�Ѵ�l�<�]D�P�9�����w���l=��c;��c�$�SHyr3��'kP<�VOv���ф����m��������H"KE�F��O9<��7�n1���j�<� F������*:c>Ns��B����h�H�����݊����x)�e7�v�3��M�~����l�6�AA //e�&��3q����ٔ�(��I��sU[��(^ޯ�f(c�&�/v�*���,~�җ�4xe����(ٲ�k��f��>�Ɩ$�!Sky�Itco���QC�������ؾJO=�7I�q+����d���!��H^���7���k�+��r#f����&cGx鳤�k_v�)�`�d%eF��7(߈�"3�`�69{%/�����~@�E"p�����L$O�K/-u������5�����'�ŗ9@�$��sӲs|O�ҳ�4Sܔ-g�w`��ޒ�$V��>uf��:u�9�R���3l/ 4�J�/�����b^~��tEYy�\�j���h͜�ͨ�8>�R������d�*��_g����*Q��`���"?�v��.[��1���J��Ѝ߷��N�'��k. ���K^_0� �'�"�
r+���4�����lЧF��홻���f(���͊Z>���풠ƫBʏ�#�x�hM�;�Ny��Ị �XTS*_�hQ��â.��p��Pz�(on����� �Ac��� 6�����1��;�+?��M[,&Fo����B4P o0�o�X�8�(�m�Hk�����8�Zd���Bx���sQ��? �ӃVݘ�cW�Q�S��T�9�L�@�<,��Sjk�"�us��؝-k�K�U���)~A9���C"xDI�f5�C}Ѡu��[<׷�ʁξ��6�;���t��ۿG+�&Y����mG<�H��S����d�y����և����JsIfZ�z��J�T)/�V��J��x���(T,O�W��7Ö��K���҅��-�Cp��諢�:x��K���<U�u�X�Q�A�\5L}�� b��y9�j};&�%Ҵ�(������o�D����`I��Css��㓜��5���9A~5X*9wJ�{e�F�n�6��;���W��j�u>�Ջ�$j�$�"�6W�.�$�9]�I����U&Q�~�l:g�ZB�:� -��yD��c���1��P,^b�i����|D[���*k8�o=g�2�D��W�M��UH�Bؔ}�p�p��)2�0F����O�>Υ�4�^���oJ
[[�!�'2�!��l;�,]��qW��
�l�y-k�ӏϛv�י�"wώ�{[���MSؘQ��Gj?_�\�+�Cy��&DC~η��3!��I>��=kݎ>�>��A�x3����å��w)^źW斍7�d4�>�g�<
�1�E8���,�~]�o&G�Ha�	���C�8��:0<�Z�田v���UО��|��5�ǘ�l�8��z��u@NΑ
��x�ShJ���d�;M��<�	�:��P�@)�Y�vd�1���J;�6�~o�Ƃ�#��O�-)�<xM6ڔR��������'X;����'��l��l�f yi%�����0�oW� �a��\]���  �*�#+ҁ_��i�]���\vƛlQA��)K�A�+�Ӧ�E�#�f]>5��F��L�f���$q�N�Aq��3O�u���6&�#M�77!�#N��ЛB��t��Z�A�yA�7��sS��<��(��#k���� ɼ����XH5 I�0e�y�%���F�������-�a�;����S<�H�a�#u<�)����Ѣ5wH8�c��iU=
yl<��ф3:��hHE>��SZ��v_��^�;��>*��ɏ��o�1�^����&a�a��zS�n#6wn��������h��M���H���K��n�v"�6(���I$~ه�@�kv*��J�O흁��O��T��߂M��rWE*�ţ(��[3p(�0�j�(���ѝ.{�����`ӯ �*~��U�����=��xZ���HP��q�bf�g���S@�}�%�/���}���l�Pep�Ď�%�},���,���6>��_	6�F�AS5�R��;1J�r�=�������*��4�N�	��-s�¯����֗fY"	x0���f�"�xe�ZfߩL�A����[p���N��f.4����&s0�IaB͌�	��2ڸ�&������zk���ՏS�����X�N�DM3]�6�K>6K�	H��OU��B�r�4;�%�p���G ���M����,g�@�3@�[Kq}vc���/���-`�bP��y�g�V�GL�}R[��lH�(8R�X�����]��*������.1�({(�情�[�'��_��s�߭9qV��w(�"���������J�o~�}lV���7�I�*��w���&p��G&�ޥ�{���es{p�*�UJ!^ ��0B���AE�-�+��*P��/w�������E�]$z<n��O�6P`�C�z����wc�v��ͺ�ꋣ�<:=^��j���l�x�#L���9Z�83�oG'����l�FȠ��դ.5'(~�I���.+jG���^s�t�}��.�' L����,dHH�Ý��w)�F{VuUC%'f*}���n����>�a��k��$T��\���=0�7_�Q�<ռ2^�%vm�e}��]��3�r_�p��q_~,v�TD���.W��������e#������PE�/;�ا��ow�]Lm0�6f1H ���U���"��e����d]��A�(�����=	.�p���i$��Id�q��X�1K��:*�yTz U�hv�d!�̻�@�M�ɩ��0� �hW��J��w�BȞ��(n��A���%�'����'���X㹄v��-@R��ba߄!�6>��������RG�A��+ʢy�W7������M!Vm�ybM��ׁ��zfx�vk���)-� v�B�`Z04C+
���v�m(�7�����Z���}"� �\�8�F$���zV�* ��f�;�!��Iت��S!�n��;]1�)ņ�e����\�W�L	�����Xt�w�R�qA�Ч��Q�>hjٔtڹ!�7w�'`�wX�e8���oD�Z�zCK묓�?Z(.�\+�"��;��Al��(4H�k���.��U�HM3�4���4=��)��Y�$�w\|�`P�\
,�c�G(�T��,-|���y�����)s�ml�cK�lC�!3�EhZ�d"J1×`׎L��^%A�)�d7!l"�������w�����{ۉIS��;����6__��/jq�j���5����9<Sf����yBȮ�5�ͪN7�KÃe���Na|u��` d_9 G�H�����=�Sa��8�2�%T�O;m��:JqJ��a��ҳ��=�G�-ݲ3���y�Ӛ���"7%�o:C��7fxӆՉ�(U`t��J}��*˻�oq���,v�_�[�B����xo��Yz����o@�{�q� n*�����Y�9.�3�i[�J,��Y��E�|�+J�t��ê��0P��~.�k�͗��j��q���xbǓ�?����t[{�H{h�����S��m�B쮴�l��@��� �����0Z�FPp�Y_��*����V�:j����u��3.�k����5�qS*V�Z�=��0F;_�/P�Q>�$8Iነ<�Q��&�$㩙I�ό�0*�mP`<����!�.̐��;םn�� tx��<�oޮQ ���ۀ+�Wt�)�"�nY��i|<̝u�?�w�LdY�eh�m)�Q���Z�ǅp6�E�D�m$-�(A�`���ʗ�Hдځ�GPU��Z~�Ѥ�i�8���	=�R ��0hQ��(�?i��	��mĻ�6FrG��O�?��r�6�&�Z�B�bx�t�ɩl`�\�{l:��b��R5�s�Qx�?� �p�4b�vNa��л�����~�Თt�C+<
�"�LI1�`7uk"�C��5�f��rM�%�-�3��)����BO�݋܁;@�ygO���7��{Ӽj�. -pX�r��R�9��S�����-n��wC��gJ�v����rIk!N��_�0���-��iС�>�Ӝ�v��9�L~d"/;��;��^�*P�`V0~��� Z~�F����B`뎺�;V�qJre��'����v>q�k�^i��s	�s"?E�׼=���Ųܘ��
��� g����g�v ��De����9�� X�J�2uʕ�*���umu��]ߊ�v8=p���ES���-��~_���y�l��7h�����tA��B<J�Û��ю�uF��|��H�.�q|Ĩ eW������fs����˚y�=��ݞ�ռ�iSvޭ�?�B~@Z�,��X�l�@�&��b*N�E�ϻ$��������R�
����䅺��\�;M�p�_���VC�8á缻�2����л�k�:bkL��ݠ��h�'84���^�4��X��*u�n�����ұqĢ�� ^&��K�˝<la���ϐ�u�}蓙������Z��%�%��3O���#dڑ���*�rqRUlPy'��K:�a� ��HX�ʾ�#�qE�����4EG����O6H��[[Kn���/�
ǜv�xTŕ?�մ6.CW�P誻H��Tw �L���ďk�`���7M�}=���ZX��L�:���q��=�/��D��QWn$�����"a�3�آ��M��
`*q�S�.��N�o5)���&���H��)� � ¿c}�*l2+����)�<Z���� �pt�4v4�ٻ�U[6�.(6:J�l����`=@��հ�� l'�%X?D4c? *��4G/��2P�]��>W�BR�ӌ�9�Sbr����& oQ-oo~3�`Zj���\ �~+2�����gAji��U'6���<�e���b%�Jq�~�Ӡ�7����eiVN���HT�Xa/N��Yϖ`�$P/���Q)�FC*P�q�O�It9GcGZw�CȨ}>��J���vt�=��|�2��1��]F_<Aʽt�ù
x?vn���B0$Nϒ'�2=FXU[+�����z�"'[�R�3��l��������Wׇ{U>X�xM
�p�+�H��0���mP��N��X����R���������3��d;��?���|�&?�S��k��R�^kA3��4�҄�|h�G&��i�eľ�j��:�9{��Ԑ���YH�Y1�.?+��Ç�{�Lǭ��R��(<9r��ۇ�Xo]�/��X-�+b�d�]��6n��%�&c�f���Q�)����Yef,՟�z@�\�*̘�+��J�1������sY�a.Y��֬ʒG#/�M�p�;'��&�H8ѱ~��r<0��*pi�;��[FX��]��}�����nm7`iP�`%k�i�Y���$'�(�+�N�����eU&�����][G�ʃ��q�̃�/^���ʬca���j�l�Cd¡
�>j�Gȧ��Zg�8R%�x�P EՃ �����k	Ka(x������v���0rPa�%G6�#��s�)Al;�[�W�u� ��.�w�.���K�O�:""����Ō(�;�X8T�4c�A�<��3�m���ӳ�10ي7lr�4n!�%�qܭ�ͪ�¥/G(d=4��Q,�q���J��s�a�k;=����K�'����
9_��=nńl`�>�������gI8
6� SV�����9�N�P��f��~�w�}��1R��χ���K֟�F-R4�gTS=�qU(��{�A|Sg��Gm~������B�ĭ:�c��,g�,�������F��t�5���m#*�Ը��(O<҆Y=q#��f���s���Ntv�R��}�
��K�Іq���'�݆�&�\��9���}A٤�v� ��E�\.�:��vd�%L������EF����Ї6�;?���
(��4)���>����E�A.&6Citũ''���[K	D)4����]�x�/��*@�?=�֝�k�̮3���vPk���_D1�R�Z��8����͈�4i����V��е~p*�F���`�����v�W��3�l��r>*��5f�&�$�J�@��>�<4�jY����
l�f'��,� ��ێ5�	��e�)����P�Ķx̮�d�/b��SN0�R�/���?E����!ɼi���������5�M��'�����"_�q�ƹ�U��(K�� 	ǁ�ɠ���ٖ���T�g���1X�걇I<L��+�W�z��)��>Gd�k�|�m�G���1]%@��4{�?��{�(��m�U@<�Mu�<�wT�#��ݵ�H3��� r�;h*~����U��֔Y��Q4��.�z�	��e>n�ڞ��g�P�1f�/�o�j늾p}�xN<��s�>
 Ľ���TT>�9��zjs��{S���9UB���Ο�`�`�@��ǌY��/v�����W��|v0�wh`�D�F���1��J� ��ݭ��X!����q�o+-F-�m�w�֌�Q^�ٖ�N0'~�b�L�H�f�=�!sI�z/���-n����i}�Rj]�b}f��p�Y����e��N�(f��]S{�T���@���l�,$ �Xk���Q�Q�O���s�[�E�Q�5�L�TZA�%��+[m�$s��t�d�w,b�T�%�j�C��Kڜ�x�(Y~����rRe
�(ϛì�Z-��}��4�V��$7��&�c�A:`F��^�A�E�-!a�Un����O�d����'ǫ=|��,W`��(1ѡ�)q��.Cp
�y�wܪ�H�����W\����4�Ut!��7�~�Θ:�F�� %U��	Q��q�̓��vO�z1
��yq�����/�bLNM�E�>(���Jv=�Sm@,9����Nt��/ݩ�7=�ػ�Hol�-?��> s��=���ONY{�/�@��`;�6~���:���j��NЃ]oޡ"�z󰩔i�P��fX���:�ߪ7 ��
���1Pu[#���u,v��e��h�V{l�DWr�u�-��3�|�q%}oQtͶ��ݖ��Ƭ�G �C�e"�>��98�a�U��?aex�#�IJ���d=�ywǾ���,��:0�ě�]�ԑ��z��1�Q��s�����{r�旇-J������o34r�)��c�b�&����n�K��➴|�?����<��*�B��iF�~-���h׃��q,�Q��)�`��x��YV�)7�5yU����WQ�k��W���Aג�/��	�{��ՙ�<!/r�	�u`�E$,���܀O0+#؁�Y��&u��o���MWā��l�@��(ʕe�2r�"1������qZ�$�1=�}z�6�lű6�����,Q#Ċ��@����Λ+��(<ޜ��8>ӽ,V�o;ڗ�9���v������`-�L�� ����2�C��o�r}��@�"���ܹ5��Іs�@A�^�Ԭ,�^(wf}1<]_j�&g��Hޢ��>�����X����哀i&�� �����3_W	)�h'�R#n,�{�8����S�#F �_+��Y���Dz:G��m}�]0�K�@E$�܏��uyZ�[p�Oy�=���P���CB�3�_�������z̍��y$���r���c_l09��q�K��9r"�p;;�H	Q^���,��Mo�=8��X@�gm\1\_����E�Z��3�����'YE4a4W�Ѥ����X���v�P�[���� ń#��o����P]�rZPW��#T������A'8�ٰ����"�А�����v�L���;>�˖�,0NCIb+
X�m�}�I��gf�n̐�����N��j�������DJSJ5��7���[|=u�9}m&u^���r��
�+����bHׁx).�$�A����ǫ�3��i~`���&�	7ٍ}�[���5��6�`�O�]���_z�3?���-�u�(8}�V<�cuf��?��C��;�����%��FG�Q~���6P�\��פx~,���4,�v��Vv�����BDC�� �;zk]:U(B�u������>��Ʃ��xZ�m'�Ԝ����ťm�tև�O�S�A!`ڀ�WȢ9ѸM�t�qi���k���D>x�F\�L�|~A�핑�ُ>���� ��}�7{�{������V��ҨaAMW��+�DH�����	�!z�D��}#��mӓ8�`��t-��-��=�T�rS�������BCe[^�q��X[a/�؟��Z+\(��օ(�"��ł�Ҷ<�z�0�ɽs���&Z���n��� N�~�7pn��!���xXE5�Vِ��_,�����7����m=��ƭ�ku��)M�|SB��H4rړ�#[�e�͜�ca�M����J��&�ip<^�L���Mt�M*Cp��7�w���T�R�AM��H�'Qk�H*w����d�&���_��C�\&�D�=!�����h#�n��P\�����ѣ.%t坛9��8�4�_��8�;=�r
N1���> З�d!��S}3�j]$6��a�jb�\������"�PE�֥b(yl�,ݖL4��:rY=8�Ѹ��P4�� _/�M�k�])������>~�oz�<5�5�=W鵒ԏpĴ��szm?��� �L�B�<̬@���S\?
X�a��s�Bs���y�zC�\t�Cl��\}[�H���v�s�p7x#�-d����S��3[.%�8~��u%[��|���������]�ۄ<�Jsq�ڜ4��$�n�Y�*W\0��حi�Q��NŮ��^�
sK�����)N�v�ԕ���pb�Df/�6�����oF�&��JmV����B���#T�U��OK�f�W*;�rH������}�M7�Σ����P�?+uAo[xͿ�k��zWmvońB��wj�ȅO���\�1��G�����`��_Ɣ���Y��嶒��$�jB�lؼ>:B;��e�p�X�i�������y���*��'pgp5��M���������m��NZ�G�� ���6���t�Tݙ�z#�Q�j����ڞᰃ�3a�ՉZ�`W]��{�&]&c���a�9�u�'I�:au�|���"�pT�F���W��'I��5fn�c�`�ggLP��ci�~G��HVH�a��X��,*�'�+�]��L[§(����v��]<S"��0�8�+��RIy�6��:���!i�0�cg&=��2*��tݢ�_;b�5���;�����0���js� B?̈́Uj��ϜQ	<�o��Pj��.苈6z!��>�,��Z7��}��3Wg�'��2ζϔ����^#.D%Ub�+��L����#�`�%��W��������P'��y��������@�$��C���̼��u�ȥ@�V�g�e�?�|��s�K��~i=�vB<J���ᒂ��1p���d]m��9|�^�0�n�;y�ZӾ0P퐹Մ���>�ѿ[���n�;7�U�����(���,`���3y`��aZ��T���m"����q" �G�O_5L�Q�W��P�Op'�>QZ:) ��
� KYlg5�1���W��K/�Z���f� (!st+�j̡��Hn5��
�̥��U��Ȃ�ם8��$�}���`��_�I�A ��QKs�U�GK���.���s_�����\���Z�!�=��(I�&,�OX��	���L9��B訰�.F�xN�@b9<����zzW5q��m4.۾?�~˩E�{ӷP��&~�Y>����ˁ8���v�X3����%��ł�T��D��f=����D'�b�m':�C~��-�$�f O��--�HJ��|�U�I�c9hO~$�q\Ť[M���ݴ-	�g�5Q�'%"��)zs .�$C5�{��1���2&?�1��$s���(o��M�(�wJRA�;�C��v.ф����4GhRlM��E�dBy���K��������xJD$�pU���̐ƙ��Q������=���6��'�J4���c�$��M͜�gc}���o'�`�u�@m�O���%n���5g[i%��k�~�T;/L�����HIV�Ȳ�tB��6���P�'���D�������DB1�����ju(�H<P�o�y��0����$Ҕ�n�
��2:�ډA� m��IC�ۋ�R��eo�f-1�����;}S��j�E ��D_�]��v5/����sR�X�d��4[r5H�������\hj�25�@�I�1�?��w�1끮i8���4�F_خ������xK�O�cz���+Ci�X�4����a�j����T��a�Gw��7��'�5�'�2�@�4�`M�%���QP�A�`8gF�Hಆ��tZ�J���/����E���TQC0P��3�	EW�5�$J�s���}`����}Su[�Awͫprs
k
���4nK�ip����kƄ%�u��`�Hޅ
����Hգxk�ZŤ(8I��|��!>R+��,E�VP-��Q�(�� kV',A��4mL/���a�ܷ�\*� ��Ъ��Yr_�C�(���y��Y�&>1dQ���s{�\�O�컸lV4��7fs=��{�2`�*�.ʨ��+P���{`n��o(�"rH���$���!��-�͑����eė�"�?}4:&��V�5��a�c��)!bf�<k
M=2ic���gߎ_`&��>��O�,�]��Z�詥�iZ)�Ĉ�m0u�ǔ6��R���2�Mo�c�u4�+?3�)ymZv�k�ͺ������ŝNM����� h|�z{ߦAP/�Y���u�pan��rT�Y}zq�>���4�-���>�4I�;���;ٷNtϹ1����jQ%Ȩ���NE=�Z�a���^�y��{�u�J�Y��d=6[O�Y��w���]<Z���x&1� �c��y������
^֑���)Y�Q�n�f�W����Ő�G�6�H��j߽���WF� U,1�y
�0�����~n$IPu&�3=p���^���������]dn���ᥬ����TXQ�c����cti蕵��R+� �!�i�{/ւ�o�ϋ��Z?I�5����ϊ�h�כ�ca��Б=��xci��"�8�7��7v�3��O�m
1��js�o���l/n~f,�ƜUa! ��g�yI���ڇ���3����M�[;(P��%:G�W��q������iڧ̅�:�M|�=T�0��	�6A��k(P��4�ު;6�h��{�5(´���ȿ!���Rޫ�. ��|��20sݻ>:.�ܡ�:=�����o�y=F�z���ep����ܮ����վ�7��>��@W�����p�)�61�B7yփ�(e���ǖ��?��µ�}�i½�aQ��a�	�`�I;�g��+�;'��y5�ǝt_���6�u�W��]���c)^��xS�9PF:c˴!l�|��l.�O���g�e �8���C�[@! ݄3'�W$P�O�־Ȑ����G��QH�>vjCa1 d���I��!'2ݷdB��?��a��Fiܝs�f�(V����_Tdɡ l��@?2a�\�u66���ڏ)M������?l]��\~j�A�6H	�1i�&�`��R����|s�i/h)�iw����@����˘�]s��s2(��o�@�
L��6�!��Ds,'*�1(��?9�/y�~WBHB5�1�̥z��F�VE�F���w`B$Ѹ9�>���e2)i��K�i� ���P�B8��v�RD�n#aӥ��d�%�B�P@~U	mRAʨ�M��� >���nw����`��C����`�§������k���z�b�	�Y�l�U�A"�Ǐ2�C<��G��
� ��/~h{���Rg�+t�蠉D]a�~)�Ma`\��e�%RZ��>7P��8ѿA�;F�&���;��$����R�ڑ6�}�ږ;f9��Ģ���v�P_���W�Coom*~ē�46pU��g��������廰}j�3�%� �}�@(#�ϝ$���6��^a�dm^�X�Cj+�:L�1x�3@��ؔ:�秸����~�㭲��v|�\ ��S@�!��q���7�۔8H虓s����g��*��V
��� ub����¹��J�.�l+��>��ʇ�
ӱ8Y������s0�_{ɗ�X�z�3�t�bb�����k����g�b��k����:���W��v�Cxxyp���@�>���P+>��;�*���ǘ/���Wmg�̾`635y[��#5֊]�d�
j��������ݖ�?�mx�jw� ������g��
��O��R̘v���߁|���q��M������?�+L�5.�H��_5����Q�d%�Ǩ�g�e{j���ks�]}|�U�k����:C ��+�5�V��1��@~�{��ƻ��z�S!����RA��k�R�������O�`;�@�����P���?\oS��(f9k���O�8�ռ:���~�"��q�懸�4�Հ�X����4O�,{8d��u-0ĕ���Y���w�1řS����h���t��<lt%��q"ch��"zQ`�� �o5S�c��ɤ�d�b�S�7.L,�\R���F���IJ�n�����b�W٘�(f�4��`+������ꢂ>�w�"o΋H̧@�(������W=]눊����������<'|8��2�eP�H�����u��
O�V����
��|�C�a�9�"��={����?��'�ْ8m'�L<�~{!s���Ok��	.Cn�Z�Cc��5�b���,��?ϡ8�C����Y'q�c�Iv!�l4�S�W���LG�8�A� [V��L��G�� %5h�*(x-�~2���/��>+Z�ܥ|"q�	c^���=G�}H6T�̑��;�2*����UQ�T<΂�4��:�-�8��y�um(�x�T�����BQ� o�&��H�xT���,��E����݃g�"��ݒ��eU������0�<!g����It�=d�}Z�W��8�	�VOVx�qlH&�)�Wr΄�jr���e�']Rq�E���ȃ�*�⏑P_81ʥl�@o�b��l�~�@K�����S�>L�G:�_9u�ArxҨFK찍���[q��4�e%*�gO3'��$B\^� �?=�����H���T^���>_6e���^�")-��Z��4#d�;9��m��)�<�EL机�l!5Q��֑��o�a�l�q{58xk��T=�tDd
sڸn�i�����}�8.o�L�="�GXG�T�2˜�,�F6#FU�
���U������*#��x�(F�v"JK��by��W#�Ѭ�h̷��~�p��g'dfP;-�*N!�L
b~��;���SK���K��U��H�!A�����w�:��ÙƂ\�U>�{���hr�L� �CKpi23�����rP�����4;�NV������"�V�vi"�g4�TO��0�V�XJfJ��CJ�,���u�Z�v�z�_��,��.�lq��6*��,˱J�_�`��ɻ$�R/n�/ت�.)i�S`����Q2��.;}���ρ�Yn9A�yC𤔛7�!$�ȹ��=Q�֏F;sU$&�0�,	�m�a����r�4��yt�zOZ��nh�y��I��;)��9�mˤ+�t�QTO�3�d���-F�uS���`{_d�l��t�$%���F����:�nϮ�f�a�<Ut�d����q��6Y)�v��s����ʎ�g��\�c{�8Q�2*�$!�.irm��3�7��;���!�M��̯K�����dj,���Ӗ�錯���˴p�[4~����ǟq�w��j�,� �W���y2X���'<q/*F�T-cO��ˀj�IР~��,�q<���Լ���]`���CV��V"�m��Z������4��X2�>�5sm��Xq��W8\(���xF<Y{!���=Iĺ���"��#���<V<�O���Nl�����L���p��U)�q�&��Aj�w�������S{�o4��|E&Z�����f�����U�^��-1�
o�f�,����TT��T�@]��@mwt��1�F��SϢ�N�0��I!�R4�­�����,�'�d�GܬuN�rÙBǹ��P�mrpX�d��X�c�ʓ�u!�k���2�Y<��z�"���q�M�y���� ي��%�)aiS���̜fV�>�?ϫ����p��KR��b��^��4��M,ؓ���׹+P��͛m�#�!��'9d�� 4�/{F���BVZg�`YeeLWy���� ��$~Q Q���K|f�v�U�a���덃=�59��"�\����,tseJ�#�H|�\v{�|�e|,3��"��렠�:;�S�� �L�D�?����)"�B"5����C~+��x�p���X09���縪*�,������;�Ϟf���u�2�}b�}�q'�h��M�{�Vf�]k�ޯ��?���\�n� E~��|�gq���΋;��Mkѓ�u�1��[J+~��7(|�����[��A`5N�+Qm�oa�|䆅�3�e#��
���|N��-���%X�P���d�C1�}�/�x�W1��:��^���F�η� �۞$�2D��q���q#��I�?�E(�W��>H�EIF�O��˝IO
���0_Q�Z�XGn(u��n5�-�1��g	Y�z�s�,�n'�>����)x���a""`�'�? f�6e����z����.¼Z�T����=�8�IN+f_�X��`�C]�h̾��[��bI.�\F��5���^�����<G��(�x��g��L���1��p���+��g��5���Fz��;�U�$=ԊP6�q�w��D���vY����,�>hY�`F�E�m��^�`���L��:(�s�:�B#���KN��-B�����OD�.Z�onRt�m�|�	�7C�DI����ÿ́K�^!b�$�s ���7��c�9��]�~ś�?�̮h ���^�Dv�YmH-�=f��TA�0�+P�i�{,�je��"&�:�#���,� 9�@��&�gr9LM���(�L��&��P��RPx�� �P5\͒U�4K�h�z�dZ��,�2J	�A	��#��_�k�r�K�d<��&�ZK-]��q��d��mb����;�]�D1V��A�߿O�r��&��ݬ�2a˩��)Q��y�3���$��uٲ�^U�4��q�xVϢb�A��Kx0�TL e�y2#v��4��egbO�?}/�-"*��	'�!�[s=?���$a�5�j`"<B9���{ʂl?�x(
2+K�ș�{���f}�G�-G>B��VPq�8=�A��,�륣��dD����WQ��uOK�USd1&\�,�AT��`w���r�!����{�߂U������
U\��.���:�"�g��wiX��!�s�3it4�c���vT|�P����{��u������0�r���(F�MP���E�
i���Ũ%u�� ��� ,�뀀�&��ɭ �x>�O,�a�ܹ��Xzz֊����|��~� f������]�	�����W�j.���ejN��)�����v�7��7&��F�}j� ��`�D?����~�XL/
v����8�x�Y~�k5�q)�Y�q��[B1V��2��
��N�<`/�p3���=�N[� �f<�*2����W�x���S�ʩn���+�hA����<�k7���,�X�q�$U����]�4_=0`��5t� _9���A���/(����l�=(�8���l�IIf��]��Q w��S��T�$�j�U�W)�>�̑�Y7�ZK�v�+�ݿ�k��y��/�	j� �/g�#�O�Vae��V�e�[�����p�^����%w�|mx�@�J��A������ZO�����kA�!��i�H�aD˖,@��y@�hHzGg����D��)���m��>9ӿU��N��͵-X�[F5PK	W7D��%L�*��U����5�8������ъ��tNZ
��]&P��
��y5�l匌�]T{1���^f5��}��lBE�D���+��lf��.�!��ؖ�S�����3���Ң��w��w4˴Ы�����S��e������>^�CZ"�B��}�%}�p�ʩL7;���/m˖W�q����=��HN7���$����ʣ�-N���0lf��*CN[����V�{��{��oᾢdRV&r��!���N@o%׋A�JסR}�$M������4�\�XM��Eğ,j4-�����	=,9����f�hF���^�?)<�r��P�N��y�]�D���y��巐ܜ:U)��P��'(���M"Ϸ�rZ�ʉAn:K�8��8M�洦�]�t��uܐ�?�2%,�_O�"Yct�Y��.�ө�s�K=/����1�����Ѭ2�r�yj�zTڒ_�mw��V�FM��MFp<B������*��ɼ�VK�b/g?9����&�Ɨ�WG�!o�y��߻/��$l�4>�X~�hp�#��n��ˋȻ�D^dɑ��XCX@��Q?�[c���K��@����h���QD�C ��2y�H�ك�,H�.��/�����>��)X˟�VG|��������'y��u�X�Aa_P0�i�X��ﷄPq!<�Y����`�3�e�_J��żId�~T̶��چGVR�1�3�7Km_�0E���5s~�[��FAf"�� ~�5,����բ������7e��]*�����b[c�*�.G�Z>��Cv�
f�A�X#��=�Үe�T����k$	��i��V<]U~u=G��S���ӎ��.��iaF��C�{�9�������-5L��[���  ǿ���{�}��%��X�
��ն�#ݲp]�#ʹ��CMq�"�����^dAP����O,�P7D�ɓ8���+�p���q.��_H T����/.=�q����[���%Z]����42��5������L3��7Y)���s�t�"`���)�V�jS.�k�L��?׾շI5;{�¸p��k\��_N��V�t|�~�_0n�{�mb�F==䆕���zް ��OBf)��h@��p�d��i�9q�[p��˙�4�OAg�N8�m���aL���8�دZ���޵%����o���\�e�e��߸�eԫ5g�W:����^���i����!�bWJ�?=��+$�o}���4�BdIє�$��J��Nm�w0 儞���Ӄ%x�pѰ�R.���:��S��-��%?sT�(&��x�,�=:.5����x�)\|����; ���?!+�l�7�f,sg_���$# <�,���yY�?��-�Y�`R���݄X�����Ӷ�Mg^H�i�@o�&���LĄ;�<�7��g	.K&����Q��@�~JS�����W���Q!���â/*�J=���� �G��"��a[����a_fIRlH���C&�����\�9~��Vk�Q����@��.	g�v�f<< ��"�.'���v �V���s'�+��&��'E�dtSׂV[�̋�!^�|��!�ކm�T��K4���?҅bee
���)�)��f���W��3��;���aT)̎��-
��=v�B_�f6鬞t(�o��>��.����1R��ӗ,�!	y��T�r\��7�a:U���\�e̴t�(<���u��݇�`�X���*�ױ�mM����Xqhˤ�bLe�@"q�c����$��	!a��T�T�r��x!m*ޢ�^�މ� tx���}���z���9@eq����k�*���4�h��I{����d6�7��K͠4�x���rk���֘��f�)�~[�H�A4�P��8��g�W���:p�]p����{e��I��/��Y��>
��|����.�~"=+j<�||�Z��28_�����%E�5>dkcO�6��%X\d���Չ���~�z�$V����ʤ���1TA�Kp�Jt����`XŢ������c���r�Y��.�Zm,	m��oK��� �8=�k���7<YO��m��S5g\?���)�x	� `fŲ���Lm>a\�52�'/�Ka� L7q�*�[î^ �h����}eǌ��GS�i�v�ň�{������$}���) ���٭&'�F�'�_m1���雇��F��a߹2~�o��8�!M44c`"��4���I1!g|�.`����w->:0]��b��}7Q�b7��`�q����x�ĭR��t,k��-��>ͅ�9��%�D�1r�Z@!�~m�7D�h�ȵ�7u���oJ�i��g��D�;y�k�o�ɕ?<�F�����4!�&��9���&= ���,nE)NbjkǇ-v�j/4����f�	����	p>U�֬C����K�fA�b�p������;�e.Bo�ǧ��}�\�R6\y��!q�F�̧C�W�6Q��/����^$�u_?���
��_��ˀ++B�P�]��F�~v���W���C���	)d��Ֆ�G	Ւ�� ��#U��6�Q:6�i#���}wZEg1����`�f�q)���x
�]�e*K=Q�u���'�C;}}W�?Z��<����k�St��i��i���O�ՕB\i��'����b"�z��QQ��|:�rz�:�~?T\���qZ&g:~_��$����O`�����Akm���8�S\9�� ,2e �a��`���H:�Zr�@��n������^2O��~?N���IhW����nj�(zC&աjf���U���� a��4ĵ��ʥ�C�,���,�w.�?D*P��������#~�1�%�T�>koL�0�(��-1�_5��D��a���_�����L�x�����CS�s	sG@�N���*K��p���<������U��O������h;&�Î�g1��A�Wo�y+P<``�3�b+���mӲz�ơ6;)^��7�m���m��"J��$	���1:e�}UϞ<	yʑ�P�X���v���"b,с�;r�p؃���o���9�ֻc� �D�C�^�dw��k�A�;�E�q8ĩ�o^��pw@9�	��uL��˂���a�p��W�����}]6��X���	%����h ~7�	�9ԷW�lRќ�xP��e�J>^��/ȝ����"~.���.ñ&���[40��(!E��}�*��� Q�qW�|��
L�$����"V
��H���l���~���.���!������@�	ޞ�\ut��K���e�#�ݍ	�M�!��a�Z0��P�}r���>J�ȹl7�
{�i)��ۑ�;&��>f�_�2�8�>BҤ^����B�������Lo_⡩����wsd'�P$e)��U\'Y6|f�@�����|!�hｌkw�_�_,��|�ֈ��T�lL
�)QP���O��v_����}Cf:���'�-X��pR�=��)�f��	�w��U�B�8�^��}" �����i@���G�ߥ�tzݾZ���o)�u����Ş���u?B.xҙΦ�سj	r��!��{k���Y)UX<ŕŦ��z;�@+�1�[�
�r�'��Q��/7�m�&$�G�r�-�]���D��m�lnzD9.#���n��F����Ј��4�:��7e��j>��)�������l|��eXQ�(@[6�)瓕�itR��2��A_"��$��b���b��ϑ\� �w�y��c"�����z1w�ϭ#A���a�t���,�Z�hPb�^ft�5�ϗKЈ�i������rM���m�K�]�S�iW�\�s<W1#�)�a������{��^哭K^CII������}�4?����z[Z��Ze���	�by�p<���B1�O�z�
�Dt�J��x�������U.�)�:%��&�z�?��D�|�`!OWsq�__�� Ż�Rʱ��oG^��#�8"�f��F���3.�@���5|�`gX�x�ҝ���p�G�Չs�I�Q���2N�fi�k'&�z�tU��s�={E��ٛ������b^����RB�_���IJRzG�&2�3�
�ML �ZZw��$Ȋ�(6E��+��PV���#�mn���Ls@�=��Y���椬�A���4nk$}?���e�-�K�cd:$Y��U�E�=x�?M��[��^l7�� t�S!1�3�"ޚ\ ��f՛�9j���ns/��R~bB��|��y��.�0�>���AO�cfR�~ǳ�Q,�2VB`�����O=2B��l���'�h>Ű[�{a��7��$ٗ,�˶�R�ɠ���ܹ��HP�oZ�n�1v̆��{u����X��E��, n7��t�o�T0T��3��=�5��e@�sm��u]�ڿ�b8�oS����baG#�hh�GH+5)��~t�Fܳ�k���L=��3��n�v~{�"�e�[D�O�!�a:��ILÏ��Ċ��%�ݹVl��uZ��r�AAdn�5@&˓ǃ!l.'�<r��mDL�Bd���]H���ʫA�OG�����+�	RI)��_UW�p�M�d�������P{�[����䅗��(���3B�8L�L�(F�{Z�xQ�U`0�9��ъRk�<���GPHwM����s���b��/߶u>M��x���*��U���L"��f�4��Ö=��LH�W��YJ��[*g(�ĳ�>+'["D*2�Q�P���p�ڒXgN�,���T�+�`z\n��U�v����ˬ�}��"a����g�-<kq�5Rg�Ds�k��x7�#4�r.N+g!�;�\d��d���*[R&�{�?������+�!E����1�O��w"�%`R� oU.ޙ�r2L5�t��ٓ�6?�pv�����.���Zw���
�����lc�Ƿ��Ѩ��S�j7ɳ)��ww%�<�/��R��I�ʐ��oVW몊f��O8u���,�@�n4����=a|=�+�Қ��kr�uU�_��w/>�:�*S�v�Q���X|�܊�e�<�I���D*�����e�^QA.�*��Hą!>�6�	�C�ܧ"�Րc ��x��h�3m��U�2�֑ �o_û���r�v �(w��TXV!"=\ْ��sN�k��Z���V} ��I٣vBs.ƾrd��r�Ff���m������J�� 2�/����Ȃ�}�˸�Aq��~=M�{�w��S��BԠ2��Jj�;��r��H��Z8?D+�	-_Գ`=q�#H��(�s5�}y#�՘6�;wC�<�׊~����ɜ��
�E�����`�{-�B(������,6�q��6)���װ��4�J̲�o�P�<QX*˼�����{�Wdϼ\8��&���^ny�����gvM���n`�+����iQ,�0���VG�3U}���n�N���Oo}x}�DM����!��BdA�vZ8�Ϫ�2�,��𕰝�e�\s��r
rf�a���AP�>�~�ЖMn7)��7EvS�w�{Z)v�E�e���u�.��"o`�w�����*���&�R>Qx�T�i��˲��� ��o*�,&�9��	}�����5%�t�mڹs�|!r��m7�i��sQP|��0����{=(K�"%p[j':Ȭ>�U�k�x�3�ɂɕ5�ŬA�g	�oCޢP���MK;��
y�kz[ �����|:H}��6�$�q\���PۍG��F�+��kB�����t½aZ��������G��<�2 `4��}�����¸�r�����S}����]�=��/�}wC�:�~�C�XyL�A7d"���y���"<���SA�TQيk����*/7Z��]�5���C�zr|��Y�T\�48�)�*�� S��U]�1���r��kBx�B�}�v��(�Vf|����~8K3Q�  ����.�#�P��*���0���<�DTAb���#4���cd���B��I7�7�?����!@�]��Tq��"�`$ݽN����k�#��$�p�7-�)�o0>W�A��֤q��h�$���v�E���UϻT��9�zf����oj�b�DW"ST���Xoq�h��PA�ZHMZ�ף>��D�i0e�=F�]�|0�5ֽ�ܔP�!�����q�?7����=��ܭٹ|��.��8�\I�?쨳�G[\{�;��`�{ET��aJ���C��nV�5 �f����#���R����vڒk�)8�C�Q}�g�~�f�uH�'����}p����)�"J���0���Oe؉�T�3�1'�z,V�F���&���AY�}��*�+����|�ϙ�����r���1���oH�0*C�7�f������T^
i��\���w���|����!�X�p~����Mz(p��o.b���I������r�ȑR6�vƉ~O#ѧ �5.��SL~����a8�,y�/�3"�6�d<�7[�S ��!�Q9�j���s`���n��|]������|k�ђ�Ր�Ȝ�ki���-��h�ԉc�|�����ߩ�N��!,0���!�6j��-:�ݗB��xo���0����s�$�H�1A�kQ��;�>ۙ��'PK�
2ٱ�e	����gg��.�(���h�͝<4|�]�4'���/{�eA��R��헗\�����N���'��)y����śs��mr <��ә���`�����5?�;�ûa�-�L��1E�����J��!���Q�g�g�$!���q�IIס^��H~�	����[$�$�N�6H�PE�:���{9����\ U
��1x�h7��mx�]�˵��C�׋K]��ƗF���Q7>p�f�g��V=�i��{_�;�G��S7�0q����� �(��PG4�A�je�J5N�w�q{D�����b�)�}b�4�ARG��vU�Y聪뿥wn��jPT_�ϊp��Ri` ����-�u�h�4����G&��u�D�pاS�;��kt���&�u���&����Τ�f%\p<�@�686��jV��IWo���r|��v�\X͋�$֑̑�2�����Za�_�}������X�/G�c8�:?�E�����%ٳ���n ��۰K�kx��b6���� R�EԼ&ʶ����_M�w=�PDPM�0v���I+$觉������+>Q瀩�t�4��eÅ2�+țBfaN��wm�i2~�:�$u��`&a��%  ��fa(ͷ��n@˰��T� �bl"%B}�Tq��a+R��6�>�\D�����oͼ5���m�U�)���:���<�tɱ�p)��r@d	�<����C1}��om�$�=t�b�_����	��^�*8C -�6x�2c��T�2G�Y����"�c�Pd���2v�#4a@�W7�m��T�?������S�G��m�JC�/���<e����I�$��#:E�/1�f�pq8�ø�5) ���Q_gY[$�f�&ʌƞ6����*(/_�4~p���0@b7&p(�#5�K[�����g�K�f��g��Au�0P ��ßf��8��yJ�5����M{��
��H���~@*��@[z���mI�nJ��������G���
��߇!V��)F�̲(g�|����5��{R-W�ŭ�YP�7z��A�����~��dx�0��VZ���u19]I;NƵn�T�����
�Q�c\i�j���2����Qzzaq�q ����@/w$�V�ɿ9���'pr�a�
DĄ���:�+�zk����º3d\���fi�Z7X��O1_���u'��r���4
���(�4����0����P�n&Cd�ۍ���}��Z=|�Un��[*�%�
��;K�ʜ�ƚfb�����P36f��f��`�
W�D[���.|�̄�׾��ɧ{x�,�:��W��4p�A��6����1������4��}i�$z29@IO�o�n�s"6�I�U��v:E���0{��1|�gX�U����@jɠ���lz�����4�L#����ԮV#!N�pV�|PeP�r�^b��)��'���sL�ڐ���j�Y� n& �g���q����m�]���~� ���tZ?V�c�z�N�?�)���M����g�=e�?U!nPt Q���3*W�
q��p+r5���q��p��������߈�l�_�Lx�7�5�����**�z
lv�@�y�>�F����"l,Qo	� =F�~��T�O�a9|�4a�k�%}#4
}�T�{E��qT�A	(RdY��2��E���pQa�s+�~e�1TA�+�BztOۙ��?x���*��0����:�($J����[o�}�8���)���Ǆ��C3��t�"7���_�&4���5~��؅���{!_-3�@���980���Ǫ~��l
���̀�mG����(���s����
��}[0�؄�X��;1�g
���/H�7�d�p��"e�
��.�<�5��'��n����i8������1��?�%D���_�c�
^TQ�{������l)����Asl�`>Қ,������p�
[F��[��t�K�{W�-	'z:9V�#�s�%O��^�� ��L�~_�:�1�Z��#sM\Ǩ�=����G[̝�"�|�Rb�N��"���\��~q�0��JP�,�^ܳ���ivO
b	w��;=a�f�T�3Y��A�8'���a�7���Zj�C0�Qn>��!��%KƠFR�I/��{���˞�Mђ���y_��H���K�OF@�� �Ý�?)�@�+�SA��,�a���Q��R�c��R&^X�9���sϿ�{� �\�D��FMZ�]��֧H!��-K���<��ǈw�����U���W=4%8���m0�5
�왫���X�D1��y�ȣ��}�ޔ�Ns�/꽡_��m*;�_�+>=���5��z�?C���g9-{dG�Xyo����9�xEbY�g̢�Ұ��5��$B'��@�&2Nz*w�GS�Q��J�]�YCK�3����Z�P�"�+�'���h����~���PFMpwN���H�H ?�%C�u��r�1:���1~;��şPj�?N���z(��I�/M�Z�R����M-Z�v��$P�U�_����EZ���8$Y{Sc�� 85���nn~����S?o�39�$�v�&�}Z d�J��;�[_;�	�l�)���`DX��t+�ll�釳�^�?TQE��M�X��%6h����O�q�J���[v�PWGzB�n��͘YO�5ENGx?�81�ä��Vr�܏��)�		G�_N�Ûg_�xVӆ>y�h�������q�[`�ek�taO���t;@��}k�\�J�Em���ݲru P,G?Mq2�iL2�h!Z�4�u����3;��l���I�ё�&�;�}��:���	bmzA��'���b� `
`��
����tvW�7#��u��`�S��U}v�� `����1Y���z�8�4Ş��A�+ɥ�S��:g�(�G�a�<9��k1tL�����)��5i��<b�O��A��tTW����Lz���{jR@N-��O�/�P�!�q*��*[��'l�#
��3�օ��L�>��: �"us�1a�l_��1���ؤs��t5܀�Ъ�h�uT��5�t�S�s���vA���b���s�d�46ѐ�'x��P�3⟻I�U����1W�LDZ�Z״�Q&��ܢ�|�?�j���D��o�b��p����O��O|�)�J1����)n�D�;ݨ���j�
w:﵉ �&+٭�=-��9@��!�v�ΰ����kǡ�qx=�D��/xĴPYѯ����Su�T�ƦU�`�,��������8o��9�B��T��WtR��1���殡���z��icM�,2�$44�v�]�����>��໙���!�gFQSIO"�BN�k�q(�5�;���xh����b�B����������k������М��1������& �68z�Mǝ<[^�]�ִ�Pd�a��o����(�o%��35�o��H���37M���sہ$|���Qt����%I����3n�__�ށ�T -ȗ)ɀ�Z����~���X���xB���h���x�Z��]N W��-�p@�^�;�i�D^�o���y�����?4�\��u:�/�{�㯠Q #1l~���:1BK� к<�ꚚR[���㰎xKA��4�Rxv�C�K�l㗷��+���?����a>=6�6�c[���g�93�),�q*юj����Fs�X��E�5vE'v�	�;�(�#ʥ[\�pp��
{m�Cz��;4cl�L�\s����ϲSH)�0����_�J%�tԭWTϻ+�oT۬f���O��ݤ/��䝘�i=�^'� �R
/v�S�zTA%��Ҵ��B�����܆�&��,��x��fKm,
�L�M�� ���ح��_G]�߄��\�ms] O�U߬�1q.;~mi��3�~�����WX��M�������$�D���R�E�Otb�����4�C��c|�⑂ċHGְ-�<��e�Q���VǥR7��R�"�z�FE�څ�[	�{�E�.E����x� |(�m�΃j˳G��i��c����A���]����yi�Z {����q�D��sd �� ����ȗQ��A:�.$&'?���8v�����������}J"-xخ�Ӵ ��?.f��W��zr���$-i��F&��*&���K����"�R���*Q����U�T���0�Qü� ���n���|��9]y&����NOO�i�����g�c��ΏkHm�.�~���T:V�	�_9�#��8ԏ�����S��pw��p�v�
;��+�s^�D��
a_��Z�?y��/���=�	� L����1e��R�4��l�#��=�)�Jz�<�^�����(�%'���b|�ܯ+f��X���=p�A�����
���|�1�le�b��&)g�vB����m�hbX���#�tz��[�e��I�f�x��sXy�����C�o�������ع�X[���9Fq c����pG; ݶ�@��!Y3No�m�^��P�)>���H�s�3���	8٨�$�����4<%����i�;���n.*��s�z��
U�������#YG���S]�F�m��Sܲ"�`����g(�R	1ERZ�ma������,���	����?Q���5	�T'?gdf��ms�����xn\N8D�������n���I�Q����P]�� KY��~tA�߲s�&��v���S��"E!!}�@�RsM׆��c����E�G,C��g�Y��
��F]_K1��$Yk3<K���T�(����9�J���ur�	�,�&W��Ô �M��ͻ���5t ѺsȔ(i�ZO�g*�����Qf��;21��*�>�D�~�n��� �8�>k�Gm9��ʊ��I%}�����QM0_��_Z���"R/�q�hq�`=#�0'`:+��bQb>`�����D�#��';��I]�H��{��%d#�0K�'�ֆ�vJˈ�к��0od���t��SYϛ*�+����e�T�F�2�O2�%(44�
7ܙH=6��ʻ�{}��2S�A�q��������DKw`��?(9�6x1ޓ�dnj�/`���C��<8j"|8����ys��C,M�RJ���z<��nm:h�$��Ǩ�n}���Nzh�q���Q���xP��\��sr��ɽ>�&�kT�cfT�T���b�-qLR�Bҙ�:x~��Y�����%����^�C$�a��(_& h�݂J�{���n���V٥��D���	�Y�?��]We��\������ 9�L�J��3�z�;�]A� �L�ƙ�Z�h�,h�H��JA/P���M�Bw�o������1O&���ę,�"V�o�v�y�t7�~��t�������>��&hVr�KE)�2�?�@W-����X��Y[��o��r �����StMp�`d��0��yn؈w}x5�˽�I񠆆B�='s��x�B���c (�țr�ż\��wP�j�d��3�6�_�Μi�%s[�}�K�|��2�@� H0Ga���bx���eQ�;�"��̍jR�/7�P&*�Io������=�����I���h���R�"sǿ(J
�n[kRN�]�vx�lL���h��LA1�����;W���~��k��EѶ̳p#;��\d�/O]x�rNZ����/��`|ߛq��l� �g��l高�"F�l�%����ҡ���7��S�����o��N���j�M��3�ϙ� ]k��E1�+)G�YYw亢"�>�بNL&;	/ ty{�cD���;Kd�ӥ@om�W��^!��%=�Qj��Ƹ)bË��9����PQ�I��ʲN%��<[�xZ)�j��VJ�]�DQ�Wdr�R�2��[�6E�'mNeE�?T����R�>���jI�%�g����6�3T���hdL?����⌂S�l/ޭ��di� ��x���f�-�Y�2�RW5b����D肜��Ǖ��B�"�T�t]�q9�b�tZ�/�A�	"{��g��-��,s����I��l�ɚI�3Z����D�>`�+2~4���$/��"���us���xU�]��̮1�)��[�|��Z�$/d�uK˳i
yv�z��9������z�u�����+o\��c���wjTN�ܝŖ%��o��Gg*�Hl|��@���"�&���VY�G��tiI�j�9B��}qϟ|�*oA�Nbʷ&���⚱F��!�f8(�����8Y�*C��V�h˝�|z��+�lS'��@�2�OLj��m�	
���+�b �O�	�P�t���TθN�C��d4>���4}���dL�.Ԧ�U�|};��TʶAɵ�Bo�b-��%�,б{�
@�{Ĥ	�.cq�|(������7L��6Ԫ��V-`Җ����0I����Pq�i�m]SC �n�	rd�p��*���� �A���[{h�y�F*�����(����H95!��Z5a��.�# �IF���pM
���y4�7�b�Au�8�|*kɵ���X����B���S��1d ٦G3�P��&}N��2;��$��q 4ѝ~�K����F@6�i�1�"%�g���у2��_K<���<�_@����+p*B���<�,Y%z�z �Mo`!Le/��T���z6Iz�F4�Hk���Yp��M�w.
��0�/s_/F����)������?\arag8�Lj��q !�>O��Z񩷂�m�ڦ���R���
 �.�vL���r��$�*  :x�&NEv��̳�f�:��P��?��&��0#0�Y��fᄕ�7��1�f{�<���X�����/�ab�
+!.�;R�/�
븠'>���;�ua|��F@s�9l��� �K�ŐG��������XD40���ǚ���_����V�=Ή��E���~�����R{���KTc�}5�:U������g3�!��q��Qu*p�t�'�F��r��~\��84�Q2��_�[{+Bu��r�ޥ\F�_|��㝹I%��'����G�/28���NV(�zW��$��.�E�\sQ)8��nܲ%����}w�/7s�J`%Ŕ�ϟ{7���o�ZS�"� ��6�	������]�F������)�ǀ,|'�6y2J�,����<��g�1T�o�ڐ��J$V/N�ь��aa<wE��r�hW��.����>n��P	P����H�Sb)2��!��/��f�A��uln}'s��xԩ�s�݂s�2$m��>ˤC�����pLv�����A�)�ph(�W��R����8�M7������qLk��c�4�|DᄴW��)<ګ�̼�+H�L�>���>���O�)�ʍ��m�ǈ����?��@�t��9W�ˋ���Zܵ����h�2��H6�C������ ��w�m�;߬'J
pֆ�������/��÷�z���2-@�[�06��*�D0�qI�L�m���i����EIT!�=�ya�M�q�xڬ�HB���,��E�4Z┐�|&�h�
0�O' �ba����19�yu9P@�Q���ki�iᆬ���)w��.?ʿi?W-_O�r��������;�C�m
&��L�����|,�PS�K*@"K7x��v������mI����rS���)�9��6�G���؏K+(�9D��<d3q3�f�$��r����,�`4���a#*�8�3�Z,��}�}oˑv�T�	:����ꄽ�8�o�M��%I��!��9e���i8����.�Qk��;��=������d��+���$�zQ�G���,[�L=m��<́��i���L�3�"oO����ȩ4Ξ:�|$�b�T�����G�4EVl6��h���i�D7+;����<��߆�mo�c@�{���Ź�����G�m����=S�}W�%��u(���YF�Þ)�ɽ�1���J��z��:��I_7c2X�ML���zfxf�x{wNf8��YHn��!���֚��w�7E����Y�ŭ�I��[�`��v��>~���#�`�UY�XK��������3�4	)>�>8�Q���⁁�V�J5�$�aRB��k~�#_b���OU�i���sK��+v�7LՍn�0ƅ�k�2�Y����gQ�g�b�4��K̮.�fC�E\��B֢�n4���1<�qi�V�I ���ﰚ����$aS��M�;	�s�
;�?�Ӑh0X��O��0�t�:ނ�*mR�J����y�F���"g�F��2�
��<�N�.����˹r�U��}x���������/7�Ꮈ���+�5-m �4�D�<�*p�JRk�ݪ�B����h�ʿ?T��6�tG�4Y��D·��E���t5��T�ZZ=	j������K���ӷ���7ռ|�Z���yaw�O���ҡ�М��޵�R�g���-�VA���,���M>��������-������Z����@q�j���ÌĴƆ!�Zpԕc�O�gL|u��Xʞ�2#ɺ�+S�tV��ݭ�������N�9���'s�%�n��Vx�����fȃ4\J�����'ÿ��g�<�K�K�
�x�<��W���6f�9&,�@�.Q�4|�bi�CY;{EP-�ك)�U�pth�n~{7ki�T�G��{�XY�pMO���[	�cIM�K��9/zl�����*��k���s�ܵT��=������a��:�r�@�6�t��Dڔ
՟2��@|yPzb��(w���cL�Y��ԕ��������/�ᨛ�1��6C�D���̆���(R�,.;ba�j?���pn*����aR7������!Gw?^����
N��6�c�"h�e@��+�0��;�=]�=vP�v��������{
�x�CK��w��b�_+��W�/ϓ�����<�n�!��E�Yޔ�op���"߃X����63;��^�+���1����	���3�tHI�Vqلq}_���0�u�KE�;�U�G�$�D��S����̫���]\(S�N�?�6�z���A�x��`�LX>��<{u��Wr����(U�H\�ɲI�^�h��	ڣ8
��܍�-Y��©�r����O�֊��x��!�Z�&N#���� ���+��Fh�8���	LB5H�Z_��;/	5���Ǹ��ۋ�w/1�jû����]Ӑ�3���I��'-��)v�L�:K6u;N� �Y>&9
:���9d���ڒ�5΢���n����H���6�<��)�u�����xN�^����ۼ�~����c��hլ�m<�K8�JƬ�,HO}���"��)�F�����Z)k�Cp���1�N�\S�q.����o��<U/���O��ʳ���ᲃ<�cM6�I��t�m�-�/_v���s4��&Q��}�bX�J򦜳v����nc�S�c�a��r.�gڼa�s0[��>p^)�������wC�Q@E	��lL�k9�DY�!90��s���il�Q�(�X������� �@�/�o������B�GT�l�aQXP��%I�FQ%�n�e�*�E����6g�$i]�9�#\��
�Q�cŸE��bJ�Ϥ�.�S��m�3^aꏓ�Y����_�}�.>Nk@9�7�[�����9�OG4�iX-R	r�L2M���1��! ���������p���zs���~��q�,�{Ȍ�L��0R�4�H=�'�*���������8uƪ$F��1�=\�C���58")loE��Z~�(i�g"p7�S"�:l���Yg��*,KG��T��@ٸ1#�́�w�"����DӴ}"��^�_t�!��5�ɼ�:�˽����w���5����*fXO�&e�Ȥ*,P�#� ���vZ�4�/�����)�"�u��mNx�t3
n�(���¢�����+8� qC]��_��ZZ���pMX�0^%[���@�P��UA�K@1K:Uz�} t0M��f\h���^��i0Ҟr���k�*E`�$Њ�����]ڸ@`%�ZV�*t]��vrֽ�}�kk*��w��Ɣ�T���i}>�ӇG������K�y��&U۵�S�pc��ԁ!��)��ᘖӲ}� �R�.m�M^5!��R�B
�����Oc �a����˄7�SD�X]��il�~���������\밥O�˄K�[l!s-�����+������ڀ|q�� vĦ�{��i�/�@��T�s�\B��!��4:Mɋ��3������@Vȡ�0�J��U�FAd����gs L�@�S���%4���_��I;�LI��n0sR�8�&V������ ҥ2!ϻ��&��1d�;��ڼe�ޱ�4������,)Īl�F	�`R�������K�t�q���d�#��-`����m.��)���Sc|3J�_�����!�Tw*r�Eھt��F=�>�S�g��(G�pt�u,�C�כ�P;��w%�+��x����AkҜ���h��O �W���K\��ORzW�A�U6��G���y�ت����G����-^���-t�V�(�Uel"��"�N��P_��lHo����m��,,4�Z��e���z�$��G^<�8
��/�ϲ;Eߚ�c�f7���hH�3U�Ο1aeZ{��P������7��²��b���<w��h�|q��e��j9��cZ��Y�����M�pX�!T,��k#G�^
����px�>�RP\"��ЅA:~�@�y��6�xRɇ?Kj��,�Ӏ�c��xӠ���j7�45���G6�ԑȋ�.�;N�zo!f�:��m��J?]��U.���m���$=�C��$�.����`�n_8�օF���Os���uG�uE+q��C�R�A�^���5e����Q�z�w	;i��e���at�0 3'v��T�#|����9��?��m�f�z��`�J��Y� vN��)k�V�?��]�Sx\uQe�ۑu ��+����(��g#;׌�x5��՗O�b%�Uk��:�鼌t���9m�&�����t7��F�����:A?Y��G��p�}�����Gu%/N\�A <si>�6}�?��lJ�~4L��lp������?���#�>����[Zv��l��x�-�`'�sFI(��:���"���}BQa_OM�J|IX{�x�M���b��W1=2�T�N0����>��,�%��~�z���Le,�Z�$&X�R=%3���na�ѭ�`o�Ag4��eP=���
�����ZH��ןZ0�J���`o7Ew��>���?\�]�HR�~(U�^��b� @'q{��7Z����I�
x�Y��S�q�.�?>,�>=�N�=�9S�z����6�n��2��!|A�i��>�ҿf��D������̉���R��Yg�No�\����\T�kH�#;�M�w��5�	���LPu�X8MJ
 ��j*ƩzO��M�`�Z��:�Cp4�`B��w�U��gz9���]l[�V�]��\�\#����J`V����<����w�lg[������ئ{����3��e�D�?�AMP�~��7'��Ci���-U�'=;�n��^�v�?fT��x���fB�SOօ,�{R:݊=�?Au\a9��h��'�N{EOc�d.D
�VRuf�V��6c�
DA���B������(�̈́1��Y8�$��꾳����Lo� mm���+]�����9����|T[,)fWa*ҹ��'j�T����H�q�4�t/%s;+��ﾰƬ��<xV��*,{~h8Oi�=�QWh�ݜ>)��i4�,��:�[�V��_C�8�	l�<G��`��`�l�w~�{��6��_̈�^:��;��g�E<���(�Hx8���'�h�d�k=&̋��	0�����`b6M(0�4sة��I���w�l<��(�cD��Y5&TZ�{w�,$<�����T�KP�Hm�h0`�*a���1k�%I�J�&�L�a���Z�2�x@g��xq[P�i�*-bl�Q�ʎ���R8��w����q&Ǫ�_���QL�]\�:�����R;K���n@5�Fع���h�t݂��:fh6t����[!�B����34A8�
[�4�HC>��.G4�|u�)C�p������L���ݑ"�*�f�GU�#X�*c��djØ33Q\���(������f�7y/CJ�SeA<6&jM���a���ͪH`���>>��׏�uv���uz��j82.��_,���o�@�q�6�m&�����J�++�q�H�E�=h�yS�$�C���N�iՊ��)�G�)y����Pg;y�m=]A�M�8ɘZM&o~0n��\�.����'EO���˓a�8�jjdL�⮡�V�L��Ҕ�� �Ю�B���=8��u뷟ZD�g���)~�t�>�\��Zz6�����B�=CX{��rd�/,#R�T򗪊��x9q�b���l�j���A��7ܪ�ƥ��[ʔ
�j|���x������ʳ;V�7���"�(�����[*�O���KdL�����U��8T�� �{��{4j�%^��ʱax0AY�槚ń�DOӓ�����ɑ����S���·���7#uJ��]r�f���_��!�M{��;6�I}�|8��zr@`"��,љ�X�ʴnDab�x�y����W7X�p�	� �g>H��x�(ǻs�x����3�@S�)���=>��s���&�����[��vD�֏�nldи+ߣpLyL�� ת�d[���|h�����ք�@}:}�>�#�0{����M�os��e��`Ģ�����r�M"k9��J���b�Ɵ����:����0h�
GT�n?�=���2ʲA�s@Չ6+��&�:=E{�iz[MV�g:�tH�h ���f�ys�O���/���d�;J��G���2��o���~{�,�+6H���D�`m�V�����S��V��@Ģ�s�%Y~��M��8l�ò�,�U\��LTp󽭰�A�B
�b�!���Gӡ �ig����Z�!�W6���0�sH�P����� �MF\_�U�xe��;c0I=�qCK��p����vPi����Z�e�������:�.�w��F�=�ݿ�^6G�+O�u��*p��	���*6�}�Gڙ�Ωz�?�8BѿV]	��k+f���C��O�f�8p�Ҭ;��x�G]B��U.q�|�1�d�g O)��ұ�fG��J���5K����3*>�SϟP�Z�t��]����ё[���r�Ek��կ|dό� �#`-�SG �)X�)���'�W2�����-R�F�A3�RWj8��Q!�`�Y]��_�<� �=�ֺ��i�la��PMD4�ǍFn��Kq�JG��speLTc/$k)4>`�Y��j�q�
J��3��'�C��TlXub累(y�=��i+��눽�Qv��O'9�g�"<��,��뚏g�*�q�!~�>\|�c�͟K�'�>���(,�_�P�sYnȅ�o�L��m�����llR��<���l�ʰ��G�F��� q�
E��co��ץm�&-��x1�*~G��5��y�O��|9��/�gyV��LA�i�M�W�vb{Ŀpj�{(���a|�R>=���I�#��KZ�l���������'�;gͶϨ����Fڬ���q�y0��_�h�H1,�=�m��T!EN�#���IZp�<�:�T��~F8Og엱ØC^~����6���kb�	ƀ�!��ʆJ=)�{�`Zs�q�X�x��1��іC*�_]j�a�ѯ�L���:��<��C �����#�6^�;���mk���M�-o��@b�A!�=̼c�����3��vDs� ��3��S~p��21���vt������e��l���U�GI���lw�P�|��ֆ-��[�4��C��vބy�qa:5#���g����srbD3��7�D�w<FFQ��wb�+�4��&��0;��)�����6GJQ��"M�3����\��_4��z =~(�ţ��-��Sy�t�@�B�D���w�L9b��⊵	���Sմ�%6�R����+䖢���3�����(�6��'6D���#��G������\!Z������~��O	d����0:&�GE|���(�P�c�=����
b�*���	�N��o8��p�p��.��Ť?dk:dt	�z(��7���TU��x�@�k#P��¨H@���7����N'��л���3D����v���g=K��%��2�L��y��l���+���o�j�3�~^���nC���/�w�xY1�!`������ƿKOP�\�� ��6��GL���K̐Z?j=/�J�'�#P������,=R�Ιpo-�LJO�>?���.�k��*��R �U�e`��Wj��\)���$7�6�͓�mN8[b cS��(:���l.��~6�Q�9�QY/�tb���C,_�/������|R^�.��_ 4��3�R�g�؜4��d�r���wlր0�Ḭ�1�����BB�ZSW��JA���n'���R2U�D�#�c=����!�M0'݇�Nm��m�1؏�9kB�6�uw�Yy�P�q'8�G�
�C#�Z�̄�E(1A���ĕl2���{��j;pc�\��c�΋Y��|T2���ĳ��O*�=^�q��H�,�NFi� ���t"���-�����R�R��=���9H9��Cx�ذ�Ի DKr"!���2��-�q
�X�WRv���5y��j�	Z�p)]���az�<����K[�4�s[�T���	�G3����Rw��[Z$~���}��!���g�F�$Ӡ��`��Ǘ�NU6$|;�zݳߥmP_6þ+O�⧣��@u`r߻��LO���Z��*�czY~�~;a)�]��1�o���γ��zʓ��c:�lE�����њ7�h��j��Ȁ��h�n�h����~ҥ��J�0+�4_م��\��N��#8�)�"q���_l닊a]�N]���+�bv��O`5�pa��Ax�G{�l������W�ދ\�@�9�h�F���]��w�<����F��씘8�`����$<���f�/�-H'��g���?��.6-C��0�8r�'褼Dc�Տ>��vIJ��o�8�J]����bWUH6��g�f��f4U	.�?�C�ƀ��c~Nr)���e�x�UW�HW�P)G�4�M$�N�Jc����& �3��ͥ?s�i���gV�f���]v.	�o_�{/5l�Scj5;������.6��yԤ�ǯ$�!�o����>@��)	\�\V�b�|΅�u�}B �Og:J �eT�;�n~-~����%t�8���fG?�F�!�/Il~�E�jN�L�"�e��sW�7}
8��=�#/���T����&%G{�kXu��b���Ċ@�4�Y������>N�%2ţ�<K>V�{��H�ח�E�%�^{�[�$s����,��&��lg���͎�Ǧ:�JzWJ
[s�q������1����?���%���&��d����Q�Ƣg�!x	����G����H�r8�������4�M9���S��DňU�`���'ϝt�\�ʞ�M����;Ɉ�;�Ը�֡@�JFH���
gzKY�������Ybm�Ӻ��s]gT�,�������t&����.*��a�ׅ�Z9$���֏�Ⱦ����w��)�Ch�� ������	�&U����=�
E݂����z�zf�$��iF�o�=�>jr6�ӻL��v�(ENf��.�n�	ka��(�э�݁�n"D������E����R�<&�-;7�q �as>���c�7���2�-�@��(
?ē1"��n����%��Ѐz��<��b6�O Dlډ0-����<H���{���)]ױH0�iE��tr��W&��+�9="aΊD��	c��������|��S��<�'>{1����3a�jb:��A�u�Z楎��$�Ԍ�$�dđq�wE[2>��_M��Y��=�'�Z�˫��a����#rbK��4%."�p!س��ۃ�z+а�[HI
C��g���-��/���	�8<���n��s�L��݇��U�L�4@�D�yl�f�{v-��;��QL�w?�eزW�����T,��{p35��ɜb�����+"���I~���A��Ɔ��ȥ���,��OÕ��^Fo�!/�!~�{�a��z������O,>Et���"�<�.� ��u8�����a�~R'�r3� �ߏ6��2[�K8{���N���TZ��uquᷯl���\����<wf�aϳ�2}n2;��U$���@]E��0�6�QY��U1���t��v:�|i�O7h��}�H���N�ฆ�(���qC��I��T�1>C:"����C�8D�o�s��><��c�����䴁���!I@ȟ��M*عN�U�Nc�� �$�RJ������a"2�ǽ=$���2�2��jB!�"������M���ָ�&r���g��Kή��!ޑX�wr_�X�1O8e�įy�퉇	2%Ϋ���NT�w	��<��pz\�.�o͢�+�����s��y��R�j;� ���Ӎ�c��=���(g�<�(��G��O��M���b��~Rr��9��^N��L+ː�ƾt�ײ��]�<�hF�����WO�U�z�(���R������PO	[��;3�F�����H�˂"�Ed�	 !�/��ɾ�w�x�����Aa���r AhZ!E+]��bx�U�.K+f��¾�~�}��΁�t�=�h�԰���� V�'�Eܔ9q�C�`}Y�����^��-}\�vťӀJ���mV�<~~���o�뤄���Fٻ�\2���*Y	1�X�y����e��n�u5�K_Y�(�4�����_�4ôm���Y�6���O���?&�6���8!���6
qgM+ �{2��B9`��m_p�,�a��7G���P
�l��&�²�e�L~`9\D�h�0����	-BAF2��gDڑx�B�_o�?>8�Ei�t�3�q���E�4��|��FFk�!�'����ZL$�&� �h��WL�\p�ul{����n�&�Xb a��&)�qs��r�;�~�|&gī�YY1��C��h/���� EIlV�u3D�G��a�pec�a����7�h��pMf"1q:�����I������i&���r���I8[-L��9I��n��dul��yO#�
W���ɜ��g�l
ҚG���X�9��ވ�,x���Z����/���#��ц�4��x�<���t`O���W��6`��GDLu�eV�2��̂��qm����6{d���գG��TM��=���S�)�a�����:˘�@D#O�g$�vI��.������}�z^S@��*2����0Q��.X��]/��P���*�[S�

��T����_��Њ���s7Dڪ�dL�ߡ�	����"��~`�9�1,��GU�f�6j��&�>��=�<N~�]���"y[��M/
}2��4�[�+sa��<1��S������EC�f7���sϿ�5'�ڭbs�	va�]ۢ�L�Oª�O� k�,��v0��\
���zo7�}��3^B�%Cx� ��"��m���)%�tFi��{�8�ݨ�XY`�y�҄�Q�����}�����,� �k}`l�HHZ��ɀ<�SB��5�y;�����$�N�)긒�!}o��P3k�f���]�@(�-ʭ�u��8O�͋���;�3��w/�aGҲk�^h~�gv5��y�YG�]_^��[�|���c���_TN�~�9�U�V{;�+����U�ZM��了m�Z'ݔ��$�szs	�	x��x���,��A����%��i�h��N��z�K0�į\�ye�Ff<�� S��7��MM1��N<��[�>5y)�o��h^DQL4`X�VZ"5�
D��b�FI�x9`o�Z�]��9��[i4��7�KK(3O���E����0�3�?�� j$���hV�d�w���|)��>�؄��-k�g |���|�A)�5R�GF�R��3���k���9J�T�U�V6��'�꺣TdR�lG�u|���G�ӓ;z�y�%W�M�
��>C-����2cѣ�Iy���\w؅��1e��e����φč�+y��HQ-�p��PO�!6�������$T��ױ�/ڸ?�O]�����Hk+��`����O�b��޾D�x����:��^��re�Ә��V~������dR�<F�VdP�E����X�Wͽ �[  ,�C��TH@���b�Ĳ;����d�6U�c�}�΄��<0�c������(��0!)��p���sU�+Ɏ��*����rЕ(^G�J���#Hs�]D�w�M���f�\�a�I���-"�C���O�[�[d$J�&Uc�`��^����r0��]���?J����Ġ�;�o�l	���'B0	���ȍ���A_���14٥�'�&l�,� 4M^�D�t\ٰ~��Gқ��V׶������:�N�{���P��`{U�pYT<�U����5����I|��9��ʈX����h����;�b��XS�c63�%��0�MNC	7G:��ǒ�C6RC�#t�f9M*|�p�;��֕��o#�t�0k�Q�۝���B8nG&� �]��������.+7���J�`>_�S`d��a E��hhu��?�|'M eo�;Ltqn�%������lkD�
�0Wy����>t:�{�� Y�U�k��cw%~��U�>�w�#�;��k���<πO\��:�hC�K�Mp��"�
N�i7�K�}�k�-�����\�����=��u�dt�7����=����pc�I�ꨈt0������G�a |�3d�sin)Jg��܄�M4���@���Kd[�҅/�C�'��ս�_���n+f�d��\�r������{7����0���8�,\���p¢z518!ś֩3G�TJ�jͻ�W\?A�ɫ�q@ә�>������+�|�R]�+HN�!�UFm�Ԛ	�x?�{�~Ow 
\2c+�3�E�T'O��Ek����7�ߴ��BOJ�<�9Q(�Ҫ����j� ��rW��Xmv�t���F��9J�=�I�۾��q%�j�Ra:)�G��`��W?!��_��7��+(a$Q��1"Ź���3P�H��/�bc�� {HVw�Ҋ>�W���Ć>��J��˅ȎƇ�L� ���GW���>X���a��um����djO(��^� ����\�ڱj��ςw�ׄ�"�HUd��B�y0"C#`�8;@!�n��B�`���끘'�Ў��ю�n�+"�ɜ;�M̱�3�aho��&���0��LC}0��đٓ;S%Be��E�֝�K��X ��i)u�:�@��%�7��Z�e~�MFe� od/��$�)V��e����`�p-��'�Ѭ��4R|�\Z��>�.��¦O�Ҹ�~!}]{�\h�z ��	�� 8�H�I�?� r@z@�<�*�9��������jk�����q�F*L��8~˳�W��T�tȩ��$�)�UMIe* K�����4U8~�9e���f̧N-�
������ϛC�"�+">.B#Ծ9lx /���qp��41��!H(��nJ��o�cɭ��6�u�a����gQ���(��S)�R����ơ��?SQ3&:�~m{�X%�ɱ��/�`��q�n�@�	r���ߍKw���A�fá�bQb���>�z�CfZڈ�=ƕ�P��#��(R���`e.�q4�P����,?Ҭ�᝴�<9�m�*L�bɎ�w�%��`�Izh1���7���$����_za+^�.�S��^�ʷ�Y��Z2���K�,|$|�xBA���S�m�:���m�!�!3� `��'4L�J�cP�[���{��N�~�u�8�OGn�!/Ly}�g�.O��B��B��FD�R��F�<	w���	!�p�!�S3:���W.V�3��D�1a�n�`?c�t�N���O�,�9�l���v���y0��]��i҉�MqS7ǵ5�s�%
2o/"Bc�қ�-�^�Q��@(v)�x�=�m�Xz.⧒lV���m���Jk��=BK�E��3���8:1����d��0I�D=��駼��j7�z�֦���C���9�t=n;;�c��z���S��[I��R���{MX+��c�>��� ~υ;˭��T t/�]��[�l<���on.óE����}i¶Y�3�WD��J2d�]��1��v�K���g�n�~3���1iA2�� ��B���RBV�o[�7;�4��.�8���dR�ĐxU����5�c�v�s<��2�K�(��� O�{��ǟ�C��RL!�H���in�?����Z)kTy��-r��B�P�Ѯ��L)��=�ے.�lK�9�'� ����ڃB/��pI��3����l��wO/�#��V�J�2�Lpr�|����,P�|���Bhۖzf��A�\��M�i�_�˜����8<�XI<1G�̴�ѳ��ԑ�����l���6ϲJ�#�����V�U	�\m3�s(�87��� ��d�	^�w����8� '���4�����7���K��Q�E�����}��vÌ�k[A�簵	��3��1@*xti-�����p�d�YGdg�.u�=!1IȳY�'����q/~k}}����O��W��m ��0U�]���ۭ�����g<�)��Q;4:���(N]"M05���ߩ �9�	�J�)����9E��JTN�3�?縈���c�c�1��sx#SV+����x�)��2X٧�>�N$g�na	NW�t\��;�)K����+EOp7`Cȇ���٣?���4
�� ��S���k	󬵤�"��7�ǧv�&2˙"�[wi��!�w�}B*�L��yУ ��o-�N��~����62�릙������D>�e��1�*.j�K~��(�?�$;I�<�%�� ]훏,��Ρ�K�Լe��I��ܰ#�7p�х����ǩ���T$�����h�k;N(W�`ճn�?�	�Qe����{�?	�e�:[���qcn.�5��6�M�v	��>��l�uR7�1[�e��M�Hr�1 3,B1؍�kkN��O����H�'����&�w�]�o;�O��z���c*��:��ȇq{��`j�~�^�	E0��e,�	S-�#(�J��q���A���~�� �G����
�u~Q7~	�v�q3򗐴�~O·�K�O�d��L5��єC"}-�{�|�Q"e���f�ۀ�_+���2c�V�e�F���ѽ�P)"���TƎ2i�������H�ƽ	I|;;��6�
U�����v�a���#���mJ�#�f�Y��o;~�Z�z��c]3O���i�I��'��S%�f�;7��?������-��Z�G��()O�|o�C�eyЊY���%����e��>!�pE�ZhT�`mV�nuk~�(�ﳃ�|-Q��'�� I,-ia�m�$��?�g��ȕ~����aI���B��oCB�(�h1_����E1�>�&:���nL��� �d=K�#�ޤ��o��b=Q�J�1��YX��=H0�����ص	h�2��ȟx1�ǈ>�*5)����T#r�cn��;�����s�Y�@cz��)���j�R��r�d�v �<������ ���d����먀A��Kj�H6�U�g(��
냂y��T^'O�*�$��8פ5Şc�����q��.�ʧ��J�)��7��3���]��7P6'�����!�:�l�ubj�*}W�(�UQ~��?"Ic��.���'J�zb�@�E��=J7�Px�&DzQ�DիA��J��C�E�H�emJM�R�<rxt�����>�:��~����9�?^=���k�T��}�j�P�G�0�c�c�Y|��H�wq��:]I>8�RV������gA#�2�P�p���ފd99������؛��p�Z��Pt!x[�q&�U���Y�
������R���b��kqa9.�H~����B_҈�9�m p������Pw��Q�	i����G�Ә_Y���%م���^�����}o�7�8�ֈ*58mK��Op>�i�X��S�t��X<[�EB����Y"��u��H���������&�a�k\�6��Fup���%��(_?��0z�:o��*�ݭ���/����䙥@�5�l���ct��9G��\G��_�f|%�f�2��A�y�����"S�S&͒��7K�IxS[��T0��d�k�Fx�~)�E1�F�7�T���q��	�e+ [��� ^j��PwI;e�����U���_=�@�75�o_c�8vÎ-��W�uA�}��x�+�`H^���4u�a`��XbbL�Xc����7�}�^
3�8[O���$CC_;��n;��_֖J����h�xX-�'6e�|�$��k�*n�b`�+ϣ�~�"�o	ީ_N�E�Z~��7x�GR�
���F�r��W�\'`t���t�P�����C����[.�m���߿��G���侑�b�,<���� 3�y�ޱlI~s�l�����#*e�&<V���Man���u�
�\��a�x���8��f�B@pڛɉ
���Ԩ��B~���i?*�XH�M�j�����QBC��~#�\�n���Iy��"
�h_�����h4$�:�:���앩9�V=s���_�񼘭�DW����s����r�7���ҫ��mP�䴏�Vd�n�fB��uG��1i�j��0ޯV8to�����y界��S��6`���L׬ztdXc��_|�"�w���yL4�B���xdɡ8��o{��v�ð��_=8ֺ1�{~P��I����x�bQ�o�g�J�7=s��K">�V�I>�Ϳ���x���D�ҫh��?�yrCNFy��$/���������Ea������?ŗע#\���_�<Z�7����4U��k&!i)q�����׎�ԣ��d����{8l�9�	��Oj)��Y�Q���[�q����ͷ����ﰑ���*���QM�\�I��g�ڵDȡ��*�ܦ.�.#G��T����p(�Qʸ�0q��ƓB���Ļ�����xv��0�`O�:��
���\X���8�5Ҕg�1�S�9ZS���
(
�d�p�����d�S�*"7j��9i�۫=�+�����|d!u�Y1z���A߷���Հ�������Է
j�����CE�!D�.��Fc���f�Mb����B}��; |�iSZ��A�g-�Y�,XC�'�hl+[�h�3>IonU:ʆ��_���S$�L.�V���@⫾w,�wF�᤿����
7�VX�G0v�8��&��i��Ac̮�Q�Pe
_�'3���~Š߮#ό+�����"j�>C[�;4��0�k����Ir!�=i #�ж�%o!{�!��G�~F�P<�Fi�>IZW�$�1��ҩ��)��{h"K	9�哱�~̟,��������Ԋdgh�U��!j۾��(��'�2����� ��z���?"�%O
���8Rl�3���j�g�}J@����@	�͘S^��I��}߄��,.���p�h�z���AcN�K��9�������X���{ڕ!7��"�$k�3�J�1ƾ[���N#�D���[=�@w��p�Ȱ0;:�?�RU6�n�E���0��e��QQ�Lp���l�[F�;��9����r$XxGPeKD�^��S'q'#9M-g��0x�8�N~aZ��E� h[�H��h��Xk�-����a��Ej}na���|7/6����pn�h.:&��{'l�/��쇤t*�'3�8Tl�ρL��V�4^�.�'��H��F��:�VX	Q����G22!��n<7�=o����Uje�2߳�d�����ZR{Pjr;�X���D�����Z��.,2�s�{u�V��8BJ���}�mQ;����]f��&A���|?8$�d�`O}�K��]��`�	�3[Қ2V���J��)'͛�7{ӣCa�͛�()ݑ���dE�؏m>ǋ��,#��pJ>fݙ��h���|d�wzŨ�����?�k	��?��/7Q
�9I?����Ȥ�.�γ��l�)0��:�i.2�(��	s�jݿ?I*����f���yJʜ2�Q���ng6���b$��|�'M2�I�;�@Hs5��|	�&��$���'��u��^�(J��P+O�ɫ^����-�8f��r��z.�yZ���iq+ �:J!% Qtr˥s�~�o30vm�tIh�(�Ԭ��J��}˓2�l�L�(/�ӄ0��v6/f�Åj"ĢW���k�����	{����~��1=��cg��.�M*���g�Z �R��jJ�KA����yڻf6���K?��^lS�mA�?�#�\�H���"!��J(Bc1L��{T)�f	���e�妷՛�xD�8(�+���_����Lz*��k�Y�Iw��\=B�o��"?ƣ��R)+K�]X�9]t1���8��rZ6#���׫��_^D�^�B7�i=�tv��g�N�eĲ7q.�$k���$с)<H�ˠθ(������~QB�߉��Z�xES;*�k��0�\P=wi�1�Ç��D��f�_���-bl�ߠ8�E �Z�b	�8O� �ZTX'�_�C�D�W�^J*�p$���N|�s7bz5��Jz��u�hF2����J�g04��w�dn�(*��͠��J�p�XphYHʌ����p��e_��+��W i�6�z�E�~)�8�:5q�KZN���%������B��MZ�Dy*s�C9�]�U)� :�l�W�R;[���'��ҧ�����D��E0�`��x�@�N��F��Dk�D ��Ơ�N��-��;�¢t�^�7��x�y f������>3�Ț��f�Vt'��S>�'A���Țf]�#H��)�D��ȼ�~�|�E��`���͹������\�PY&I�H9jr2����HX�b�a�)��X.��B���F&|�@^9�lv�eHS�l��qȺy�z�y�g��P�0ې`ѱقYbJ*�`�`��!�)�b�TL�����91x������dcB@Q\�%�_^瘩0�u@�#E���Ë�V�1N��1�JX��8���PM�q*��%R�����STr�,|c�v�؞�A4��(�7CAi�v�ֈ�w��֑���Y����RG�	[����x���I�	��|�$gWh�e�m!��~Yi�@F����pgt�ø�g�M�Ѩ��))�h'F������r�����ږV1��ȥ3����Q��pNñn늸���-��7/:�������`t��鑇'��L��A���p���4��۽��\ƛy�F#��4�2�~���e����d]:�g`���GN�����Z��>��O�����^��M��A�j^|(}]R���P	�C"/�d���&j�sE^��GO�PL���M�����H-��3�K��wi����S��:�ܤ��-h64�_ �"b�n!��v&��2,�{0$R��-�/"ng����/4�w\�d���D@%��i������]yW��06Ƒ����t�l����6�
�@-���W�O��TTLhX�,�*b�S�;Pd��I�آ�`c��5��?B�pR�PĻ[v�G� �K*r�3�����Y������_I	�%�qtl	u��iei��r��g��yx~v>��FO-f,��fau"@�4�!Gs����E�C���j_�I��}EBze�r���q�+o��sE�����Z�d�p�V8�����S�iu�>>��[t��e�ft����5C�[nU��,RR|�f����t��|@�s	�a��c�5�e�=��r�mo�S>]n�LSפ�YЀ�R��s<�N��%uԮ(��*f�!�UO���U�a��=D!�#;H�~��m�% ����H~sz�5pd�������47���n14|tp���$	}�p�t���r�����PV�:�/4��T6m��3`
!+>��^NS��K�{�|a�G���"��C���=�>^#;�&O���ip�,5&O0Q�>Uu�'��-4�1�g�M�e�4\�ƪ�ر���|H$�B��C�|�8T���ȭ��6��t�9}�T<�&iόP��i�E[�_%����Mf�Ke�6�7y+�{I3�KF"݅YK$�ss��@��G��e{����3¶�>Tʡ`��1v(Ųtz�����y4��Q��򵡫� �zH+�D���,]J)� �@�=�ҙD���L8/j�hV�^�i��4E�����M`[ �T4���M�H�u-͇c�)>)����}���zbp�	�E�.���f�=ڛz�YZ�b<�<i7�4��Y��2�cѩ�{�о~���.3��뱇���Iۢ�Mum`J�����^.���K��Y�J�8X(m�́�?D�N�K�Ĕ`i�=N����oo0���51YF��n�ٴ^�)����ɡ��$$[��n���(#��
�	�~]kRÙ��Qp=��K����4���%�(�҇t�X܆���7���t2��T��8��t����)�Z���+�ޘ�� +g<m	a&D��7Y]�!0�u����P�`����� ��q��/oa9��Cx9����3�U%���ݾ�6�;�{)���o�+���ʅ�(�r�	��=���p�d)�p�L�B�q��Ma��j�e��d�����1��VAoԔ�`��?.A,��<Up�j�4�W�K�(p^δ%���G�ؙ4�R�e ۽S�S�l��ZȺ��1{�ƙ���o=��L���H^�.�}��h��<b����tn�M��v����MV��"޻�c^��"t16H��O��u��p(���3�Ss�3��W�2��r��Y[,k��O��	�q��u��1����)�4(&�R��	P� ��Q-p���'�$�;�^�ϲB��2������͊��>z�k�LÔo�%����;=ǍՒ��vs��&�䢐�^�K�Vհ����gM�����Va��f}[ݟ6e~��L�*��	�w�T�s"�r ���0xݏ�/���CNE�b�%09�a1M�V��ږc�>�8� ��fkGQPC���O�VN�Vw�40O�&2�u���%�(��n�i6�J_��m��"���dY��`=��[�{�� f?=£�##�	�ӏρ�Q���T�M�#�A��TToC��n��^���/�x��\겲\�_��q�)��dPx ^��Ǆ��בx�?2"��ħX�n��'wݕ��-�t��1K1��������6�SG�6�{^��̮aR�:"��m>�=rع]k�DHF�"��H�ҖM�_��(?�Hs{�s�K��������멸M�ҳ����'K�'���j6�s�M"^zT&�Z�Az^1Z��R�27�O��R=��Or����㏠�@�5�ҝ�ȉ�Sɫ�!�F���T룑����	�3O����0���� d���ٵ)��6�ݴ��IMc���f�S\�n��5��]����oe�"�J�b}]*g�F5G�6p)@��k
׿�\]�x��n�1�U��k��w��o����c�1^tȉ^&�r�Sb��Ju�ЃBsj��Wn|܄B����|M�8�2����pu���J1��ȃ�Ӳ�a�f�>gQ����.��b���X�p�ZĦn��A��W��\�C��vk9hֻ��,#�D}MD��������k�p�%�;S$�!ZB�D��[`k���Clt�9`o���\��q�H>��**U7�뫡c$C����}��W��
j̍&�OL��E	�-_=��ٸ��{�Y�24>�J�M�0��=v��i7 q�,�v�D5o�8t���堲�!;�0y�a�\�>�f�j���Ǉ3t����2\�u���EN��d�J�&᪺�GE�z���P���j�#���i�#$�bZ����V�{=l�O��G�U\"��%.��y\�����4p_�#�B���Q��I�FK�nŶ	'����>l؅�[9�q;Bs����\����,��x���IU_x3Ί'V���!gO󑀱��Лt���0@plNȩ�"m�ʦ�����|�t>��&:R��b�v�OǓ��\����힖; ����'D.�+sñT�<t��կ���33QJpkb�l�����:;-%�sk���1*FܕϽ|���m���� "��)�iޞ���Pf��)��Х�4��]�-;.��OQ�BtC|��{8����*5�/t����Ϥy�)��<��F87������������9d�&��dK�De�+[���I�^#Yq�t�ܮ��i��X��8f�Y��$)"TL���>�@FX�#������lNϼ���L[��}�CfĪ��v�3��T����(!υ���h����L��)�!&&�_9��>�j��RgY�&7G�H��}7�pq����z�+E��}ty"�@z<��|��B�oX���[�~w�e\���+G���{�_�m�>�̱z�x|&��Ĭ��\>�~P[�3�䮆���OO���;D|�*�L�;Įg�OS�������TH~&�@��R���-������y�0]��sbB$�T�nG&8�\EP��ML϶w.�fX�&���������Է��>�o�l\ �C�Uᙹ�Jtc����5�iDXW�s���L'��^��#��w,Dv_��M���+��hC�U�~�a��|}d�A�W�ab�Ƴ�[*�ys ��uj [,zD�o�D�X��x^��û�����xn�>ٱOu8"��`���d�3_��XM���5ӫ���`(]
�mb��TB�z�2D��@dG1ِ7|�?��<nQm��GbB�oI1������'Uy�Ì�����b�Q��n��F��]RM������&`��y��΃�R|T���V�
���~���	��5'���w#��>�������#���+>���<�&���fEU�~���g�A��K�3Pw��))8��#\��x2#��d��x��U��q��q�Dx9��K���גf͉ip�Z9%�����ABg�<	�����E/�Z��l(�Nq�j��?�7d��v#��rf����w�6/�V c9������z=>����#�)�$iG� ��Tl'Ю�w���)��φb�W�H�7��{X8�����e~���Aetfl��^�N��@1@�8�DhY�-	)jep>A�d.�dߛ�?̳'�F��SMQ/a�+T�����<C�}��
J���)��!��"�'w/<�P[�Y˱�}E��zMA�1ȦA_%���|_��Ԟٷ]0N�Z&��*]��}Ϩ��bo2�/�!`1S�ģ�]�r@��<`=���:�"��"r���^����+~��K�l�W8��X�T�%ꀷBï3��#���w�1)�-��lƸÞ��֣���F�ۡY�
��oy� NS�}��:,ǘe�I�Pw��郷ꠖ�#�(!�i����KF]���"���S�Ǯ ����ZP	�z~|)lh��޴θ��0	�ߙ�'J�|��gt��[p�J�X4N�\�x�+[�����n�����°]'`M�c������Aw��M�y����|ߐ`��ؾ$���i��!��J$�o��<*zc���,���=�m�������#G�r�Ur�X�W�P�d��dBn���"t�C7��;U��n�_ܩl%!BG� ِ��hc����1��>�h��D4LlY�%� �2yd��O���?��l�#�xUE�H�7���v���9<����Ko����!�cZ�,��Nv܋;��Z�Uk����o��t�֟�SY*�̥���
��"��4u��hv�m��7��Qd��W��ʫ�&*�ffj^��~ntګC�\�<�-ڷb>o	3�?��d�o�����S��&�g5-u襸����g^���(j��2�=� !�Нt�f|%!�V#��x�Jޡq��-���yR$C�&�	x��3֖d+c���9�Ky�,G:��`�ͤ��/\��B�x|�V����2
飿�F�SR�#�{��%�${��ET��F���ȧp�쨍���RM�B�l"r`�;R`oqxɏ����&g�
���Q�:샱�h��ciU`xŚ�F��E�@i�6��؟#)���ce(��^���!ڦs������򠡁��Q8X���y�u'2ح��%����n�A�8p�fq�a8�J/u=e.�w숲
mg'���)]�*�&#'p	 Z��UW�fb�� -,���<������VB�8
KЁ�g��zx�ra�4�W7� �P�r/��T*JvE�ŉ��d�®�AB)��Ժ-���3bd�L�,�X�ҟ��+�����%ӂy��[��<٥
jWZ�?%f{һ��V�$, �&wLᘑ����0�3M����,�(����+&�E"n=d
G�u.Iu����M�Uu2B� �}rx�A�ʜ�"�D����)��葐�^KN�9��HuKzl�qE���q��ky��vw�M�R��.��S@V��w#K���ߎl�k�
C�-%��rOu�̿�4W�q���>�%OZ��v�a�`��=v�G�X�Lp-����! �!-��sj�;�Iq6}���`ic�;���s�����а�M��\�̱�>W<X����bǳs4�C����DF�w �GRIT�4$��_�[Ʉ�|_����Ӗ�dESb%��|G�_�����Pn��9�X˻dߡm�\M����I)�BSa5��'�>��^�*f�S����RM̲ż�C�'�Y_o�e�:#JpF�Ʉ�����-�(��:��3��hphԍIP��t4Xڝ��N�)sw�E�<�,	�koaG�qh䪨�:��TB�>N���!i��[�i/K��uH՟�E�n^֟�|ԉ5�K���^|�h�A����K���~+#:�Vc��K�����;��֐�.1qs��n��\��|Aq�Q����?x��1�t��׽��R"���ԱDB� O�y�ώ՜���%��ٓmA�9����S��~>�e8N�0'�s����:\�a���북�)��j�bܫ�(�6��ë+���R������?�A��[�g�s��>�wF��1�R�0�֪������_ϵ�i��Y�ADI�A`]�8O�qw0��J�H/�P�?�M-!CJ���1(;H[�,�1��}�9�f����?uL?Vt@�H�)���wU��_/�!����4~:��R��iTt	5�H0ޗu�r�Q㐴����>�t�U?�@b,.Q�@"�D��9�t^��6!Y�~��\�Y�hSh0�n�Z��J���3��\?���4��Yz4:'�����aGVx$�SiXgD|����*�͖���p:`5c�FY������V��*��m�y�py�l
�5rk{��Ӹ�Jk'#F@�T�x����]w�K��oǵ64���T�N)��:�(�98��~'���?Zv���?.R���s���_=�����;!P٣��;�%�8>�~�{V�Y!аi�	�F��N�ϼF�ѿآ;|�h���륿���v&���טY1X&�鯄�f4;����ɲ�+P��Ʒ�Z
k��-<U�����ƍ��o:.�����,/ �
dy�)��Oˊ�[�ƌ`ƥ Y'w��ޒ�Wd�(��H$� ���ѽ�E��� ^����68�>t����"R�js@���i�����a,��?�����ʷ�;��[����R��J%�7)#Ǉ�Ǳf��E�l/���(]9���aʡIע�t�h�H���s�]�D[c�(�JVF4c�g6�a�-��aG��츼�b�q&D��۵FM�{~�zV:O���ڂ�9c����v�rXR��4�qA	RJ���.�Y�����>g<��\��?��Z� �Q��[�u������ZS��~�V�W���輻m��& �
m?��l��w)�,��ә�
��+ˁ����u;�1��i��9f��I��K`�*=Rt_�qe>g�@�!c���z)�}��l�@w��]�pY�R�^A��\ޠ��T�.E�	��c.�'�M��0������Ȋ"�"�;����M�t�{d�l�ퟝ'���19UH<L�A|�#*}�'��;�x�����eQ%hm��
��VЗ�����;1�0a�� fJ�j'�{[�+Wl9 ������;��!���V�R7�o��kM�4��]�'O�&���:^#��(���)�3Z������i� c\��N�E� �p���F��<�
��i�t�	���}�Xe
w,��J)[˷sNƠ�o���nI�!{c�DӵPL����&�'�
����Q�
<r�+|�Co���H%7F�F~<psZlw4+[ebK�NƑ��5�x.觇���]����p��!�����F+����[�f�o:)���Z��3&�r[-O֧IeZ�i���O��*��؀ŮNm�"+��$4��C���c����M�E�|h�KBm���
`�7eP k�^HD�	�{���4'D��(�V��MƋ$�'�{�/x�5%O��b<~5�>k�_R,/���l@Ǒ��H��;l������ឆK����w�pH�#�] �USr��4�����:�	��f�r��V��z��BQu�H�4g���L�t���1Qw�R�φ�U��9D�I�=��8Pi�*��|4�j웤y]2y������b�G�c�dHd�0D>�����bs����w�pg� 3������&M9U~��<��#$��L!����x�y�.��m�Z��j��U_���9��Ƈ+��D�Ֆ'�ʮ��������1��yx�O�5����'=�u�j���{����z�%�����	�66��P�g6	<����DC�wGJ��������[�Q}s�9{�uՠZN�5qq~��"W���<�� nP^ɟz�5F�s�m�A׀*[3i4c�?[�h�@A��.���ķ�2��vs8|��I0�a.-���kH d�]Ui�C��(�;�K�{��r�����.��R�Vw�8|��]߯�/��ʉ^�9�e�]X)TlH%8���36YG<H�s�C�֚5��ۈ�?�A����fV��-���iԪ��1h�K���ŨOP�����1@��*��'�����%���w�)��57<��y>yԓ��aW�A�C��S'���e�n��(,`99jq�f9�q
���(����>h��0�/�]}Ήn��Y�Py�2X�Z�"
�Z�q�/�\�X
�$/CĿv�Y��K�,Z���*._������	j�0)�F�m�_����io_���w�^��א�ٸa�|�Z�1�c$��[�J���pؔ�]m���o��	c�y��JF:g� �{��+�f�]M=���Ht��ObU�dt6R�ծ��[
$@�Zת%hԼ0!hZ4?���<�_8&�@$�}�6
h�_��"j���J��zB��>�H&�����Iz�V�*R���~��)o��zq��Ѓ+=�OIG÷Rv%�>f��G[�A�NYx7�����g,���҈�9�=>��H�|���a����2K���G��%��՟��֊���A�J������e�a�A�GYF�PG�ä�����E�'2�'x�nw)G{o��r�_�`�O��J�F��"�5���UsK­G�6��lT�'����=�_�8Y��i�=�?R�bu��r,I�SWFz�bJ�Gѷp�FE(�è4N����_6�))"2S;VM�ax���ڋ�=P;�`�8���]P��'E��R3�R�5e��;@�IV����j@�a�@o	�/F�C�\>Wٿ�G���p�y��:�7P�gs�3���>C�`�6�
�l.D�ڈ���9w��W���tb��S|�.g�]��mS;����R"�2��"7�8z�w�D��,~_��{�B \����T�J��j�r)Sh����#�Ŷ�Nv�ڕ�iر��y4�szs��R�Hw��Φ��5�y]�%l���\p�ޚ2�̓T��[�X�"�XUw�pn�$�E�a�qL.�PG9��k!�.��3���sZ��(g G���M��$/z@�SkT��Hu{�Lq�N�'�9;B��}Fs(	p�w�ȼۇZ���?��a:SӌC��7R8�đ�h�ћ33��̰#����s�t��q��%�Cf�>�Sؿy���?���M04A(�Mz� �+�o���hL�@͸)��gS��l��O@���)Yz���a��� �٢��\��/^���H8g3	 <�S��ڧ�f�"iTT3x��K;팟edN�f_C����
�䜅˒X�i��7q�AL߃�qv�a���>.ˍ4;I�R���Oo\��%.gR�]g�<MEP���� Zo�G��.�	0���V� r�>��²�}I�
�t�ʺʑ���&[��H�����:i�լ� �y�?��%�����K�|�к�kֻF7_��O"I���@�Z��n^�[ޚ�l�Ꞥ�?i
��v�ڲ�}��5Q�a���H@u��b���	|�,I��E���"���[Bx�u��:	��Q����٥���XP�����!��T��}}V
 .dQ���iQl-g��8�I�F��Yn@m��۾�es�J��=��]�2���N�
��-�0�,�"�q�i�
�aQ��[�Q���p�4�0���<�s���3��)���w���q�Msx�������>̿~n
�Q
�L��(�m�R��ޮ��ؓ�[YOT�2~������~j�@��$���X3�d8�J{��]�*޾�"���� ;>DA��h���|,u�#T�:K#�Ka<n��@:p�&ed��V~��S9v�F<�������W���5W0p$��p���!n-��*��4	�k�r����/�]���w!RK փTsJ��묅�S��}�}�*�"us�4��p�"UJ��;FU�8�W��{[�*y���&]e'�!S+�H�+x&���ꙿ��9��K�YB�z �+�����W���i�8�5S@Zڮ%!Į)�^ϸ�#�\! V�?Rګ�����c@"�f������}6��n&$�HK?\�w�s^o?T��̏%�suY�0����W�y�KlF��"��(K�k)\^v��	ȏ�-��j~9~et����ݛ����BI5|�T�F{)��L' �k �2��W���C>�Q����wǮ��@���nֵua�xvs����'��(��~�x����tcd�\o� R{��H�y�D�x��Q���u4Y�[�
(y����.�H�)M�{�g�㥱ǯ�up�o>��#�uJ����EG�H��͂�j�55s�b-,g����_U4M��.ȝ�|�d�Ӈ�6�Nz(qx\�7�����.�2"�у�R� x�N	���vP�/�W3\f�mKtZ@��]�DΛ���-D>�Fm�d��EJv��%��>��7���Tr���n���)�b�9ʟ���b�T�E]�ؖ6U� �̊����]Ȼ�ծ����D�+Nm`/4W*SQ�``��H���� 4�Ϩ
��K�̎5�:.�����U2i�hµ��W�<����(�t�����~��`�Ά4�z������.j�=�mdg�P���T6 iwP��e��i*1�#k�����3���Kt�$���W=���O?I;���ƞ��1��퟉b"j��/V��������`��濆��TX��H��jq��ȫ;�����
6�Т4c?�)g���cQ �¡��[��;�� I�F��WI����fr+�+���v""�x��BBu@�e��@{+tB��)��WaVKTG�M�^"d�&*��s�����W����2f����h4S���cT�����-0�4������S��s5�K]%�z�K"��݉c�ĺ3őb&0]@͵y�nͫHU�Jj���9�2��M����̃IL��M7�x���x��!�u�n.�{�As!�T8�UC�F�3q�
.x�5Y�̰��MO�X,�����X���[���,f�fV\�6���Z�x?��{���F���O*ㇻF��\y�^���s���B�vۊ|e[�%�=�C�#B��М��ʽ��Tѥ�! (��zvc�1ȥ��Ȕ�[Ҁ��Hb^��0,Q���l��7 4�BC�]��_�\�'�3�/�����6À�&Y��3�)q�66�҉�S��BC��������X�T���cKBbA>�-�ˀ��0�W��i���Ka +vO�g�]v�N<�q�i�H���,���0I�c$�������+0���E$�N�^�n7!��H�c��ӹ�a�5���	�Q?=���5}�<q�ٚ���ڱi8F�s��V��H�Ox`���+����A��Qܘ�I��h^}e��jt��~=VeZ��f�	69k4rwg��Hdƒ���v�Z�H��v�Mu������Ŭ���Ϝ���������w�m��e)�Sa���[�tF�g���\2�>ܓ��y���\N���KZd���Dh��?݋�@��%s�_C&�����%�H��G�[�ź�'H��؉�9 �?�<)کr!�)A7�`�O>���\
�,��� �'���%�ğ���9��B�ri�WG1���[H�n��#$y.���(؆�M@EI�\)̧/��AC�XRL�]�[42�q(����p?�'�yF� ����r�1�H��g�̵M��a�� �N���I~%`�Y�y�K�w�Cl���̯?7�4ݿ���.��a������
=�Pexמ�)t�P��۲s��N�
#.$-|Ԇe����!ٝ���%��6���˛�mxUM`?��;<�Ѭ%-�"��z�9�d+W�aj������kp���pOѾ�*�ԹM#7��3#�H@�1vj�9)�6�Um|W���Z�:N�?� �v�7��%^6|M۵�����i<6
b��5��Z��o�h�p��Bl���gԀ:-b�O�7����v����~ޖ���p~����6��Hsx�f���
?"Qc��������U~�ߐ�J���v��B3w���s�M�c��̀���ɚ��`�����ͽ,]0���dL�;�S+µ�/D瘀|�SM�\Vwm��_?�����4�ixO���Ǥ�.H�6�;v����<�Q��V�+�h�W�=?�B&�3�tBW:F�K}Vf	��	����-8��F�ٝ4,,�N�C'Yn��g�T0�X� ]A3���m�'Ə�d�%��D�V���´w�Ò|�I�HP���MP�?]�n���z�X��"�,z�򧋘�ĭB�� d5��4�;g���~qyL�IJN�;���c�h�~�1ϲ�4����+����[�Ocr�٘���i_c-�������4Ġ7^��G���ĊҺi�[��xd@���ͬG?��M>�#@N�Eb�O�0��E��5�
>�W�J��}�g��T�"���VL���%�ɡ��h����w�o������"�hℰ�'x��k{�LZ>�������ө%Z(���@���5��c@�E/vj=�b��$s�l�����m���n'̨g�HJF=z(.��(��e_8��D�̛B����cZ�x1�S����?��^W��~�a8�
Ԩ�<�C���aT����	��!;t ��2� *�n�3�sQ���W�tpY��;��yJ����q� T��N��V�
Q��#D��h�МZ��Ӳ���8����k�o	��$j�_����'����@>��g�;��J��tR�Y���1'���'�V%'+FXAj���}�BƂ|5w���a�t6��+,�񮿲��C�Bm��^�?��$�25��k]��y{��Π�E���6Ze� ���}Z7�~Ў;<mp����D��!F-�3C��rڱ>`�m����X/�2/2y�XA@��.�C�Q�w#R����3�� Æ���,;rMt׍�B1����**N��}�d�PJ�Y���!&}7�@�B�BW?zq�o�C��#F��\���� 3*�*��x�N���R$�+���/�lK/P���%�#����v}��r,.�h3�������:�Oyj��E!�BB�b�H]��#!����]�M;�������o6��uS���0�5�,�VU����f��(°l���d�'z1ȥB�N�#��x�	Â�w���;��^1j &�K�^��%��njk��3[���.%�A�p
��V�}�H�oA�Vi�*^�Z��$�M�~�l�#V]�qnt��[���h���|pQ�_�%��C\d[�eJ\��Nv�	���+@�Ċg��(��{[�6�Sy���}��ƍM顢�c<��dRH��+���i�?s�6�Wk^�A&����W�e��*N��k���n�����nж���$��)�}�mE#�+��|�w�W@W5��I�@�ZW��L�P�J�XLs�o*!/v_��U����U����9��O�]O���.4`��?,�z�q�v�
M�C0ώ�Xh�ik���8=y�H�fU�'QiԋV|4X�f��Y�䲡]����k�z������/��l��fє0mY�F%c5*�q�0��GIzB��ֲ!��:�˸�E���6�����1���w�9�ʳD/㤗���O㍣܏ܼ�u�s�P���Ў~umB�/&��#��͛	}�� J�n{� k�J�r4�%����"y��DJ`ۇ��w�͔�6�+�jB#[3%)_�)�Q�:	O��z�g�le��Aͧ�?r�(�S3[�m����Cv���a��da�%�ll�g�!��[U	H�5���|��̐]b3�9:v�C���+��G"���C�8�
ϔI����'/C�7�ZD q�2�����1����~lJ���>��И*�*!�����z��تT9�0�	.���v�Ik�-m�r�u5���M����~�j}2\���r���zvH�1����auO���Jd�.)��qﭼ�o��|w�a��dW���f?����M���|�9�t.�@w� �k߲��k��Lf�ցKT_��Aø)�HFb��/�'�;*�oW��M�t�������
׬хSj�b𼽍p!>Ay��]Sf�<{5�N��eG�g3)���#>�-���j���Y"�\��
x"qEH���k~�(��4�	O�<� �d!�ߒ��6Ev.�pt�	;��.B_E�@��S������8����3cSֿ`�è]�&�P!Y�ւ��s��x
t�����)��E�|��5�M���Ձ�7Ւ�к���)F�� �v<얮�KlY/����L���[�"~W��E�ӞH��˷�� ���
Vc�ׇ9
���p�`�l��@�|�Ua��'��0 �՘X�½:ٶ����ݧ�#��H|����(�h�����C:�?�_�q<��A�쉧(7���1��c�.Q;�W��Ѕ�����H~>��@���e{�����M��x?�պ?]7������X">��
���4�&Q�J= �{���< ���N�pqQ��x��y�Y����ǋ�|l#�]�ӽ������"����M�]�'YW�R؜��N�
��<�OdD�H�����l@��A���B�۾QAy8��ٿ[�O�:w3:�� Z֞��LR�ژq6� n t��a��j���|_�'d�읔iX�d^\/��� @tk��\�y���WE�k�U�=6(���"F��{6⋇�"����W���pdYc��Hx���|0?-Ͻݚ<?�����)�-R:��`<�_�T����C X��?5E|EaqP<��}~��n���ż�,;�E���X$��$y��6�ȸ rǆt��x�W�KW�\.��5�4�`'�ەM�2~g.�V���l@��)4��B&���2�s�1x��/:{[���{0(�E ͫ���1�1�'���
*׭�h�4�/7�\My�G&�3>e^���'IVZ��O]���+M7���7��i�Ȑ�"�۸�]_j�~�e������&��{��`��t�C1������pe=�&J\�� �S^Ä�j�4�q��m��;���� �����$"����ig��y!�6w#"^�\����.2tT"l��F|�Ɂ_��`��閔oݹCM��+A�%U��-�`�9��L�ai/���\�Y��Imb���6ejH�1��"p�](���`�����w�׽�Ӂ��Ƣq�� `�̭ڭ���>Ha��G LY�!̈́�u�ѝ)4�OR�x�Rw;�T"mΰ���;�G�;�.�(��06G�Kf�$��l� ��u�i�s$�ܨL����׷�ԎN,,`L���U?Ϭ��D�#���B93��]�P�>]Wd�*o���zA�gB&�����V� �N��F�e�i!�y*C�Ƀ&�XC�b��5*D��89<��B�$B���U��BMqg��z:K�$T�iǠ��W�����.i�
���x��xܐ����Dy�Q��?�Ǒ*�4� �ʧ	�JH����^�<�X� ��5	��!�1�\����1:�x��Q/|�xW}�`��OR��İ�#�J-��"�,�CV�W�y�=��Q���ւ���x{X�w�ɯj�q�EI�#L[%Q5�]M�Y�]�U��&bwI?MQ9{���D�W�u� ��!��\2)��P��ƞ`$�p�Za���t`�l�����Ǳ�;����;[�qcȁ`�"��'�ͽ�4EV-KRz'2'x�"����־���Ľ�Њ�L{o�N����!V�h=��*Z�0f�T�zl��-���˓lV5-O݀Κ���_����2#qV���%�aqk��i�X�h�� h��lm��:GP��/�ԓ��ew�� �k��,�
�%sn�o��]9?�.�o���E���A��B`:D8gݲU��Qޒz��ˊ8l��L*2�
Wl�n�:��N!�-�mtԯ�踙L�`h��$�����գb��s��!{�`�������a�_��Y�0�J��Vi%��1B�V��jnĒ���|eHA�åp��z�I�T�Y&�����P=�H=r���9����s�Q�O�t��̩@5��s��8_M]���cN��?il��{☝^��#"XJ
���z�J�[Q��N��l���8�o??�\��U�(n���gQg��w*X�����b�%=d}��,%[�C*2B����h� g9���/�^3�q���	Ӏ�t�#�u��l;�
�1��h-
�f�՞�� |�E���T���lmP�$���`:%YE��i�[�ѵ���ӈ������P
������	Y�fZѠ#Ud����F����&e�k�l�Š��T�ʮ����9 �R�y�[�s"<�T���i�~�h��hϠ[#��L������~�fKf�<��DZؾh�f ��&��L�j��u_b�k_G�gu5e�beS
 "����j=N~΁�r��u����3�A��:�Ob^k�"�6�o�Mʤe#�v���:A��5&�P�&�S�$�֨��9Bp�ًGM�ڣ�\'�G��_��A^@ ���9�D������]_y��{�nc���H��N�j��og aX�G�l�QȘ�2*s?b>��dp�Xw����Đ^�7ʎ���D���������r"P��mS��P�vױ��V9��;lg�.�����>Ү]>�_I��������0'�Ed� �N����-!x(pa1��=����.�EW���]E�A�L��wV��
���AlG�(��5o�u���,}���� MJ���ӭ>\M�;Cah�w��S��ZZ����
��\��#wC�7�����mM<��������Ļ�G5C�Q���EjH�s���H&��c�t�a�� 9"�!ϒ�H�aK�wX��_}R �|�\~MKNv����^cJ���2�4S
2�l��Vd3ny���V�n�ͫc.״�@������#�?8/	�6I���`ZH �Z=��l]����I���9Ϲ��(�|KZ2�;����@�%ӵ�8�4�Iq��:�ɜHp1u7�g:h��ns�_99���@��6�r~8T��7�z�9I�!s��R�r��l�nJ4v䠸��Y{щ��Lk���Z����0?Z��{CK^��y'��J��X�e�d#������y)�%��l���G�S�����t3�l�;.�ȭs�3���&�	JJی%aq�$ٹ��;�r�����i ��)�nc��uYV:O8�;`���	�U3����	�VǎӒ:��H 1�a^
>��Y������<��������S��h�ʆ^�
 �;	�����jjM���(D[z�z���ix�:^�<��`+Tb���),J9!�{SB�~���#�o
�*$9��7:��e�w���P������r��o�����s(4����+�>)��̾9�8��1�	ow#�J7���ꨫ	��왫���ǅd_�W�%�µ�����1���-���X�N�A��0�"�i26�~y�G@�lƝ"2Wîpz0gM�b���N9�VH��:]wg_[��x,��������n��圜���*��E�2s��Ls�M"Оo۵5��S��`f��Ơ����$3	X�93")�6�����M�0�U����05˺�ߨA�"f�����)zP;ȥ��g�_���Ԑk�j� �P�K��=�jLX"3/T��(��Ӏ�8&�酏ե�$��B�Z��&a�<5|�՚o���go����8ID��,���i(V����.|ȿ�O/��Zo �� `Hb������<�j�P�G��,���D��Hkj�v�n�כ�����8����ʆs�˰VK��w���S9��9I,���z(���̨})8P)=�\sksC�� D��I�N�'���x��ƫ���tʞ�bG��x&�qQ�n2u���剫fP6v:m��ڛ�y��>S=�S�=�"W��k� ��������5��)�_�n��Ȩ!9	a��A`���+k���u��r�9rs���)��#�D4��G�µ0�DG+G�TI�t/�˗j�s�bo�������)}4���p�h������d/���Yb,0ͪ΀'�Z���H9Xb�
�Kؐ�t�}4n�n�F���'W����BQ�Q����3�EB*)�����?XTr�,��E=)*��S����f�͙�!�T'1
Wv��W��T�u�*�<+��:;jh� ���a3��s{�x�>ֿ��#�AØY\���&s�ʜD�]��I��w�ND���T��eSȶ�/���-V�c�}�rt.3
E�p6Լ���xU��Y-���{X�ū]kx �����)�ؒ�OA��%�.��5F7�\vК6���n�,��xN�D��F��zJ�KV¦�n�T�����d)���iq/��K
&�����x�;�%��ެSB(��7T�h`�yyζf�~V
Q>����N�������hb���(��m�����f����ԟ%�b�����:�[��2�X�D�nH�Y_*�pV���sx��3��CGhB��e�H�2o��O��"���~I�� ��
"fC<���"=]�� yƹ��Amm��竸�h�@� ��@`Aα9��|T�wR}7�-�M�`�4�@��TD�����ҹ!<"4��}ԖK󋾈����(T���b-��k���&�=�5��U��3U�#�'yJ��8���}#ߩ\2��f�y3C���Kȉ7�3����F��M*�G����r�������hT�=Qc�H� �*A1�{v���V�p����+���t��wa8�+R��w��&�b��i+�4������Ta����LmI��W��E��Xo��$�$���^��Ղ1��,
�lܾA��ф�cZ�R��J�_RSP3�ҹ���xF�*��:x�x�B�k����<�sBAC�yuŝD��M!Zq��G��73�@>��`P���Oi��������oT%#! #�z�P<�zx&�U�W��K��
I�Lɟk�H�E���bQ9�w�u]fS�ww��v0w�'8�/|#���jZ�)~�Ƣ͔Ԍ�u:(Hw�@��+�o��i�i)���������d��"�1&?�	�R]^�����<��.jLY�8hZ�-��$�����t�P��}M�pD�e_G��#2J��xYn˯3F�з/C��c2��!+c�ˊ��\�1��q$���Zc�%G&����q�9 <���ht?o��E�Fq�P��A�74��w�A�fX��m�I�-��9R��᜖��fd=���!H5������7�ŉ@��0�,�� ���R�)k�><�T�=�[EVD����ڐ���/��J|�%pʧ��y��$�=Rb��tR���~��?�ۚJ_Z�� ��w�.����������zD_��?Aښ�y�V��'��e��8H�:�,AݮL<�F�(���SH�SzJ<��ˏ:�����UX2� ���'5X��aGb�8R=K@�Gm��]�#J٣����x��/�&�d���X���W���@�Pk�%cؠ	c�QFI�u�D��T*s66>A�T�C%_&�f3щ�c����x���Gy��0T��&S[l�R��m�ek��1Qҁ

{��i������M��E�T�����:�2"sy)뿕5���D�⏅Y��O��r���hM��x��;�N���0�E=�6�����&����:~�p���+��`�M�"�U����F���?�{�R����}����1�3��
T��z��M�[&`���KQ�,d�6'�=���,�pxw�`��0�\�B�L������<�Kv�!\-]��n�cuqN޸)x{e��5E�D��-�i���9S��L��8̝��xS���Q�-�m�`Uv�9�ߪB`m�?��_�{/IoO6֎�lђ碬TJץW�����g�c���
� hi9ܨE�>{X/3�*}s�j�vB�B<�c޽xե_G�a8����
3Uʰ7ٟ�)hǚj^�7�N\%$�ct���9Q�7���t�iL��-ɨ��L� �-rb
�ץ�dJ���dv�%�3W��^b5����������$f���ڋo���Xo��@
*�l�E���;��ݜp�1FA[kV���nt9,g��-��c����6�M�c,^I*5r���C�M���q3e�D�UB`���le?r*_�П��%�f~��M}�C��qm��o~�AD�'+B�9����+FL�ĩ��D0g\��m�<��:�J�!�K�!k��˲2���Wu�\�T}\`�����1�Fȑ�5�JHM^����R�z�������RS�-�p�$\榈c�~_Z�?�9����&� ��#j��'Z���4�#�$qN;,���ш	�"��q�<6P�	����#]�����=��~��:骣��b�GC�}����^�t2����%ؗ�VG��z��-�4!a�H�Hܬ�N:L��\��E��-��@��_�~��%��L@t��=(�7�]��u&�&J`<�[ƽ��ַ�Zc�%���R��_ ����>n{o+!����&�K�'��W�j��6�z �
�����x}��%�;�tմܧ�s͔"
�?�z`V���{�ᅡ�.}]���/��=_�")���qץ!����[�EN�W4;����ۣ �]�)���N>�E�Zd��ȥ�n�v�=ao#wT
����'~��ڶ��7�ܵ�0�>Ghav�����d��%�H . 茫Eq�,�5�A*��=���C���UX��1���s؊}Kb���?���##E�b��'�R�#AK�$A�-Һ�+��� �-Q<pz2�����<N�`���A�����t�U}pxz��G���c���H��z�ѝ/,���K{��0�ڛ��A��̖ɗNR��4��5p�2����Y#нL�9p���T�R`����5�l��!�������{�UA�%c����?�'C�I�5�0�bzC�s>W����C3�ƌ�]��Ɗ-Uº:G�nxA0\s�oGmi�߬]��B!��x�m%��o�oo:FٞKx�3Pcā���S8����z:�Uh+TztMS���U�� c3!��,~�	���ԀpP<��^����!���3��P��-�+v�Y�1���y�v�W�
�<�E�0�ZBx��g�����=ʳh'0����4d�#�%�^�.�n8B`w�"Z�������D�̑&|�yY���'���	��W��iP x�'L��|P�% ,�p�e�,s�w�S��S��HBA;�} � �I�����1`�yQ��:��m�AcaC�# %/:ů;�&oѺ*�K��4�:�4���A���Wŀ�q'Ry�������1��30>9Տ���}�[���o~�e6���
DHytHCX�3�I�Kt��ӝ�5f��"d�V�Gӈ"��+"L����	��W�h��y��#Ra��L��%��=��F̸7a	#�P���Ѣ�`U~�{v��ЛN�hO��98��ߖ����o���Ϋ�+�ݥ�pcqo��Ӳ��v�\�ϡ#��D�y�G~,�4�[�$��r=B9푡.����x>QjJlI����<ىJ����u#v(m�i5O�si�v�J"oц�pZ
��ak���φ�x��ܕ�e��*��tڡ�8���Ҏ�F&aL͍����`�ʉZϾ���D�4��̅��`:Ӓ:C�0����6YF����laj�;��d�h����#2���{���� �#�������e� ��(�L���By�S���F���p�DE�A�4���0���	������y�g�i��I�����vѐ��2#1��H��{ꠀ��U�Jm#�A�����uj/�H�h��%3����B��3��8
����N��t�?\37��Z�DDD��4.e��Q������[aӅ��X�熁��^=ǈ�g��cз�@��z��r�)|;���U���R1�Ny��t ؜���K=\OK��ىb�*#�Q�خ� lQ���pv�4q���7��d���x�E�y\f�k���j�A���n�����	�Ј6��<������RZ͝� %w�K)椴��mݢ|��;�l��@�DLE�$�B� ���&�k��T�fYElAToJVB�lf?�X=Y+�^��0eE�Kl�"�L�S�F�j�����Y�a�޲:.�
����<�o�D��큓�N�B;���XX�s���6�����$>���nv���ظA�L�NH�R�ZP�p�h2]������c��8��	Ú�A��|��3�?MW,ǵ�/X������^�+�<�o���2�I����&�r���x��U�e@��Vl�C_Q������K=�Q�Y�j��\���� �5aQ!�A��A��4�9oŤt��3�PVLr3�H��Vg��'��z˨��*k�^���Ɣ|	�k�_����J���i^l�8�p��ˣ�M>i��0gK��Y#8�C��ٔ߷�Eu����?!'�J1�dEq3xho��Q�~�EQڼ;�%���솈����/��jgN$��8f��+������G7�NӘ�Q+�gsLj5���(~�S4�k�n�5^6Q��wO�K,��A�*�6U%�tb�Z	�
�*f����}N8����mLz(D������]]t�6�y�'&�
�H��|����\_��%"�5L|�ϿN-C���3:���7ǽ+�+���
��Sӟ�(� �ץA������vI�d�-9u������Ys���N�2W�C�	�Sp��ehK�;?�6�0�c��X&��W6�@�3�EeA�OmQG��E87o�7�c������A,��b�G3�jÕ!����w�c+0eQT$.�g�H�(��)ћ�& �F��h�'��@O���)x�k`>��=�>�tM�<��~:�c�5T��pcc�tu q�ބ��m����YmW�#׽2��:�C��Ժ) ;���]�?W;�֐�������y*������Ч�X�QFaԻ9ae>"�Pgujba��܋-��ǀ���r륉>f#��c��n�}�M��A�m��Ж!ncc=�p\�8�����-���n"����̮j~B��utJV�z�$z���%�߹X�����zdV� �jƦP:�O^6۟�<P@Vd2�=.?@����wA��{�����bu�B�3^lc�<�4�{�n��*��q�0{��.���}S�86�#,�:���Z[=9�R�p�W�3it���dzS�z*�451�x
:��v��?ΰ�A��\>zX�ޚ�B�!�5^�;�ZtW*� �C����7~إ|ud9(8q�l`��+�wէ�Q:7����:񍩍;[�=6�d)�K�_���]&Y=��L	� sT��s�O!f��'���O�)� "���s��G��m�O��hL�|E�	�#�4��Zu��I�����I�J-o����+�	�ڎ1�J�Z�J���Ar�g_XZM?��R��W�_ʨ�+�G�\¡ph���)y���s^*���z��= ���v���m�d�LK����Y��{v�����	I)W���X����L�q��j��̤l���4��]K�	��0���u�+<��R�B%IU����/�ؕR/<^�D<�K��u�b� �
��8gLE�������Év;��2�K�ޛb���H=����$��K�{��8�+"���?��*���Nh�t��+ ��5�*�^�hAS��0w����d<>���r`�1�74E���'��~�I�6��^�In��ך�J�TR��Cv�\>����t�k?�:��5�럅'�QSfK ����IUN� �j)��t�&}�I���~����]��R..4Ev�����Pb�?�z��zыX�1�Z� �[��1
�����;.���y�Y�	����^Z��n�8{�Ϟ�����CN��h���Fx�S`���M0T�q�Y-�Ƥsc�vd�B�� �<]�e^�d�Xk1}­�(�ٲ~�G��+��{�\����K�'ǐ�K���I�k�p>�^p-ZV�ٹ��\����F_b�$G§��ٳy݀�aJ@S�����n�9��"w+���/ZU��6������)i�[�PQa`~{�R ��eܣ/��q��E�	�2�(*W2N�Ġ�������O��[#���^_�~��ս4��2K���$��b���hI� �!⽒~$Jl�<#�d�c-��c�Cy�nx�ԌZ���5�
��I���;×М���.2����(KSA�*�5�sӼ:�N)@�zZxtfb�>�T@����ޥ��bE�B>�:Iء;�㾳�8��u�3�fF-��*��(����w_Ȁ�7=7+4;���մ^L] yh$�NK�S�$,K!��(0�}�>O9�R*�������D1$��ќaIjf��-�	z��{��틜�Fǳ3�߽�򬕮ߓ���>���ÕI�n��V_��դ�C&Y�Q�uٗ��y�
X� ��*���ѣ�?�u�C��),޾�����޳�(�F_����=o^�����7Ά&��s$��K��N!�:Ew���n��S��y��%���Jd/��Q� �hӶ�؍�Z��v YM?$bIb�\v��a��N���Vk-)�{]r-��Ҷ�ָ�;Ҫi'jV�lS����P�0�.�����.��Q8���2�ߎ7�ny�w�m�|T��3������� ̖�)<��]�/V�z{:�1�҅�`^U�I��T���1����|��=���+dʅ�3���f���P,�bQ�$�fŭ���:+g����v �P��U8�
���l��p���~{-}����k��V(����C���MQ�'5��c����8�����2�v[����Uk��2��*D2�M1a�v\~q\)�,6`2���0��3���Kn/�A�o�`  +��|�A� `*�:����	��W�Z������ F�6f��'G��>��M
�����9�K�ܣ�5�i\��GV�
���ex�^ �'�������v\�N#VFx3Xo;o��*��].�Ƈ��hu�|Q�z�.�,�?~#T�C�]�1%�]�|�g����	��JK��:�~"F���?.�#)n�^*��^����?}��������_�6�=��DY���{���As/-��?��F�=9n��6�����y���}��0ٳ!l�ՆFǫ��]I�O�����;4��v��=�6X7B:�TE S�d��e�2}_e�,�������[�� ��mm�C`��ϰ05��O���t
*;�f�&�-�3Q-��C�y:˿CS�A�!.�f6(���ѿ ��0Ԣ�,>�֠�7JK6'����_�Xr�, �� �,}G!�ҳ�@�g�v�����p���=�%X��}ѫ��'N�.��|a��h�.M@u,�-���njmcpܺ]=A����H�H˩�$Aîo$�����?���X�|�����1�Wx�GR�y׉%��2��u��]=�N�bF���5h�Ӑ���}̧����s�@�{��a�[{��~J
Y�3��Zɂ�^K�漆��z^��O�T��,���`�E��n�dei�|�}��Uy+�7�`�-ͦ�z:�]�k	$YG�Wm�����O��)�r�Iw������[\����_�96GB@��Ӽ�"��������&�R�k�Uq�_'v�������L������:��:��h�_j�/^CN�u�$�8�"m_sb.U�;zT�S�/j��3�a�1� ���><����� ��������8oG<׿���q{���g��niSI�\���/7[`��\5{Ϲ�&=�?�?��h�"S2S*����_	�/��IV]6$����φ���4�尌��~����
��*�Qu�_V>��t�2�8͎�����ub����aO�s�)�#ю�!l,��_���_��p͜�h��^������^��V35a��	���Rx�j�8E�?5��os��6&#�>���U����,;�׳��m���7�l#x2�A�ƪ�>�E�\ƨHS��2���p�58�)!����e�� ����2T�_ԍM�(�9ʋ�`؄��@��񑦠����f���1�n�����A4���sRꮒ<����ԓW�C����;���\X8��Dx)d���-��O�*��]ԩx�z�e�,e���qW�oP���MʯH�v�f5Gb�fP����.+JF�-ۚqw2�՝�f��:�cK_���oF��+XQ����#�Ϥp�b���>�b<���,,y9�n_�>
)�92����
�h��d-�JX\ۄ[��|�g�I�&soYy�:Gh\v����+:9�9}}
�τ�7�/�g��W��.�節/���J4>%�������FeÆ�D[(C>a�VY�rr��6`�h7џz�0���W�n6���� %���?O�Ͳk?߶�mM42��HЯG��2]�>�))�uS�;�Ü�]����B�;�b!缑�?[V��CD9��}���e??�j�Bwj����ּD��3�G�0[֣����� 6� ��<+RBg#�?��}l���11t��I�J��dr�mCCw��$%A)yP�������
hz���O�K�f�0�OP*�Ly�����/�M.���x�1���t��1�~|P [|1�I�\ w������TyO��N�\ ��g�@t��rFH�n}=�\T	����Hyu�&��f������YN!%���{t,��1���G#��[��Ё��>�B}D��5���-j7�x��ũ��Wu��.,YP�*�	�F�(��a#�3��{�u^,A75\NE�Lu�S���o-���,K�L拵�'�j}�ݐ;��y��q\Ei׭n�K�d�?Vhш��">�w�D���&m�9#p L��l� �Ǭ�YI������!���ɍ2��FR��*D̘uߏJ�l�ۜ�=Ӻ>y`���k�햆��.f	����o8�d���}h=%�I�)xDY�e쌘A������\!],;A�'H��0�W�a=�tP���\Nr�!��1����F�R��"�Aàʜ�iJs5�1�^-�r�Jy�n�r�Ϯ��1B�pl��QQk���M���'���>F/��1��Ue��v�ʤ���4��[q����a��l�����]z�u�7�^O�\�(d<���4Ք]���ұ.��j�/\{fa��A��5��B�""Df��n���،��N��*�s�O$�����4 ���vXD�(}���jS�c���CX2�VĠʉOr�Q2����=)tJi�hxٹ���hL,���O>��y��zW�5��͒� p���`~<����4��+pq�ϯ��q�ѽ1P�v�&IU�7���v��z��3+H�o�.�,�9�l�Y�xҽ�R+�ސ�����˄�ه�@?w��}+�C��M�3���V�8<��x�� T�Mr���X%�	'�[DG!S���R�\���۷rE����I51$�㎇��ѕ6Lh��z������uf=oUl$N��L��jw��1�W|d~t׬s�U��R�,6yeh�.E��%��Q^��Y,��V���"�v�;_���x,��
6,����ĸ��zТ�;��le�H���Z�T���H�՟QI��qIWT\���ޔt��`��*9}9�?��a�b����P��i(C��}��a^o"���	��ê��U��R�6|�\�5;u�w���O�0Tt���:D���b-!��f3�I������9!�m_�[�U��]������W�?H���2�~��a�����s[T���G�@�	�f�L�$�ɝܙE5c���T�4ے�XeF��p�C����!oH,2�����*xg�f��X��Evfݬr̺�`L��{v��H׶��"m'����$v�֞�*&��x���21p�kǡ����(+B�]���V�\� �ߥZ�c�M��:�9�a|�x/�Eh�{�T?3�N�}���moͧ�H�T��η_,'C�:%�z�v��]�Y/��t��ZvRq��e&���bm�^z����
Z�.}��?⁮��l�B�5�I���=�H�� f�Z�y�g��߷:Q���w �?E��)ÜV��a��\V�"�ۧ ĄP�:ˬ| dŚ�t6|l �D�ަ9��{1v�m��L�)ik��\�x��?��:h.�e� >��j2��_~�xS��9���TWԳ�U���t,���'�na҇���ג�̚�,;Ο?a��U}�]���C�n��`>����z~i��ve7�3�Ez����k�/���G�0��!�����
��ςNN|���h@�DE�t��Dv���(|���g3��$0ϲt"�s*���@v3��s] S�Pe�5�h��"n�(�Q4*���Fi�����o�m�aد�J��\)ɢ��\ur�|h�n��-Fh��y��x�=�4pd{: ,�_X)�b�,�y��=�_���|3چ����P����?��`"�9հ�����=���ucW�A��r����3hjoK��V		�^�C�R%�]�.�8�E����q�>���=�����d��)j��a�tp5�F���m)��O:���_��b��o�[:��S�t����`X=2JJ�䷠w���{?y��:�2৖�
#�Z��-s�`l��W�<>���99�iŹN��Ԑت�=~�X��@������d�_M�B��ts�`RDk������C�y'��m\R�&�缏h��N[?u.A<��]kte�V)rI�vgy���j�f�ٻ:��S�~���
z��\�s#Z�6|��B�s�I�����o�q��-,�����Ҹdk�#�e�A�n*F�!:#�T+�/m��3��4�'��]��ј�A�kx�Y�de��Ѥ���>/��%������M`nÓ�q_��w�s.��V�� ��M~���,�~�۪g�	7�=�F�z���Bc=�+9�gATFI~o���Y<TU��XO�5��;�6H
�&q�)g��&��û�]$��U_.��́��'�gc����X	���Q!Muy�����4��d��2;ɭ���,�����9ـ�a�����a�L^�6)�͆���\�m�����Ă�~����x}��,��P��������4���b-�d�	��i�U��C?�vލ���?���jy��|��3}-i�c�I2|��^j|��"&��U���LO��> 2^�M�C�,,8����$8���}�T(�bγ2:9�V Z�����a��/�MB�+Luo]?���,��N~��RV@�������p�<�h�34L��j"���Yk!���=]�ʵ'�H�����g��U�+z��K�E5��A��\B���d��S�S	��9����]�=��s����]�w���*2��"X&���/~�[��?N��g�5��r�=%�Ҍ�5�jp&��.�����~��qHj��MjH�QT�X�oGg&��2a���	�>˟s��uM���ӽ|�}_2���6��ը�"8�Σ�9$1�6�H�g5���}�iuյ�J �Q��9G�᎟x�kǾ�I�IX�R[�]�x1�&�N�
>�s�h�3��]`���,��(�ޕEv�����s��*s�3�GQ4sov!�ʟ&�R�샅6{�2}�v�d�K��pyH���g�Q���Y���������:�t�9�Lx(�V�J��� ����y�!��G�c�e����9�<�Y�p���$���et�=��0�S�2K��N�\���x���0��6�������F;`���x�U�(���+g,��Q"`+�������׵����6���!^(�����YYp�NA�6�=�>`G�k���:o~��ё�_��jI1�(q 0񃢒��P�*d��^a ��4M��|���A֣�L�Σ�N@�K=t��m�2K�}p��CA?���MY95���q�
6(L��^����r�ߞ4nG	�Ë��׀WR����*FA �Y�����}S����тO�c�I��y�ʷ8���$�	���1T��䦇Z[��A�߅�`���Bb>�j�3���������^3�vX^#�Hg�k��N�ޔ���3.�]�
6v����̐��,6����s?�2�f�L"�d -�s !��4M+r���S׎���M[��e��}<�U�h�1z%�R�ك�����i�Kj1TJ��*�є����,Y��S��a׈����\(	et��Q���␻��B�r�2�\.R�6@WMo���<��]vaq�=V�ʹD�����X��
�nn��"ʹ�	}.�����sT�i�&*�@�<.�ꗜ��Rr.�XK�Iy�l@$�;���������8|Dj�ʉ~��eلG�!�#����@�5?� �{�C]i�R�	ɋ8؀|�L��BU��bL�r���Y��	�7���h�k"�bM-���zsu"w���T�oq�a��8���f�\%J��ǿ܄�����L��)u��:����-�
_�9���9����ő��'Jm/̚���c�0?��H��f�z������`�8T�c-2T�A�}��9��	�idZ��o/���Mt�<�y|F�$����
�F�i���X����3��<�)��=;�!.��zS�_q3|�Q�7mכ&]v
�7T�R��XFP֞://�[m)�9*���]A�G�Y�k�[T.�-A�b���IH��]��z�����"�fq��?��6� ۷�c���,����*�0�k���x��"+��hg�����m�lJ��`�U�.�4Xud�I�<�k�W�ak�-��C��=u���Z����s���\[��0<T(�h
��ƈ0ݡ�^�S$9���7��C��l(F��G��Ct�y �^�-��׍��_���j��w%9<T���?\m�� �D��̉4��5��������g~�^u��i20�|r<H<����؜"��!�����]�� ��ZH�ь3Tw#w-��^����]�A�ϸ�B�u��ޯU�o,�4�MY߈kq�"+���\;@Ȱ�ƌ K����Ei��jpBu*��'��[gBW�:��H�I��x�.����E�tw��'#۽�����)����hi�\��7���$~�h9��i�m�@�����Qe&dhfAh�Z���gп�#b�D�ݾg�N&Ժڿ׻n7^#�lB� ���ί��s~xSXqe&R҉˷:� ��,�q�����/ҟ�D;\Q�#��hxL��B�&R���b����#�}^Q�q��[��w�&��N�o��3Gn��5�O+��YG^����a�Ժm	̪�6���;]�4�����!O�f,��O3w����fS�L�ܳ'���}���� �)lE��b=�ϒA8ő���Ӱ�RHj?��@A|&�I{����n|@091���Q}��vw'�uN���q5n�09Tsz��N�)�L����A�i�g{�5+X\����������Aٴ�`��CZʣ	c6'�rAX��02�Pd�w���O,�<8c!�HZeW���<U�km�D�Re�0I T�b[4��ѕ�i�����2D�H���0�_�/���ծ`������_S}���,�vU��.[����|�'�������n���i�O�Z�9ɠ�a��e�	��v:�&2ͷ�8�e�V�2Ǳ"�`X ��mz����5�C���46pֹ�몇	�i�g�?C��<Q7@j�d7O��M{���B��L. %�d�EE���L�D 7uMP(koQ���^⍩�L� 	�d՛��y"��ڸ��*m҅M"(�\�cW��A���D�l�0�~�>�s
T���:?����v���@_`,�3�� Am���
�l�ܱW4��pZ46�^!X>֢*����l�3�`����* &�1ER/�	>E#��g3iY���=1�<*�arҩ&0�����S���3�)3�~�@�_�p;BJr�ްN����W|sҚ1�6�� 2��@�u��"#���K�T	���#ڼ/RlάCQ��s�m �!��9,�5�7���!�x��ԗ�>���R�@�W��~f���)e@���ܶ�O��л6�|h�� 	����Up��\����rO����a
���SBWjI@14VL�9��Y���I� Tz�$Q"C��ܫm(O� �~@��-������k�B�(���,��XR5�m.y�
T�!ӵ9-B�mД�G����_��CP�|酻꼙�\ �Y�e�X�lV��L[� ����1�t8-�b�ӟ/W#�k��K5c�8Z��"?M��h�&�,6z�ʡ��j.W�G�ho�S����?�������G�Y�	�?a�l���lL.IP����M\#����$M(������%Q��P>Y����9�&���L��xm��*�-��F�ЏHl�~ZY3�5��jC#���%ai��L��]�;u����ڔT�!oBö�ۛ;>�5�y�D���r�[r �����h�.m�#t=��C�JL(:㡓�rNl�V��XSX!<ӭC��'�{m�xl�+����j~�ڔK��o�ã{�y�tii�:��sAw���Kv;d����.��I�\pؒ�h
�����ɼ�G�ZP~7���x1NL�k���h�ш�g��)��v����dM4�wPY�9lJ��֌���՟)����j0>r���� ��6B-H5��L��m�l�J^�J�1d�Vab�(6zE,�$�Ѭ��x����?��7���y5*k��ɔ�D����Y�*��!_����DZ1]K��WIbCx�������J6��0V�%���Z^��pM�&,�r~�a3���2��Sg�f(H��|�bL��xf
k1�Ru�F�e�YC�_��A ��AB�_�CZn4�r"b�F�o^�.i���5�ʑ�R������K��� v�K|�[�n"*�q�b>n��,���e���`n?O
7�F�(ٖ*X���'�w�/�10&:7���x�,V&�/Nz�WL)�l��%2��)���Š����c�KO����9$��V�0�di���z�G&�B�)7��J��}C�rv�X�w6����_�CX�D���k4
��I�葕qC0M�tT�'Ҹ��7lo:��3���b��z׊��3I�܋����xo`��"�;�j�6 ಃ��j �AL!%��CXr\M�EX_iKW����7&��>x_�����j���LȔ�|P24���3�>�J�i5�.�~�K�+[�L����g�FU���:/��HS:�`c��X��ԻZ��(�bs2�!� ]���-��d['$�a�ܗ�X��_W��>�[�6o��8�x�u ^�}:q�59�@��t`/Ԣ�\��g���.�7L��C���d��#���8��[�(/R9{W���$IQ�U_��j#���@d�݉��mG[��Sf��	�\t��A ��R�¥�7*�
��J���V�nsMO�^Ln}vjc���>@�tP��L�Œu~���@��'Ѳ�#U����9�6�����&�E}�G� seF�=��4�=z�Bt��W�/�Gbܟ}�w>�fi�Q���+̧�^�K�JV������hx���-0�u%�) )�	^$뗻5�ik�K,��&�A�Z��H��e�Mi&+���"�҂�*5���w�τ�OB.�k��o�.�fa3�7o�N��L���`�ck?~aE!@A"J��U�;SU�l+�z����Z��V��T8�Z5/y}[MU�u�2{�JUq`���y�,{�����%�qk{	�����{}�T��S��r��i�\��~z�Xmb��?�:��ʦ+�9�D�ޚ<b�0��I��i�e`(r�;I���|d��;��X ]np����L�\Z�b�_ۚ�qQ��g�����=�c>�R_D�Nir���4�@���/o�����*%��Z��iJ�b��G��n�.�^_��LqRq�x���C)<�s��'s(4�:��Q���5`�+l��jpA���P]�5����[ϊA�'���mfoM�"�-��Y��ϱ�ۜ�W��L��0�C~�t=
���b�Gv{U-Ra������3���4���?�36�(2xn5Z�k��h�398�� ���3��"
d*��'��K���C^T7�ru"\�r�A�Ff����)��1�!hU���[V��M����1��
��u���:��Q�q}�|��g�� �0��Ըċ�J������Hg\�S��ҹ��E����(U�^q�?k��$��yҲ*�SY�"�2"j��������Fb���c�G�������2������9@&���Aj��������;sK���z^��J"A�Ò�B��9�f���o��~�����l�u���H��$:Z��u�ț��ЫU�K����z�U�y}�Wf?;ȷ��sع�;����{x,'��2?��j&y�$�`�L�C���5���v�`��9R�u�^ȶ籸���A$�A��^Xx�oy�&��e�u����T�x��ZD�`=�7��x}7��Q����K��Y{�{%cI�<_���qϓT*C�nν�^�����^;Z2�뷄�,HE�	�{�{Z�j��Kc?Osm���|o�	J��K�Y �GX�g���D�;9��S�Cw-�`��ܠ�m��sj,"��@�~�C�<���Z������_>f�w|�!���� �v�9��	c��E\S6���|��5L��
�:�Gq���uwg|g��5�G:?y�ޜ2q`��?J+�?Ek������׊�0
u7n��6��8J�z�wv����D�|�jaRY��B۫�̣���q�9D��_�����V�f�[���/�XQs&C_\f�i�
�k{3xЊx�v�R�NR�d�@�;b�-p���r��E�̾��&����Y��g��m��TO!ar�~�2�ٯ�OQ� !2=Ǖ�mc���['("�V���\V���Q��yŦHt���v�je��ᏆT��@���THu@W�z����7��3re�{�p@�b��kP�,mf��:)ob��I����/?3.�Cn�'o���v]X�����BG؁�HG���B=��VW9���+�QKq�ϰ5Z�
����i6�����1�p�*Eb�|J^]sѻ'��+�\S�S�XAҦQ�a��&����n��;t�J,f�Ѭ����u�H�3����Fjo��X2��,�������$��=��BP�S�_�Q�+���6�������"��LW3n9GG#����;$fMSȬԘ)�d-/����ۢ�S9-�]p#w0aN� '��E�b�M�'�+�)��-�
c3�T��`+ �t�ͽ~��,����q�Ex{��#U6�.�/|�6�xٙAi�71u��AnV����dE������'�k8S�^i��K���{+P~�#�'���wrϊ�����@��7�Is�6��	UhƋ
ڿ�~eLsgW�ɀ�b���o��� ��~��=�nU[��h�֎ꃀ��"�lNWz4�=d�'28_E`)��a�6�Mޭ�N��tF�Wǻ�y"�gu�y�$h?�ܼx�ؖ��IkH�`���5'e{�����"�"5~u���z9����2�se�j_�`��я��&���9�r)d]_��X��Y=��}!�LȔ�t�i��ͻ��ܗ6��jg�$���3��[��? VH�z��}��w��^�n��}]#��
�L0@Ek!�
6����"��C]��8�ؔ�*��؝���&�#=hL�1u���̶��{��-�j��K�3�B\7���[= ɩ�b@°7)�����Ʒ
wώ~���7݊K|y�zF��(���r��A��:q#�U��.>���	���[8�r��ϔrlo��iW�V?֡=1���p�*�5�e�Pk������r'}��y�S�@hEdƝ�ﶨ��B!;�p��V!����&J�'�Q���Y%�_[�V�J�'n{n�۠����K��vl��D��}�>����>6}%�Y�)�0����F��{�����r��K(enI�r�U_���N�����H_Tm�`c�c鄢հ�HX���9W�xU�_�j��T,���kg�u�P���4�\t�\��NZ�XV~��
n��H��=R����M�� �L�5%�B��J��3��i3ݖ(<�9�/���Տ5�Xj�j���gA�K`!\���(� ���"���}���U�}��Z�`K5��t=�����3*x�:R 1
,gf>�>oi;V�~�8qɱ6��>�D��)��1>�W�8��:�.�ܗo���V���x�����^~P<j���{�e�5�W5��zW��/�_�V��κ]���#��Z��z�Lש���6tԀ���u������ÕQl��r3^��q�����d���[��x
�������ݖ��u<�*��!^g2U�] ,�]t����_&^ ��k�������^�g����t�|7Ǚv:�u͠�r2Zϝ2�ΝU{uӠX�qm���M���/����~	Ѧ:*lDw�ɥ��8=�(�X*�����!��O\�^m���EI��$>�l�XȨxU�~Q�)W6�E��!w�lFQ�X����'u��ջ����f����y�u�FH�
^ ���k�\���QQe�.�KS��(����������b�Z��pX[M�J��6�d�`�i�HD�`�򩁕'S�ͬ��x>Y
t��ݺ�� ���I^ ��$zY���VN��M'م�.�,
t�6����-�>�W�?�A�谏7�>U�������C���,�{gJR�Ӿ��h<Z]��ux���C޵?���P�)"�\��C�W��_�	��� eG�)D���C0��A��֪X �o���{��h��d7�$2��Ae-��:>d=�R���:E�c����oϛC�\C�k�������WQ��o5B��K	��>�_p��a���	f�8�&{I��[����kO�[ũ�y�{Ŝ�����?�O�w���lJ�0�Xm�3w��t��q��%r.2@*������^ٸ���,�����o^�J��7�e=P��Pp]���,#�>�n�`+�<���JǪA;���#�����&M�dv9�Dt��B��@
 8XF�{��v<��y�'0©�����6D�Q^A�g6��u�s�a�o8�Vhf��(��PEV��瀀��	\N�H�DD�޿�� �=�B�|��~��d	�v�h�/&���-�)]�s�&x�3E���C�m�+H�Y��b�)~���#j�>�!�%Tžf%�� ���ʙM!�Ǐ�Ȯ��xx�ޱ�oS�Ha�sD�~X8N�~kˈ�M�y��)��'m��ln��)t_��1\��(�	KG�2Ӳ��(�w��40R��&-l���#'�ܪ0��^a����EA���q�*z�ف��r�^{۵�L�T�>q~st����M�7�����$�J����M&&�~3*Be���NH�7B��![����N�q7�˩41��\�ﲅ7��;�������r<>S��l�w�]*mf[�S&Xp��i���[���4�K���~=����[�H�l�L\�P�
�Q��#�]����3� � � G���tg��jVM�E;dB_���R3��?]����߮��Y��B�׻����*]1���|*�Yv���aje�	��b��»Y�����t�{�J�g����k�����|T5����t����Y�{(Q��[�H�ԣ8�R���~˦�mm>���7��t
����]�M�hs&)��-Q��8��3o�^����vf���}����>�L����	�)@*��_eL�̱�6[n�TV�����,ޑ��V�9�u:.���1��8�p-��n���E4sf�1��]3?���9�.,��;��&�S`���C�dx��m,^R��Y���p�W������2}���"y����<�K/j�֝�C'��Y��E�h}=��f銥�÷%]�yow�$�8Dbyqͩ�v5�J%�19� Y�[H�u��DX����;�V=�J��w��泒\8O%O�&`��� ���r����@ɔ7<!�L4�1���b����� `6[Z�B���C�br2�2%�`L`9b�5�L��PJ���qXʚ�֩G�nPP��|����eC���Z�,�I]�pi�R�_{�Ȏ�Z�g7��b��F�>+ƅ�8NF0��SJz�m�c�@A���a�C)�q���JG{��frȘ�l�b��O{�f`YG�¶��Ā�ݒ',�N:�!��b	]n�Q���e�L-4�,�h�����}}�����;Z[�Dֽ��#�N���F����}``�$9=]Oi�ػ���I�
7a����c:Q!��\��-���ٹ!,۴�I�Z2/�%��I������Q���3s��I�{��I���)�m���� %#N/�u��C�V(f�m��0��3xJO�������Gv�@���~���zL_>�M�����Z=����m�3�>H����_�*]0"��~вxʯ��p�9�57�f�O`���	�{���:/�Ǖ�z&�H���Cv�{��i<ݵ�����Y�*�H��?�J��v?N��M,.�-dq������1đ�6�د���c�ޏ㑌�p��<�⨐���/�
����C��Y)���i@�7=���?��ړ�i�@�PI4�r����Yü�7s.�w��$,�E�
C0A��"Zܟ�"I�d@��� ��Ŝ���A\I��1�]c�32�Z�k	��'�z?~c[<;�!g��F3�����o�4�DQ�;�w�5������ � �<�k��d�zv}2۟�1ŻO��Þ�˿ڦ�~#5�c0��0�!�-I�!;�=��&�8�>Q��'��Ԝ�"�S�)1«t�� ��q�1���7�;�d��T�G��#��/�q~�� Cz0�Z:M�s�����'�?nk5�B��Zd=�6�"�$����9	q�s0jYLE��(y�x�䡫�b<+�p�0����Q<���^_�͏3���N(z�� ��_�c�����uݠ���Wkx!p�-�|r��mI׳�����d���9^$��� ����8�q=��ߐx �Å��d� r��$���g��@��y0�.~��5G�������gU�q��� �����\�X�6���
L�����SS��Q�0<t0���F����|�� ��Gӭ�����P��ho���
�ĦM�\ �L�s��:7��Y-:���D�¥�kK�V]���i=���>�z+~�8Wl�����:'������=A�s��x���bCϠ/�ګ�uɭ��\�_����M\�=�����=E&A^̯֋��96P�
�m��:��7c:Ah5��i�B�oa���
����i)*��uy-阙�"�K��_�g[��L�]�.�0ϩ�Z�*�������\�"��Hj�:���Qh����ʕ�c�yŧگ��8�G�fmZd�(�(Oߤ��2��Q�+bC�����}����᷅�`IǞ]�xbǤ�z�0�h�X"	���"�r�	�p�A�ٸ�B>��4H[.�uY:�}6q���c��rO��$֦*1A�8�|�}oa&��)��k#Ap�k#[���Gm�b��b������~���h�lѿ�͍]�~�+_��Z�ck�5f���Z
�DI��YK�x!��{KRc�S]�f0�.25\oz������b���^����g�`g���4�� ��ƾK�Sx\V����h��rk�:Qz����~�ot�ח�m7���9 Z~@db=:�(_��!�(a�(žu����W��%��}Zr�F�p��i�Q�\}qקԓ��U�s���BǤF���=�W�.Iq�P���nqY?��#Z�����i�!+����h�����>ȼ��M̍�Q6~��`Y��s���"�[����C_(K�5�aV�W���@���]D��Ǹ^����\�D8 }.�͒��&4�QLl1?��SCw��z���G��N1fP�ś�ͼ�:F�s9փL�W�vJ|�B�m����~�n)��<"�Dp�Ե[���W87\§]��!~�`I��7A�����i�5l�5C)ЌI��<x.Q�:?�(���ɓ6j�[��:LO)罚��Q,쵃�;�$ӘO�p2!��O;G]wD��A}�i��
g�=�aW��P\"D�A~M�ۡ/�����>�5`��O,��������#��Ky�����wN���`=}q���@��п�*m��!����8��n�̈́K���s��I��E 5�ƚR7��_ ���'�օ�Oмt�:G���X2�� 
��[\Y�.�e�d���3h�7�@�e�RM3��z�iYeJ���������|M6���̝�M��7��܁��7�����>�-Z<G%+�`���EN��Z"�-n��+�fb�o~���'5�
���^'��� ������H��XQ��
lx��}������l�Q�)A��
�viH�(i�.��}p��z+�a��K܌��ćx�'���u�������-5��*d^�#Y����L�9H��U?�^��Kg�G7����� ���-e�=+ɺ=��.��K�ϱ�b�Nt�N� �N��B��S���;N.kLs#n	C 
R]#������P���a��)��'_o�[�+{��L��0��<n�Iՙi��;0g_�иJ��mq��-$�^���ʬ�O��@��[�uy�./s�l��CB�
!�����{�ǥ��Q,�A�K�uf��wG+�!V�p�s�t��#)V�����8���<�B�r&'����P��qa�p��M���zS�a��ܜ��)ˆ.��iF[G�ʒ�H����l�49q�pШo��$�[~-��~��&��UH���UP�[�ܻWq\���$�W[qg�g���xՐG����N0��	ݧ��T��$7.�ޚ�I^k��k�5nD���$�����@��!����~���̰��+��C���!Y��z#ib��2k\nQo��,�G�b�M=���� W&P�Id�?�>��# T��8����:���=Rh�G��V港U�r)�gxB���*�g��J��ڐ�:�P�r�w?8E4�v0���2]������{u���x��.����sQ�H\ؚB3Г
ZB�D�O��;�8�2\�����H��L󻹮�߅/�	S���8�L�Fn/Y�%=���:�UT���0Ġ�EdD|�jcRp��A��� �Bjӑ�j!�����S�D�T��1�;�N]� "H��5��2���2�.�%�\�|b�E����QQ����;��,au�ýbhD��Aý��Ƶg �Y�5��N�8��ا���G�:)���Ƭ�[�9:(�&D?������ɶK��� �(�0����H��z�Y��/�5��,Q�+��iS���pM	�	գI%�1Ճ"A����ok\"h���2�r�	�jm�V(�vl�Q
����)5�R�_r�G߬�/�.�o=K�Z�Y�J,&�޼�vka7�O6�(�/����kϼ�d#��u
��4|O�^ss^��+b?�FET��㭮�o�+(��$Le��MR/��X�NѮx��n�a�8EǑ�T�]�{MA�@@�j�Rx:f�ˇuk;1_="�)Jg���D`�ɶ�87J����D��.�r4Q�e�{z������ln��P'E��M	��_I3dNF|�V��e/.5�w��_~�B����=L�V��w4�5(/*�}Xy�!'�K�Y��-��z\M��RZG�-��ɫ�-�j�g�)�zZ%�KuDN���e?	����9��ER�J��XQz���P�Z6������o>�&QW�Y���d�nUkjG��|�nc{�;���g�*��:����DH@�{I�g��\f��B%@!��lª��U5���Lٝ{F!�x��M`ּ9���D��?@�Q%�e�B�&��(W	��|'����|Ǒ�/� Y�'I��%(N�9��M�"b����!B!ӽ2����C KFݲ��@���~��p��]���l���'1����i���Z���v9ah�nnOj]��?��o+���^���ъg�W��g`2�f�g'��ЄZ��h���g��YÇ^[����u���+RXr��ل�Q�.����.J�Ng���dt��Ҡ�Jn�����.;�xj{�\`J|�m|{����V��� �J�f~1<�~�8q7%�n/�[3IͶ8cd�.���+ɜ�yE~�zR�$d#6�h�F|<��D����{:%^=��ô��:P_Ž=]� bX�Nm^�F�Z W"6��p�ؿe���rP�/�Q~�j#��.厌��e��YNp�_��� *"�K�us��wc槨�S㇡��P��+Z�}��|'hK�9U��-������!���^~�R������h�i�QHl:ON=5���9��&�CXG�^Y.7�$m}��~5������7mJ8���L,�2�>Tc�qƈ�z6�f(��=,��9}���!��h�xy�KP����zZ�h�`��v���5�
���&�=�v]�*�3��*�j,�9z7WR����!X���}̬�Z_�����iiZ�[c�����&8�Ǿ��))�Wk)"nT-n�v���X�ϊ֜_BH��`(���v���xh[ }��<���Lx�Q�cS�s�:�)_���R��r��_0՟X�؂����q�Ś�T�u�����B�z�ʠ��`�����A2�Zٻ,u{F��>��Dd�A~-��_�rW|ܙI^� k^��%���k����lS�O�UtI�9B�?�zG)P�C�iC"�tF�1!�SN�>.�S�ȝ|	����8�KF>Gϫ�o��Yx�J�mn�:�Qm��E��@�m��}J��m� �L��!��SY�����~9oǾ[���sz_�(*�}�R�v�1�-���N�5*����s(������þ�M�+p��#�L6��R�N*�@j��3"��}1�)\|e�l*&�!{
�&�~� �*�-��Jt$�L �G��F$!k�╢��?0��^�l��������O3G�m��.��oh��Q�%C5���dEBF���olP�:>*�� б���2:w�L�Wx�us��	ԭV$~&��L��
"w��n�'d�^�iDQw�S�8�5H`�U{G���bJ=�+rc��O� ��RYغњp�@>!�!o� �[�����FZ��A*2%P�y_"���N{��r�e�4�����߫� ����4"#f���A�d
 =A:X�?��m
:� ����kn>0����*���619Wi������J���*&���)۱Q�.�L�ѿ�w~��Ck��1q����vEZ͊����6 =��S�$�ng�����ܿ�{��vI�3�k� H�Jp�2�$(�7�Y����6Kr-�?���Ȗh��3I@�zV��ؘ\�_�=�F;�!ד�̻[��R�(�1K ���V���QZyh*�����n������/�vd!U	��Uo���M��!q`t�
�Ɂ��Ҷ��<�JW;��{'���E��C1Z⬡%Rij���O��j������<�������EKֈ�ʖ��h���E�M-�o����z�*�oJF�2���U����MԵ�Cـ)�Qis_�&(�j�p41>d���A�
�u�銕g_9�R�q�jӮ�����A�����CC"�)��A�<�g�^�1��hz�$-��4ʗuRx����*�M������
���ԑ��`+����>��cnʛ�䜒��1>~Уz0���HNF6�[k^���5�?�?T.�ڲ]<���Z1B�Sq��1d�d�����l�!O�ej8�s��yz%���C�����&���=s5�ʔ$;���j/�!E\�|ǎ�0\}���'jk01ʀ��M��g V��\%S�2`3���m�]~�u%=~%0�K+������W�[L��U2���f��5]�C)8���:��/\�a�bĺ0�zH�N�������s��"�1�Ej\FX��q�D1�c��F���
?�9��7�W�A3-z��t�>@���(Y&J�9����9�z?�b�J>�ʁd�N�]��r�*`�BX��$ٌ��ΨŦ7+AE����B�oa#�/]�������;�#`
�Uo^&�n�_��p�!���о���X� ]�E7�uĩ�K��9�z�;�<mr�FE4
}-�/�m��s�bcK�P��5��3�����`@���U,�!�!J�C���i1P�ٽ;;Zd�b�6��ŧkK�X�?����1T6�1�D�!�w,@���6E:θ(���.�<\�ʏ�q[���l�Y�a�3g����vr<?����{a�{P��_�K�-*��*R�)���Nt��m��b�
$m�:r!�(����[��`BB� ���p�XZ��k��N�	1"��'Ra�}+M��Xq�G��ɨ�����ݥc�̀3��Ѝ�6��C�V[[�rZG9%��A#� h�Q���}U�����z�Y��ð�yBwD|���cy�:�Y���\e�2�)�SZ������N�l��'	%��ۓ_�v�C��L���<021���@h�b~�4� �EP,�d�[�*��q�J�0dR!��!�׷YlA"�������{qQ�7 o���3~�v.�s��Et�3���A��j^l�����n�cw(�=`#� ��T'$E�t:jv�'H���"bҨ�Q�N��^�H]xo���~G��Pjv�hYj��zm����w%)�^&��āwlO�X!A��@-����v	YE[��X��0X;��� �D�y��X�C'
��ҝe� Ǻ3Eh�H(Q5�h�sė�2��콕*�J����%
^�|�� =�V�T���q�;
k���S� ]2���m�f҈l�Ϧ��ЦR��� ��L\��H��A��Q���h�_q�C�x�ܬ����������lp�7�����f��7��>M ��[��:8P����!>ih���7����wRs���j>!��\v$�-��]�=�se�(��s�-�е-{eEbr���0�/�I�#{��6�H'�i�������^%���u�e_R!fC�������9<�O"����z�
�h���ޛZ��l�� pY���-'�X���6#���ݗ�M��1^�ܸN�̶�������8Ь*E+��wW�S��+w�%SUg-,�8�����3���P�F]������{11~u��~CU-�ZH#��k�M��z�u[:�o��ZͿ�I��w_��YK�jؿ��x�R���I̽�>-���Q�K����<Ðq����bs���b$a#UT2
����S9Ze�"w��o���-��t�g�+�6�E�3�j�����0=K��;�š����A��u#�I�q�W��#���H{A�)�"��H7}ز����-�����V�� �0Z&�Ѯ%J
�t��B~� �7O��>�/Sj.��8q�H�)�PɈ��R�0��_]�TVn��z�{��,���8�چ��#`kL����ϥG��Q"�������F3�0RW�hx�<;��|�Qӣ*~0U�ߖ��b��|zv��>���x3��{E"O�"�&��������2X�+���!+�p�Y	���4����g�B�ܼ�`��ږ�<���H�C�f��`���+4:�����%������z�	�M8qۻe��0w��G���N9ϑ���v���`6OT��3%����R�F��������QJЋgsXS�x��v`�^7�a�����=�η��qbxr���	a]��=��Q	�w߶�����m�����w�Vp���t0/39h"�j!�����Z��zY�b�'w�f�>���U����!
��/b�"���w����$��}"(Қ�s�<fr]A�p���������Ռ�w�a{�L-T���f���Д�Ub#��h,w,ru��^+��ʤ4�!�23,̃���}���ҊH��D�V�C�� 6�v_�G����ZaW�����x�W�(�#���9*⩳�&��&�ZDmE*�����_��$5n +��DU�LY�� ���+��^��C���U����M�e-ٰ���5�gx�%	�.��n4'[�+q���b�E���d%׊����3}�NsG�F�g]��qK�J��?�����ba��k�o�x���3(@"=,,W�������o�&���/3?�yN��H�i������8y$�b�`�A�N���޲��9^U0��G����̪����I�Je�!G�3"�W�\�f5ۿe]�V�ı���G����,��+�e7�F�t,�<qC��1u�+=���	̪+��G*ys�̃���D��i�yƟ�#_�P�K��Y~W���{��0K+}b�,՞_�h�XE���?�T��w��� �a�*Bw
����B.r��5I<F�p��em�P�Ծ����xq�8��,��AP�[(�/9�����ڴ<^���6�<�?K6w�G��ѱ�}	���FE�M��d'}�%)Wy�O�&�;�z�4x/��rE"�b*a+�c|��RM���V�}0z�2�����N�H	W������{��H���iD��"'C	04��41�>b�C���4�f"���y��!�i�<��b�V��B]�ލ���D+K�y$��7��˖V�&�Do�l�,?-R��s���i�&���[��L�PT�"���g��Cn��3�F�6���	��ª�1'���X�g���JeZ&�g�H>�S.0�I']��X���^��zz��$W�w����lJd����(d��P=q��凪�a���$O�~�������t>�������^���Ɩ8�����!�
�5�"�� � ���"��ؒa��~C��	l������]���S¿L0�cyB�
TN�2���L&�J�`�3jp/$쭨r����.by�I_0@�CB1�T��f���P8��lp�ui��A���0Z���*��X+C��tN��%7Z����c-_|�����H�c�����mc1�動h���@	��ⷧY��R�݋�,y7r���Cch��n�ITSmգ2Ų,��F1��^¢�>PՀ�A��ы�ư�s�}#���7��L]ި(�w��]�v&Hô��9�6;.nV�A�Xi�jP824�<h1#Hm��1�ݩK;���r��`����_���O����]���>���6(��a��1h�����LS�T�P��*&/�rE�$	 ��W�<�����!�&:�����(ٶ#��jy�����!w�'�����)����]�8��˓���M�ph{���:��#|�l�A��je�Q{˒$�m���RI�	'��e��h�7=�K������M�Y�� �m�0{$�2�#=T��d;%���'��Ee�?z)G�u_:�\��_L؜�=<�Bc�ċ����/���|gT��dm��/��b]gPI�h�Kr]���p�&��e}��_0��`(�i��2I�~h�D���}�a�&w#n�eUl�`�p�C�b	JѶn�J�ݓ�yG!t�;W��H�R7��%Keo��"t񳂎ؠ�}�VZ�9�੨�቎wk�K�$�y��s��ֺF*vaӽ��
�KX�FI��!m�?��E$M%Cc���?�cg�X���Vͬ+����暤��e�P ��q�*�����zD�OY$��( )�� Ƹ��Y���KmK ��t�nZ|��L�����	��픘�L��!F48���fc���Q��`�3.~�����`��}׬S^�izB�6&��w��io<3�,D:���� *��p�@��B }\˳�^l
t��Z�Ѭ
Q�Ab� ��YwV����:(5H/�Cfv�:J�,\J'�Xa<�2�Q�s:����:��h�b��fhl�%�,��V�X�o����?Y��b2��ﴚ�Gg|���&�AY�:h��v�O��xy��[43��@�e��
�)�5&�ُ�#PP�_[=�0~qNb�zi��z�y
���{���R�M�}�m�� )&?P�ad�;`��ݕ��
��}�����k��,�@	��dm#�@z�9�m��x�_W�7b�'&�l�����,�˟��Hz%u�8RX&�����
1@:K�>v����W�F���e�.�Qc��tc�����8v��s�W�;�!&�|��'�c�/�w;�Z��c�o�6I��_���l~�A(hR�����5a �yvdc�<N�G��%ᠡ�����#LH'��& \�����1��(�mhѝ���B��et��W<׉����od�u��"�j�{pr:C�aO�m��\��?�g`Q�<�v�k���Se�����mu)`T�h��-����^���2vy�_��H��}��#�ε�o�ꗣ��d��{3(y;�j@U��|�QKbJ�����'�Dû���4^Ǖ`��?��D�����z�h���O/�'�h;;��Ǿe� � 8����险6M�i����j�����/�#Ň"�����D1~t��G&�ӥ������>dPκ\b���l��q"t�]@h�£���s��̤~�8V$��EAW��?QY�ֿ���ڴ.F �w�F�˅Q؅����������r���C�qOL��ĉ��ϲr^�����q��B~#�2�x�<!χR�O���U�������ݸ�,����}���(m2E�E�Ue��*Gev|aʴß���kb�J-&mf���r>gZ6�kp[W/�����t��;uq҅ojؚV��#u
ow������T��jQ 6��Į�w+�2����� �U����Ui�L���I>a���5v���E��fH��b���y�ճm�ޛ��vі~!�!/�z=_�7����Ҧ�^���ݥ|�ȱri�V�w;	��ٷ��H ��� d��mug���
�M�G�#���wPE�
�(Cl�X�7*��ꟊ���
��\�1�Ĵ��W����	WU�ƧFCP�H���7W�uCat TU_Y�c��������p��*�hx҈��1e�ܰ�Et��_l:�2�7�����:�pѶ�<LiF��D�17�-��8�#�K>����> �hj�[�H�a�E\�[T2TW�6�>�!º�L��F"_�>�,�P�K�9o��>�>��|�@�Ju��̩o/ow�9\mu~���(���ڝ�>�s˭t)v�Og�N'���q�n�Kj��YS�N���趘��5�AA�2j9QF�)��M`�x��ezd�P�]Ή�,W=7u��jQ�a�tJ6�wx`�MYB�G�Qp��Hef�l�NF���u����Ǧ�;X��m��!<��[3���f*�0�,/�����O=��)�[� ���H�kAS�y���bw����NG;
�E���Y@��&!a�U�#�]�������|�2�f�[)��'@J���K9l��P���c�k2D}�������<g�]������,�m�@��_��w��/�#>���z��C�_����a�M���BNr�����X��~Ә��Ԭ�p��'^����8����,}A�[c���&�'3���.�5���IJ�@�;��h��e�w#1x����,`��S3;s���xeY�p���rbW�������� �� cWԆ���:G�)�l>s�c#p)��["#1��?D��;�i��G�/�Bm�EJ��~����?2��TM�Ǯ��xW&��6zT?��� >�v�	q��Uw�&Y1���>P��}w>�����<e��nE�,։��*A�e�F3��Z~���U��� 5�5�Vt���gY�7��+D\�W3ƂB[V�K�m��.��Z������-���Xt��^hVq�̌��S����8�B��9�[���p
%� _�������7�>jYx$��<X�m�{c��PkpfA�H�����P<��J���H�5ڬ�e��F}����s�����hэ��߮��&)����V2��R�����$�1@'�in�U�e^D�7�0��.#�����k�$c�XP��f +(����S���y�L�z�o&q!���x��HD�_"�)���l�����e���`�:�p	
���;�E��EB�0|U:�U�h��dĸ4���Km�WxϨ��8�x4gw����6���$�*B�� ���� UI�]�w��.���D6�g%iӣ2�T{ޑ�f�]P�l����1�_�,-Z�����d1W��k�����w�
b�����kU�c��s+��� t�k�MO�h��dd���'<����ĥ� ,b���8��%�TJ�wGb��r�z`���#J`��7��~e2�i0��P�����R�L���Z%�0��2[	�ۅ�5 h��x����ν�S�0�_��{�W��p������$��E�/�I�|*Q�G*�����J�v�[^ /���{�Y��AaS���{�YB��xO�)&6k�$G����_��U���	��QWe����u����HϢV�fr�2B*o��!´���-خ����{@3�Z��7�ڑL�7�t�P(����"�'4$�H^M�q�+4���WE*>Xl-g�z�lۦ�'��%K�a��LX����PX\2֒�|��(f�[�g�N�`��t|��Ejͭ- ���m�0W�ӆ���k����kO~�:��.)-�?��v�[����=.W[�L¬:������Y7sr;t������	d#Pm�����h��0�-�rۅ+�J��N����C�
Ѿ�w�7�ꕗ9����&�k�F����>������������F�ФH��X=
s@h",v�����\�Kx�Na�,��.��_E�ELS�>t<Z��6Ő���kf�,&�x
�� ��Q��`~��c�|�;OK	y������J��}�s����U	�"SIp!�0�1�Ԋ&�>n�����3N�}���UL���%�r*�yG�9?��Y3�����"-�"�%lA	�H=�G��Ԏ� cv�q8��g�E����<<p?5��w11�m���4kӝsˉ X b��[��n�=���.�j�{L/a]�F��m��hݳ�e,�X��8�U�@sp�4��$tR/�����B��&��e(���^���Yه��.�TElhqzG� ��F�6�H�eL�������,l?[�C~�gf�v��Q�r�%ϛhe/+�z���ˁT�P��zw� �Xc��M����T�����=��SP�Q��t���p���ʈ�L�BSFH����Q�43b�pQn�_��]�ǜ��D��9��L��h��£1@i���G&�.�'ӽ>I�Ϛ�S��k���qL�2�|�8��Ջcˠ�
���L�$����i����R/���`�v�:�����r,�RAWS:m�DMv#�|���0����d�V�+��;4��%z�v6�K�R�Y���)]z�Ր�{4G��*Դb�_�L�cN�d��i���"HdV��/�@�R}�7�Z�/�u�.���/#��Y�V@�d��K�s�E���V���n<���ӛ*P��߉,�ƶm��#&�_#7��hvEzQ����`W$��;dx5��6�X��U��m�Sڭ?�Y��j��j⋔U����D����u��N+�m�eT9��Q	�+��Kw��3n���e����UW���_�m��_>�4*qT����I�*�9c��{E�ܠ��>%%C��Y
�c5�$�#め!�eLC��p
7
I)҂ƍ��ɠ���df	9�����R~' ������l�q�Z=�+"�$�3Fk���n���Sr���&��\�t�o	�����/�\U�c���-7��-⫑�G�¿��Az84�E/�d�)�#���~Uk�rǃ������`BO���ڿqO�cb��X\�5�V*ab�G#�'n�h�b����g&J�a�N!���`���՗��6��ѕ&�?O-4@�oW��a���,�S`U��8n-o ʺ9�3ÏB�)X�~�AҨ�a�*��_���j�2s��0?�<^����[����qw)�K�
�]S��T��o�k���X.r����¢w>�T8º����oGcW��)k �]�h��ь�#S�\�g@&���\�*� E:o������3��ks��g��G- �M؂����^�|�=E#�ki'�U�kJ���턻!}/ӱ$)�=��.@�Y�,�pt�i�į����j�'��c��%R����UT[�T��Ԋ�=�:CX>�i�UO8�u�]�l�>CԵ$���^85��{LO��jN�Uȟ��@���/0x^��ֹ}���1�c�%�S�@��?��ک� 
4��e�xM�	J�_Tx������8��{�L��_��R��P��3�賜�P�E�	E�XC�l���Bq[�|�Y�d5��+�;��t�<��np���9�]���M�E�(��B�[�0H�����s�
đ�#�i�$% \T�O�;��EJ�� �_��4�~�;^�ɵ�c�ȄS�R��*9!��Ll.�>�u����)��.PXЈ[.ϧ�#	��S��I��_.\�j��mM2������9�����ޥ)U�	g	K^4��l�Kt�|wc��t<�L�r0�8�'m��	�s�=&$�
%����&�Z��փGߘ.�9��`�{��1^/d5��1x%�����8&�-.��rN9��Q=`��%���eb'knN�������Ѫ�5-?��U�W~C�4	����c�ʻr�������V��O�0?�x�>����m3D�pwA���)��:0�)(@����/�֫�DԯX�3����@q<l�<ą�'����r��(ۯ�f`�_&�D8-�Dwb������y��E0�ݎԯ��I��cmh��
r�w���;�\����{���0#Ln*�`f�N\��v�C{���0��m�:?[�=���N�Jx��&oY�@�`� ���s�wg��G��XApeZ���G��jv;�^T�hewr�vn�]�Yj=�,�M���Q��:�;_W^��!)d{n�����d�C����� �pS�cN�>c� ��6^���h�Y`�Ni�P��K-�AK�p��)wif��^n-�F��+<�}�C
� � ��gV�z	�Ⱥ�O��7���!T{�]��_�%|�kS��9)��ʮa��ex$#�j4>������TX^�j��/��1a|�VH~�.ψ�+%Ò��U�S����r�P�)ݱ+�a�5���g�t�`u��Ӵ-��tv�w�HW}�V��h0�£���s}B�N=��8��:�s>�n�o<�"�+;��zaa�����|U�Bq>�f�޿��C���$�Bw$�l��ߢ����c����donzX��̆K.SH���*�4[Qm,v9��S>�ѹr��b0���`��,=������zxn� ����ri �ռ�)��S��� &S��ɁU���i��b~H�>���?l�c��A��c�Y,Ot�BY�T&�ѩ��JEz#/{$l���-3g3s8�^��u.H�۞�,&�N�a��[o�{*�0���$	կ=s5���	�]�[�Ƙ����J�h�T*J��#��7����O�X�{���p�d'&��XW�Ll j���-bʞ�5�e�_�0�Bz�DQK|���8��C�pJu��W��������c\��s�d>��ۿ����WUU"s<�^���U�i�Y�R�+;�x�
� �>�⒰i[X����v󧑻V���63 Wb׉�Y�<*x���`�U�'c
M�v%����GV�޾���&Q�).�u���ƛW} �ݫ�\��w��/��<D��Js�R(h7�tAT���)�p�1�>mV�y�T�YA׌�L���1c�XQޗ{��ap�o)�L}o�UV�����HJ}&�;�F��:��%�w�@KP{pk�ʚ�Rޯ}��?�B��1��ѹ�u諿<����)RY-%���eh�pՓ�ȯ*mS�t�U'�k���V�`5"o%�r�r�T��UI�����6%��a��L��5�l���`�T徱��x��)@�&�_�����D�Q�G��7Wm��=�W������]���NI�/ ��d�y>ھ�",Q���_DV����ա��;�s�;��W's<[c�4Kl븺-�B�0�j��A��A�Em�Nij�-������ "��Jr��O����J��:bw��^���+d}o0P匝�5��dd��S���pm[<��tﾧN�i�iqUr��.�e�,R�A��ٛi��K/����,��S���[ Go��I%������C\�I�u��fA3�����1���8~	:s���s����$q���w�T�uiv�/P.>6�����3l������ㇰ����(���iO�&y���)����-�F��C��ΐ�Kr����Nv���{m��V���3A�SD�[�5Cz �_����u�<xO�߈�$� k��dAb�{.��_^F�ZE�	�G?��r5����,W��#�6��V�᭨[��3��2ϿX��\~ M��F�����iF��h���_�ӓ��Q��gg �Q]o����"߯��no��eW��u���yj�T�y�BZ�]C� �1	�z�`8>�GH-!��T	�����? ���yʕ[�\a@�e��3���0�q�Y� t��T ��0�c`�R�YCPi�w��׸$��������_w�H�.��n �S��<6�:���3��]���D�[���z�;�1y��$=�^Z�����w\�I��䃀�ź%�_!�y�����I��PSL@�bK�q��3��m(�J�mrܿ�w��*�u	&�������}u��*�����Bp#\��8Ag�ma#��!�? �o89�"�3�Ï(�&B�/%QO���aX򛪂�˱`��k�
�Cc���3�Z^���	>ou�z?,K��_�w<!�Z[|'Δ!�|�p�N��ű�P�î�X��N6*hT>]�҈���t����{�s����h�����U���q]n欘'=���]�E� ���K�Ԙs�r��8Ս�����Z�S� ����v\ rIN�=&�g�El^l`����'�5��3yT��p&�|�&� G�Z�+U����a�d��B�y.�B~���W�޻��KC��l�ѡ�S����pk	z�N�;��w��zܕ �*�c�Q��7X�)Oġ�Zr�9��<�Z�f����^H]�(��������Pe����2���U��on�_�r���ⷬ�����E3�=�i�{�C�'T��1�O �W"�������GZ�)qQ�%<�v��Y�� �?�:.���4V��V�BVc	GJ��kR���Na�MaJF'�9��L0}ԭ�j��'�f0��R�G:.�hEP4sn7M��� �3ǒP���_X����k�F�����}��L��`�\�m�������8������ /,�����wAP1�������"%ÿ��)��������g���a�B��e+|��5���w�O�ܿ����� $�� Qd!�B�~��mޛ2�H��̩ ���[`�T�^�Gk~X�,�4�Y��k�
p�P<t�\ �㥽�� R�f;���ب	�\?d���&��ƫ"Xm5�ڝ��g�B�6����wIZ�?���8�-S���x���o�=�� ���J�E!�&
�z�\�,i2�������'M������� or۞��emqX$�[��h�o�M��
��s���	��k���0�./0��sb�(���U<��d~,|�|����,1��c�i{���f��� ��X|(��2�}�`r'����A�H���H��������,W�]�����U����{�z��ڥ��"Ĥ.]x��LK��1�Z�`�X>Zѥ��-�T�&����eD�0�����P��k(TP���>Cn�k����{{.`�-��61zk��.9�E���!D�yz#��ϊej�W����hY�r;s����CJ��h���B����в�Ч��.'H��ہ�{�����o-A�B+k$N������U�C1\'�`� [��Q�e~��B���������6�u�)�
.= ��G��@��V�Z�Yb��G���<�3E�Ez�7�.CK!��M�s��NG����l��4�O*5q�ԍ �C��.��+�u�+�5��/���Z�v}'��(�Ľ+�a��
��ˢ8�\��L�'[.�e3�)e��IډE%O��D��".L��A��Iv�ڐZA�	��m/��Jޙ��7>l� ~j~�1�e��o�/��?K�[.'�>���J��XVp	F�GG�4�x��"�=�*����Xh������)�zn�|�H�� Nkv������u.��΁��>VI;Õ�2�չ6?�y|��ި�<���M�U|� �_�:jK9;Ę��%��b^�����O�V�W?9i�ސ�]Y`���ׂ��A1~k���×hj9�`c���ļ��HG�����u��6�u�S�z.9���،6�17�G�bOV�<���o�(��������M���N��akI@���m���GőŶ䑊k�xz񣇽;�8�W=��*y�S��p��ʼ\5��K��J�BgoU�ΒM��_��plA<��/ ψ�f@?r
�WD!�d�c3�'�`�e���5v�@�$�{u�o��/aA
�#��h�;���=��o����:\�N���yA��ط+�|ݞ�|�> ���=�.`���\�U��O)��送��?��g$�?�Kߨ����h�N�f�J��"P��=�[���kb�$;i��Şw��z�Ѭ��k��j��񒝹Z������w�msH�h��1���bb��!�4�@w�B�v�g<u�X��$c��|H#%��-�3��E��F��Uus��B�Ȧ���Lm���������Zw�M��^��J3Y���9y��'�~<V��4
�V���r��uG'����m�z��� �WY�^A<[�kt�:���Eo{VC������=�Oּo�xciF�kBX���iP�-!%0�p
[/��+�`o����F�}ʆY���<��<�j�'>���C�?0%�{_������2�eyG��ɽ����@E���Q���gq��>��J^�(��hO�i1 �#�x�9�!,�H�[Ř�t� �����,��*��5h�H����� VY�Q���V*�+mv� �\V��{#�����wA�x�ʮ�����Q��쳉c����`�X��֛H�H�}��.���l�An/����fM늱W�����d-S�M��k;ϳ�Q�����ܰ *���z���6!(���~��kx�sJ� �ڶ��_��9٣T��0'7���!9�i�Sߣ}��!�+���y����᏾���|(TU�J]�C0�S2~K��6Y�t�p�nD�H�'���~�W��X�[�W�a�)0��w0��^XX���~���N�L1Ɋ��S'�'48�̓S�ؾ��;a��:pp)>��9}��D�{��xY_�\�������X�m��-���Q�EF}�=&���m��s8u�Q5�����������֞A����K�4X<tJ"E��6��-��=WQ�sy%�\����£`A*�{��"�L蹈�g���,j�pM��-]e� �i����@�t��ߌY���|+{��Ab��ĕ��r��-3�bMw���	Kv	���|�����KUHӖD
k��z�]ߕrHqc9E
-Q����IVg.��ƣ�Vw��DI�v���d�֔C�"��ۛf�� bo�!4��-^��by/V@}-�/j��sU\��8"W',g �6���̜j���!�	�2]-{)2��Y�)�Qx%w�RC,ل���p� !��i�a�d��.�03AL�G\�8iZ��	�[���f?Y�g�{]b*���鑐5�������	״���V�W?��ZK.I[C��h���{����3	d�-6�n=�;'�/ � �4�b�����0�C��%]�8�Z;?~����¿��)����(#��bc! �B�����gg6+�c��i��O��;Q�e8V����se�I�8˦�C(���{t?|R��7J��5A*�f1T&F�d��g})UN��Rf?����tً���uU�=n�Q鬊J��L��vDT`�w�.�G�|v�P��M������-yq ƅmw�g0�3�zk��j���Vț�{#��o!�-퓘1�(�U^��D�fe��ә�T�9��D�0��sF�L�F ���I��ۭR��FguR��(��r�Q�1��k1�c0:�����1
\65Ж��.c�Kw��@H�X�g��`-]��ߠЫ���c�&���s	LwB��L9f�w�e���\�k��^}�]uA�R|L�O]�!(��	-��TJŕQg8oJb��-����l��Op�� س��QH�u�h�7h���:1���g�U*�T+��dݸ< m*���qQ�ٮ��7h5�.c^�ڍ	Ǯe�����9���{�0�_I�n�T�
6+2�B2+�܎$���D�{{� �s%�?E
Ξ�f��aJ��m���lL�P-���ȸ�L�.P��D��9�A}Cԣm0<�X�rЅ��,��4����5O� �����A6{�6^�{<�-�!Z��U0���T���G�z�?�](2B��XQ���O�5L%�E�����Ь[=�?]�&�~Ȑ��Rq;���;w� ג���>�~��r����Lad*����cC�8��4P���
��26�
�//=֮�ݜ#M�h~9s�X(���PGoO6��B�M�3+�փ�D�p�4	.�E�ƌ�K�5*k��Ύ����I܈	(�Q���0�s��{�p��1���:0{�x�%o�ॲ�z`ΫoWFgI�g�-�B��_t�=���z�L��
�k��^V��W,�=%B�DN����|��X�vv�f�T)�P��1D�=���AJп}���g<��U��Av'���L�w��@�#�8�'�(	���Nr����F�`�	��X'� ��0�ۅ �����a@��l����\:�5��4�	#Is�|���z�k��d�T�腞�P�8m(#�12_ ��|���{��S�Hp��^�y̶�ѭK�l��UG�n��xս}"+�c/�>Z>_�Ͻ|CoV� �:��U��1a��y���W�}�o��A2�^���&F�����Rskg(���i���j I�d�����3w;UD�����^v����W�<s�f�CK��,�`�o�B��Hڃ��֪��u�r՘��E���-���~����=Bn��`l�D`@��ƫܷ������4��KQ;�֍a��� �5�<�z����S��nѠ�^�"}��`X�����-�<z��a�~�`Q��"Mr�<W�Z>m`&P�R`���-�k��L��%qIn"�
q[�����<������l�a�������~v}��v]�A���:�#?_Y��I�l3�-�0�f+����Ě����7�����^;%����@s��u	?v�e�ubtS.�Em�ZنꅛAܴ������Ay|�۱����Ql�3��F���u ��y���v�#�f<�!����X� S]$;�0�4?��~��el�r�X���e�L�WD�!�-wT�(�,@li�Ë��)ܲ-��`�GƗ�Y�$~0�wu�7ʛv����ȣ�d^眉�9F��s+���.NEs�ؐĕ1��"<k�#4X�Ao�Bq|9�%B���y�y�=u�x�Rq$����`��6���or�BJ�{�.���L���V$x'�������߹Y��B����J�4l���
'�����v����_�*~!1��O�i��}�>�w������|uEx;
�e)�[��´�@�Ae���Rѧ��="□HO����}����0�]����ʾ'5��RJ�#��Pް����W2ա~>Y�˹u��+\����*ٿ �<�v�>*T�n>�W���I�;��fFjw��X�q�s	�^Č�{^� �W&�=d���h|�"Lk�����v�_ti.�[zy<"�aŝt�90��E�'��%��!f:��Pb��P�%�}��͓SE��P��Tw��n�@�Қo� 82.�,�X�y�.r��ӂI{���?Y��D�3!{���x]�3ț&����aI�M���>����n�\�t���!�|�����^�O��u�������V�6��fb�k�}��Ʀ��)��#�	9��"0NZ���<l�[j���y�B���j]*�pp��hk;	�J�#�����z�_������B��q���$ �n��)�>�q�!?~�Ɵ����H�^�#��E��
�`�r�Y?����׵�#�Y�45
W��KҮ�;�' �h�.^`ow%FwuA�����IC�!M�n��wu���2�DҴq�?�2rhA��Ŏ++���*���KpoH�KL@�c�e\�~�Iݳ��ţ�~�C���2z���9f�\6�Ą�I�,��ء��a{�<B%�3��j�q�'oQ���ͨ�"f�P��HzsU��^���6�\�hb�%	���t��3j����gE7�5:�,�[���2�}��H�d�����WY{h�3�!�M�i�Q��[�+��/��+����)�a�s(����5C������$��_��.����Pn^c2��q}��${������w�t�O��9{Y���5kFg�!�gd̰f椀�������.a��6�k�Lv�I1��8���)�h�ނ�`�XL�p7e��)�_,����	�e��8��	��)���8ćVqA,{}>�0�]2=�jC1��(s>�*`�8�����
��U��Jو����~���-�]�e+ױ:Vy�A��	�)M�V��'�1�FĲ��'�����C�����?B�I�W�����m��G��e��� Ql<�.���Pd���*�0HǟP����$�<L:���~��фg1�F
,b �R���"��+�h���꿽R��9OU�v����7�H��#�eTo-�{+z�O�&rc)z�`&���!�8g��( 8"l��؅��-��B�����:@�4m�,���JPn��Feǥ8ea����B��C�|���%S�w�u)��p�4峲ra#�£�pU�+ F�����X>4�i/����p��]�+��M�]��M\�S�.w��n����0j~��)ެ8�-��M�&p�R���r��F��$�^�-�6���m�*�y�gC�G�OwO�P��v�!Mr*l`~I@��Z����Da�d���=��<M���H����y��*���K�lz��}��k`<5fc����$`��Y{�;1�%�-�|��-?�TjjU�TM����-/ᙗ��pQB�Q1]�@��!����rm�0z��=v;���y��~���p�(����*�{*:_�w���ǩZ�x�~���?�j>��ŷv�h}u�qf��� %vrvX��K�tK����4r�e/p8���j1�l�~�b��� _>X�����ˬȍM��a��R�k��RD�m�����n�Ő#!���a���Pl갱�n�:	n`H��~�ӧvC�?Jn�k��nz�����F@"�l�%�/R7��ԧ�u�_��'�m��$��?)D'x0���o���˝pN=f]p0�1�����Δv �˵i:��T)Y ����0��X:^aڿ&�c>�Li����n���ۢ��s�FD�{L`h���f3��ڥ��D<��@$���[�r?�i�'�Iʷ�-��X�R����PӞg�OY�.*q���1��D�C��?���:C!���BG �hR�v� ����p�sn{��P�0���(��`H�)�2n�l{� �%�K��/߷7��W�ד�߰^M��'
��U� h�9�W�o>@u�B��7�g��,���w�C�]m�A/�eű%0Չ��X�Jsb�S���bf�N��
�"��:��{�M�6 B�܍��Nu\�^�P�i�N��M*�+��E*x�H�)�u��l ���+�|��ϋ���W�ʇ��������7C֖��[�B��ad��Ql�C@ȈU'�v�� m��w�`vN\5�1��e�S"�c|�x*荰�;<_��f����PK�nD����ngR�@�/�9#o�T��|�/�t�G@�U�y/n��_u��5	�FU��*K���Y����VI
�j?��D��$VnZ KÃ� ��ꈒ�=h�/H����4J������о����>Ha6ۖ��v����O	�Z�ƀl�19bz��;�$�9u^�|Q�0"��F�˺Fta	�Dg�e)��/W����S|�/|b���I(Y	eW�o$'0�޸E��-�; D�Y�"=:tǼ�\�j'�!�a��'���*���h����p̿��W�QG��sT�b��Τ���&�u�7�ɕ��]�GpKN!�.�QGFy��V`^p�]�f�A�)og ����<֠��m�k���`�&$�Y7��NN>iۮ~2�"���H��RV'�]�0Mū�BퟥW�z���j���n�&<mq�ܱJ;+��W���'>c��Z�g� 嚁���b�HtZ��-hmy�W_	��h�����i,��Ę�d&��U�3��hm�L�խ��G�Q�?6�)�dL�l^i0�V����c軰�d+��l�$�_����f0*˄��lF�{��ℾ�T�p�h��{fy&�zf7`^=���:s��<\�/7�I�^�í��bK�sϺ�M����N~}��㸓�P���k^lòItL�]��]2��D���g6��ЁT�c�^ǽ�?GQ��a��2�xhe�Es�n�P[�����lb��e	mIN:ӧ�ɱ��#U�����Uo,�Fk��~�����)hᗑE[G�頇���A�/�nau�G��#�Wqc���s�����2W9.�^�B����p.^���Ψ��w��C.''�l�nn0A���}O{cFL<[�Q��{(�|�a��9�ԪrY}��	_�� M!d%�cM��jJ�-@�����yei�+�8���f�3xH�ZCy�xw^��!���\b�0T��2l0��
O��o�V�wz�����TN�1�ˌ�@ߊר��L�}��<�o2�z�4	��˰�a��;Z���kތ�láq����ga���޿6�61�E �ˊ)�d�O�[�����v2�F"�jE���k-�0$��"����|���X�_ ���鏷^��@�5��ҹ����NE�ǳqy��$ǅ"i�kGHT��:�@w�M�z�/��o��暸��$�f���D�J� $~p
|Fh�hV���ia�d���m�7{ĝ��f����*�0�N��<���Z���2�f!��ߋ�\�9��׏v-2��4A�jL}d���0MVA�7���8|0$�������%���%�@�l�������g��8��O�d�ˤ+W`ƹw�4�OAޙ�Ω|��ٷ��a�{Ux��(��-��Z����D�3�V��d�2��k���qJ*Ka���U�G�B����[s�6���֟xU��K-�nYE�)�8�Q�4���臌Z�R�T�h��oKj���H���2�1��
�y	�:z�`�` �<ڙ��HEG��(��K�y��#lbX6A�4[��B|���=��ԭ��I�:>n0`�<��vy��I����H��@�+�yRk�}��/��t��v�ⷲ�LGQ���ü U�N!D:�9A՗,;�Dc&��_� ��� |�������}�^��ɨ!Z0C0��Y>��v�1/|Y�^� Ձ���[E�z}�|����Q]t�:���d���RKk�{��QqB��uh�9߭�N��-I��]�h��*��	i��Q��\ů��ٚ�:��$��y��y0�ؗl�م+wb�*s��M���cl�Tv˹R�"��RE���y)��D���~����5c"�2��N�wl�0�Iu��6��$C1 Q�Us��~Z�\p>��[=�I-���呢)�5ie<~��
>Wb�n�K�0����ZP����XE�����

Q \rBh�����ܩβ���
�w��B꿭�R�wŞ�N�cE�:25��������N�����i�A��.f���3�S���%���y({��Ȣ�=k�&_�?������P�F��
G���Ɖ>M��̴�
僷�-��A֜-;3f�����@�K�G�ݫ�Y'��Qg�xPO�t�%+�����]pt�V:K�UGeT�h^���}L�I�]I��9\�� ְ\�4������Ĥ�rf!�YT���fC��3`#�tq���VCnt;@j绀_�ځ�Aj}�$.ڰ�����G�Tb�N ��La[e�}�V��M��*7��'~���Ѭ��ܸ���*�p�i�8��J@��}1��t��O���}ὓ��������J=mp$��빖��9�P�}=@ڐ���(h±O_��k�UJ��]2MGb3�_��fe�I�!>���ۃ�)�4\���W
Z�xg���XG�_Y+��(��QA�Gu��6Hp����2K���_�S
�����o�����dY)�h�$h��J�Hҧ�������ӁC/��'ܼ�YfkӼ�R����'lp�bC���z'�Gq�u�G�5�A�>q���ET�N��h K�
�#�ɅԬ���<eѭ����q�1e��nا�z�����<��A�L�z�W���3|u2�O�{f��YtW6+��b�MO�1*�H6z��PZ���h���S�����:*G�";�6¡X�.|]�ɎEXd�k��l��������y�!��f�=8hi�O���G5%��խ��9'����V�;���Ą!#g��\,�ͲK�o�Yy|��u8�}\d�Z0��lC	p���C���7��=��`�Gsg3d����0�9u�SM7�X��a^�Q��ϻ�(#�(A���I��	s�F_5Ք����?���#�X�GK�#��v�<v���Mx��a��|���l����>��G<@�א�q#���7��[����ʄY�,���Qj��JJ�m&��P
-��}�2�Tb	t�;��Qs'ov��{�D���P��N���v@���RX��fq��-�"�nFbwyˀ�����'��i�c�T�u�ވ�C��(��: �g��l����)��k�jEned���$�㻚��.v������Tl�$���'�L]� i����k`�CX$�0�j5l+A��wU�A�,�3
OIJ>Ӊ�3/x��Η1|��ʇ����=
-��K���A� $?�A+nU��~�t�+��l��}��A�3�2�p�,w���C�D���xN;R�����PW��K�<(��eqk��s�l=�#y
�=��'�9���3u�j�����Xs&޵h M�}�X�56�>��"��7�
�����C=��%�t��[Ǜ����H�z-�ov���@�.m��_X��u��5}�?@�`�̩�D���J(�m_t�� s�ub�?�5�17@zڄ5�})�0a������a�=-��]G��~D���4�Ke^��~B��p����w�.=鲼��/�h����E>Y�)�Q�lC��d6_�g��.F�3q��9�[��(o��� �l���"�ʙ����?��ȀT,ߌ�w���U��������rL���rS�q�4*&G�K�Eٰ*�QM��a�[���K�t�an�n���M������"�b���W��Ý]�E�n`�<�aBƶ��4(�l�'6V\_,�G7	Iv�݊��ͼE���Gd�b�@���dq�Q�P	��,9Nh�L<����I����"�E���3-a;*��1���?i�U�o	���\���{��Le	p��g�Ώ��]�~��@���gk��`Y� 4�:[�b\ۻ���n���M0u`����NN���n�8�j�F��gZ����L���n�mu+1�)˩���|@QwԹH��tT�&B;qrR��=3�Oʖlo���N��^�)p�z�(v�����k�Ev������am���eq��Y�3 2"!G���l@`'0c
�T� 탯oq��L�����^*�}�ztQ|�}t�ڙ��`������`(jX�@5v!�ds:y�n�~Ξ���=Y�C/2�4��Կ*�৿E�æU���#]�Ķ��,�ŷ��TA�ͻŘ(����uUY�yź��-Q�'&a��ٙ�7ѹs�G�O��WE"%��\�G�3Sp�ٖ9J���<���Z�'���K��oː�b^���Nh8�Ԃ���h�����-f��:�R��A^q��������R[a���+)�:�~�,�����t�H��gt�FV*�x�q�ε~;��ᕚlke�@�bs4R�\ǁbe9�
8�|(�oD�6K�S£�O0P/�ݩ�H$	��������a�o����y*q>���?�!"�e���W/##�n�w&"���r��$+l?�~<u,���QD�Q��Ҳ�8V��B5���B�b� tff��v�<.��;@�$�,k*�ύ��~��Hٱ�Ws��م\��%�F=!�Ɓ�s�"�6#��K��Q�@���'5Q�F2��Ѡ/�A�1��,d̴g�ރ��)����|X5[S����]�>e�Y�U|F�UV��x�7�r��-s�:�ٜe3��D�e<�Hr亳U�k�̘Nx�p�Z�h�9Y5�W��YxG�̨�+(����5�[��t��lk�6��ߺ�A_��定���Q!��7� �y�-1�@
fv%/���Px]_���m�O��0�.�G�DZw_\�1���5�Vy(!ς��i+
�/\��;�@��fo�c�(qmF]}g-h��$��YV+Fa��{��G5�c��Qh���D����)=�������5`�z�)@��C����������Q�����ȹ�Z��77JE���/N�����Ց0�>�A�Ӣ�77=v�?��������i �^�['�6!Nclvt���?�i���x�3���D-��Kx�Y������euA�����?���}p��M�N#<�
�B̩���Jj�P�c�M�]�3���{��hGƙЮ5}+��:���蟆=ؖt��C�^m�C�pR�ֹJ�4-��!�V��&�lS�!�\��A�bY3�7���_���Oa3b]�C�z����ʝ	,�F��Wd(D��s^��v�b.9K�A�;5?�j^��Ջ��M�c�#@X�16{���)�{(j���K�.v- ��k	��z{�������w�}��Y��k���m-G�Di��W��W�d��A���!����e�>�1|>uB� ���dZ+�\kR7(*J�cq}����YnY��T����Ī#�vQ�Y���p8��Q�̓7� e�d�~ʸN��Q���6��,%ESk!��cO+ �E"�bR��;�&0�T�;S�F|�5�2`��ZO�Y`��k�u��� ��� ktg$�o����8u6��T�?���ˉD��/�Wѿӗ�Vw������A��63� =t�F��3#a���^r���Ƌ��a�*�w��*0&���{�E���6):R{n�Ѧ�F͉&�d�(.������еw�:��X|��b��������%C�P��=-�������M/�n<ve��;Ļ4x�'�l" k�M��ԁb���
��y>=��G��une�o��͡�fΡ<�A_C�	�S`��%r����El�ݣ�`����@9���SW�n!���ա�+�6gv��@(A�8��. �H�h������Q��b�W�du�Ϲ���^1�\~�{9���n�r����@�b��[`#�to&��Z:ucԒP'�"(I�c��K:2E�u��FK�8��ȇ9��?��Gll9`�_ �@|� #孧`�̝���fn�U�#<>	�i���dK�ݕ..撩�~�=��~L`_�o�H"��ҭ�F�%����0*-�x���F =��աn�k��(\SO���Q��,$�	����a<���I�Ƨqa��z��_O�+X���L��ѼH��+�j����;i���o}����-6P4�n�R�L@V �Y2z�x���-�͉�'E;�W�Rj�<X&B��k��2acl�C&R_�%��c�jv��K��Zb��3�[�h{�HoH��G�#���P��}��6t�YY�ٞ�c�z���Ӿ�V8l|,����銿ے�⯍ �?z�W��?�/�;H!�Śv���#� Z:���x�/�tZ��ٚ��ڤ6�s��z�U�1r��i�m��zPE����s�n��ք�[7�W�V�@�n��{ސ~'9M��U·辳O��$E\a�*�>���R��U�e��ݷ}�ft���y:JD�&��U����nӹs�r�kH����pf�R\���)�K�ef�k��֨B@$-�K�O�P��QD�rґ���x�:���W#���ſ��t���Ĭ��Cɿ���OJ�E�����i�+������JоE�9`c�d\G\i�_ON�\�s�ru71\�-UE�>9Э�Ɵ�=K�v�!�d1h�̼FLZ4;:R�ҰA%��Ƞ:����h|I)`�l�oQ�{5�~(㓯kq�5J�/AX^���H<Ӧu:��d��U�|裎��$��(��=,��rlg��w��e��\ǵ�k��r�;F�u��t�m�{��$t���&a��p�I��|�%� L<Gޑjp�G�[8��?;??�x�e�W��p���v�n�n:J0��7�H�7ߦt����d�DT���2g�ɩI�U�|�F!a�g(%�Q4U��,��\6󓃭��hyf�6ı� :E	;Ɓ�����M�6��MC� ��m����S���1ut��[)G����O��7��^�H4�G"���F�����ȴs��2ͣ�z���T+���I����y�5J��<���.S7��2Ik)��Г����Mm�ģ����m�Ӱ��}����Ĥ�`&��Z	w��ɶܹ��I��:���}�|����R��u��u{[↬���k��\�R{����M�(?rU� yj����ݔ��J_�~U����HS�b%����dn�av��#B����������.��L�Ɩ�p��Q����\,O���B�b�b�՜�q���{��+"3���՞{�F��y�k��u��1�u?�B�� h�K1ǍI��>k�`�^���?!�gM{O�4a�(&���1Bj��%M?�'�ꛩ�C�Qi��}$�ʂ���-��#�9��Ӱ��%~�\+.��{�B@�lM���Hx�����Y���G�}�9�!v��������RJV�b���U��O�Ɠ��H�lWK��U�M��m��A���`d�8ɥ6o�l�Ƣq���G�j�J��1�m�/ɱH�l����n�9��NQ��cr�숈�$��f��R9n�*S���}��n��̹�{sdw�P/��f����}"���T�d��WP��tv���_���>�('�aYLc$�pHV�2VY�S�B�1�������2*b�D�X�ő��PL����Ħ�|�	�V�dC	�x����Xb0������{��g{��Gj�Y�������)o*��l�!�^��5��,���dH-E�\��J;I�,��]宧�(J���P��0����Fy�֛U����(�)l](?�bGی�\�>�s�J�������.�`�h^�x�:�E�Z��s�z��N�m[ ���N'���Ĝ���B_�+�)��5�$�O�j�5z���^Dt������0$:s��7<��I�,P�Sh��zaW;v�����:fW묇��m�h��\þ@A�rU�ɗВ�y��}���~L�:r���C4��N��lOr��{�c��G7y�\6�[����韼���Uν�¡��!���8���J���đ���dw�`@zW������a
�?�tW.X��2�jM�L1a+��L�ڝ�S�u?�S�E��d�Y���!h.��[���).�"p�=�j���%֘��G&�d<���~�ڈ)!X&�1}��V�|�iJ�/�wMV����Md�3�E�Ù����h�5 FV}U����#�&��6D�;�1����o0�Y�	�����b���7���1,�!K^�ʈ�]�&��Ɗ���O���;I=on����8VW!�h�5�8�'�g���5��l�~ 0֛��A�s-���}�r�EӣR\?�,B��k�I
��`��M���NHO�����? e�}��_s�������))�U%�zV���X�B�$漳3?�tC��B�fc�.�t<��t���
������R�x��N�g%�q\J�{Db�1�k�&��p��]!����`mM�=a���7�W�߿ǹh��(܌�TaZ��9�6R(�ف���.r��+�~w�WՊ��5�-�w�#��e���j##�Ӆz�W��)O��nCC0�+�|��J��rه�,x$j&�'�W װ`J~s9�x~����n��}O�Q��%ߏQ�%awe�U��Y�V�[��C� �~������$����t�{<��އ�B5�hB��ҢBU�Kۀ���j��Ri�W�w������ ���f{����,)�x����YOku�h�t��~���
;3���?	#
�;�����z��|���6�P�^=�QQ{�h R$���d7��S�<VV�17���?��I%q��$̓�xp��Tf͡�.tce?�U�o(|�ml�>Y������8��H컢�a0CU ��A|U�I ��cM��ݸk|fLшJȈ��e��i�w=���#V?*3���3�8����i��K�Ps`."מ��Fx%>�"��Ni~褬�t�R9,��2�w���d�n�9�)o�7�$`��>�\�0y��?ӬC���V��%0UN��o
�;�b`ߜ���عg�%Y����i��Ď���v�]�Ni�vn�lۂ�����}�Nc�cjd��u��Qh`O���W�ф���n��<f�����E�a�7A�l��rM�l-�Y<}��9Yq�A�b��(@�@�n��T0y��Q[�sB�BKqۅ+3�&��~F��-)��YYk�{��IB^�t��T�aA��R�L��<��]{ P���{���v��U����K�*�I�L݊�"_�a2�H��BU�^�&�(���������f
���oS��wF������/�w�������5!%��	�:<˅��}�0������x�&U���s�&��vfn@ȷ͚�<Jw"�Y��!���h��/����xX�F-�Z�8�����׉���d���OM�> ��u�}���a���ֶz�j��!�t<2{^���XhOg9M���t����	U8��Nڌo+��c�7O�QTЏG+�KuZ��Xuj�\�b\�v�Q�&�ѭ�v�f>M��[�\D8���'�e4%t>��C�p��ui���i^�_&i!)2��$���s��U�[I��@�[f��;�[��⿆.U����;U�k�l?�Xr?
P��DCV�lG��ǭsan��ܿQ���!���s��6YT�nzT���_M�4���Z�����ƍ��W9��ߋř9�r'S�)���w~?_V�t=9yP�9��E������K����G�&����8��l#D��no����ybS����	Y��:�N�瑵��"�XN���!���� �WzQ%������_�� �FܜA�E�%��ʔ)\t�G���� ��m3�Re�E�	� %V�T�tA��2{8_Sk~�j��<אP��h���'�6���g��4:n3p���z�gPo"���0�Q���m��kn�B���I�}5��3�Q�j-Lݍ�����D7�9᳕��������=j`�3-�X'̝6����.�tҫK�f�!60�����<�m�D�#���ֻ�ǌ-H;���OEIY�@�SW����re�����}|�� ��|�?����˂U��Ǿ�c��S�8��~����4��?����K�^|�U�L�������2�����í�z,\?��C�S�ө�l���/�%�r:�LpY���O��q�*rDX�na�@e���Lk�O����2y��V�,������^�9����?
c�������%�2�mx|��Es���F�z�_�+��Mm�@X������0��L���-��Փ&��s޿':zecl*�А=V��`�)	�,���J��x�����0�?��m�?�� �4�(��W�����0+��@�a��a>�]R}.vm�}'H�,x��2�햢�o�ASĬq�yz��ׁ��� �$p6���`�(y��t��[@�$�=y4��!�| ��"M蚹ʸ���ˬ������S�.-g��H�X/�9�ϕZS��D<^L�?��_3=��5�E�(�ga�FI���7��\�\���W�e���k������k��4)5b��ӝ�a�əb��U��R�jD0u����4AP��[˺8��-M���T�a���틟�D�(�z9fsL�uv�ɟo#���6#:��bl�^��m��#z=k��#����q��q�X���m���t�rPӸ��H�|
/���v2���EB ,#r�;oL�d��V��W��ϲMR�����!..b- ���?P而T/�ģa��)vr�,�k����#�׊?QDȑ�,�� ؘ�yXM����c�� �����WÐ"�,�uI耴�\��|(��μ�˺�`�+���v��Q�СH��r�i��&(�J<���֌���Q,:��� 
�8@�k��P6�ful�=�_��W8�U!ޯk���M7zh��)���7,��5A�t
�`�Xθ��d�c5R�C ���6�1��9�&�
ʡ¤}�eS��]ȵ�܁�L�����ֱ�-6jO��v�e�|F�(��C[��������,-��,��3Uv⬴��)�1�:�<@gu{'xs$���cD��Fp�����Ooi�Ǌ;�OX�f�Ơ���'y*�/�[B�������ÉƖ��p��-��zv�O��7}i��i��[X�ʄ}�#�$�98lMw>�XUn�Γ����&vm��7����QĄ�}���;�~��b]m~+�N�\)����/�PI�#B�/�->^����ɷb�Xr����E�d�U4�
=��@���zc�YN����_$�B�^�ʒ�J���_%n,�� �� ���ы�W�#N����^>��9�c$~(�&"4$�����^9��77� �8���J�V�������Ep�l�<@��;��$׋~�
�5K6.4@��<�yX�V[��[ІVnqdbE��?(��y�Ni�E�����t� �2��48�����v�u�MpXM��*����#o�%'�v���/�~w�]i�D���m��ʀ����ш�$�U]�B��Y���]��yB,�Sk� d��Ťa�LFKM7Oe�\�Q%�����	A4�&u#S��5�� ��H���*ťn�B��'c�mdӇ%Ƥ��Ĩ���6/U��\�_��K�'��I�ߖ�z`[��)fJ�&.�b��*�j*��ڛ��6���Ǿ�4��$$��蓰*K��|v4����1C��
�WKQ7
�[�{�鶨�0�r�R��;&���H�@-y�˧�_�Y7WW��"s�@�� ��}O�dL<�ֿ�9n��VD�2>�G��r)ƒ���o]��զaB����e��^������a9�B��6��O�~P�<(������D�̨�-t)�>r�w͇�z2f�j���3����?׊��լHLU#�}���ŐG���CҚ��Sx]+-n��!X`m^d<�Іky���v�+x:�6m��ٶ� ���Y�W�'��g6�X�!����(�o烳��GU�BJ-ӗ2�E�\����6��dS��AK`�f��D���F�������g�L@��D�ؿ.ݼCm����w_g��ؓT�P��b��v��IAy-2s�Ӂ
�y>���,+�"%k�?��#�[�����������s�w�o�pܖR	!�"Ր$|���J[��8��6��z� �
�� �Y_���'qC$cW�0�2��`�Tl��
#O� 3�|[�D��#o#Uj*u�2&�ީ3h�#�.~5��~M�)���9�z�x�Ӷ��Քˆ���.G��pD+֒�A�x��ɂ�`��G¸��H��#�*���#�������C62\�
��Ｍ�S t�\vVBep�O&�nI ʙ���**)#`�#�����s�t���f��J�r�=$ׅ
eA����PkM�6����������]%��J-�O?��8�VQhp�^��"���C����W/�|5wk���-���������Gj�b,|8��R�I���n����*ިr2�
�.��%�Y$�� 7���&1��I=�LK�\�^X�I��ePqO�4y��e �&�B�A���iV�"��8rW��
[*ڔ���B��n`�l�Ng"�Ƚ<����{�����oG�VJfE�[�6�|�R��}31O�ԧK��>9�h>���̞a�x�N�読����=�Ԋ�����`��-����y�d�B�6��v��ELMFDY;w��O�Q=�5�����[e�()�
"��ā/��(0�tݭ��5��*s����������	���rH�
f�S;�r���}?��+ꩭJ֚��봉����'~zJV~x��~Z�2�jAJ�т�.v���/q��D?�ֹ��>��
P�p!���,����6��04B����͵-���C�ם�Qؔ8���K�����H4���Ծ�\eF��ߑ.�%�Lvu�`�� ʜ��?eo�T���0����q�\�/X�Kr��˄��^�q4�R`)��ވ��{����u�4/o[�a�6pRa$����l�I�G׾V��� �e�-�%��ݘ_󚨌[�ag~,��>Z�|S��h����iM<���3>T�3o���G�W%Ɯӈ������0`d_n�i�B��Z��%$���]�w��#�?_v�b��(�l�O2mO�涅� �Xs�7�|c�����˴f"~L�8���4V�19��b��|�� ��YW��`%�W�i�x� r�|���0�3�	��Ϻ��{��r��*���,���9n�G�3�+�����t;U�&��3�>��m�b�ĳ�:��X��C�3o��O�Ҫ59 B�5S���.��߮z_�b��r4�2��Z,q@��n��b�L���� �PX5�V�.�g��h�d	�i����%������qH#	A�cI�i�/�틏F��)�\�^�7���#�	[��g�
~���Ńk�PY�Nco\b4��Tj��=ʮ9팎���,�r�M�1⡨ԕ��D��5�M��ۋ�lSU�y���$C9	���sEijh�Gc���&���m��ţ+�P���bJ-#]D@#�%T�����s�; �j|��Y5��K4�p�1���*����J]"I�qVJ�0�B��s�Z2��.yy��Hn�P�ph/���;cA �L=�t.�}Ě��n���TH��k~!v/��dT��B�iG�οKdm�xk���.	�#tv�Y~��7%��(ji��E��S0M T>ڋ�Ƨ�������!���k?>z崴�.��Ow��.�3o&��u�jޒ��b���.�[�m3�X뙲2�M'�*���k���1�����I�����VC�h@�_��G�����H�G����>\��N��:5ndHa����P�y>����}�_�u�D���;P��e��ᔟ���66���[1x$���S����Ĭ<�
]/;���p|r��	�{�??�6&?\���tMn#D�]�|`Ϙ�l���7��(��ISdj���Q��E&�(�P�҅�gᦏ�E�f����0z=��zV+���L�uМ;�����SО���%o�A@>����7��h䭰�;6�뭨�"���;�`������]�&k5��+�x��}�ʰq��-���X9�Y:�����Z2j���jO�~��j�Vބ�o�p�8�\|Ex)��bL	���Ml��P��T���8:��'�ť�V�8��ENa�����+�~�İ�X�c��K�EJ�;�	H��&���q�h��h�t�+Ma��o���*T翎�¬��-�=)�v�4�>���(<��=8��47c�H��1A,�֯g̾R��EU{�s��]m9Gؖ�R{�l�T���mt��z@��'t��{��X���Y��9r�
͝��-����fs�Yql'�
���I�Ĥ��L�
���F {���� ?!�rkU_���H)�LL�8xq�YC�����(�����¦�J �#�Y
ٗ�L���͜+�mTg;m�G*�͓�ǂ]��*س���t�[||b>nJ��W��
l�
hwC��{���@�s�������[����!�cX�f�?�r	�����ˊ��rN֦���ه)ڃ�m���̜p{�?��|o�2���5�哌��{a�r�?��}���pae�CU�����Q]��3G�!�y�9���Sű�	�:t��FA��޶��%�9ɧ��
�)���#=�d�C����14���VpLĨ�e�x�{>�W�<�P��>�J�Qlj��#��0o ���'7�?�f>N�X���#\C�}�t��݇�)X=��e��A3+��Hz�?����D�d3�o��H��,f����Ox�ߢ���miX(L�F&/!|�������"�� *�lIU�h"��}�N���1��DQ�y��Dj�t������EF#���Q�Q�q��˔l�C
��"&�%��.5�yX����>J�6����Jag[W�ds�q*�Q�{��Y�s���P��V�n��n�{�`ς����)���<?{� �{��V��D�x�/�U��i.�7d_	p*r7� ]���N�<�T�7�;Â㪂�࠺'ȃ̽I
ו�L,�*��6����e>��|J�'��$D��;��KEȾX>����~_��ŷ[F{c����^mX��/�������<�v�9�$\��7� KՕ���mu��[�U�v]l�WŘ=�j�ӏP7LV�O���4Ҙ�.��p��}����}+�=�|�]��IB���a��}dJ�u�^`�&Ӿk��.��I�D;�_���������*a� O�2}�Woリ%���,փ�"��;	����Y�Ul��n���5Wr8��ʴC�|5�8{޾��Y�%9�����հ8�칥��>kMVFH &@�R�z�^T�u�iD�X4_g�گe��v8������ؚ =�K���^e:���K$�|�]3[��<�A�zL��
�٫^9�M���epr�9^�n *����a{?��3�����3�jX��*1<ŻCvatʯ�X�?E�1����[���_U=q��5e�lj��圕�E��(U�u0��LL ���jPB.�ʁml��W��c��}8�8Ɛ�QX��U4�Ј�T� .m��k���ØEd�@/z�[my��M߾&�,���t�jݣ�Z��D�Ai��� 3B���G��L� O��nځ��=y��\����S���n����Ch�/�U���v��ȶ����w�����m��|W^��> �3E��2�h=X�U�;�\86(ݦ=$I�cu��+�y��Ln�(yt��&�m댕�f�wH���0�����UF؞�j�Ln@89D0p��f8(�}<�����s�æD��V�Y��I훦�K������4��7��ĵX��,�Mu2�����f��+B����1V�4j��9�zv����r6�4�W�SN�n��>$~���a�v�g#��,8�H� /�Ά0{�-�	��\�����ߪ݆C����l7���rɊG<�ػ�z-��������~g���(s��W�;��I��J%���4�+�� |Z��L8,t|��E�z�G ��|J�z�l,=(*�Ѭ��!��`1^a TMa��b����\��_'�%�-��8D��Ć�,�Ma�P�����I�G@���p�p�l۸�f�B�}��kn^��nP�-Jxl燊Y$� 0������n�E��ǹ��A��O֒��jz��3a�u���q�Bj��
�s��D3[D��-��YE�������2hk�]�bi�5�\a�䍦6�H�Go��v�����xYo�O��[)�O9uD��;�\�x�����P�\ɢ������"�D)��LI���z����El�ؼ�����8���L�8!c	bo�!��a�D��
��4�M�3�V,�	cX{/�~�;�yn��U�^ �Y�U��pA��K�4�ƅ�]!6�k_�v�ݿK��C��$�$��}~��,3Y�f�r��`tO:�}��e�*ŗ�{�n 1�� �YӉ��c�0����_�B�ѼD��8��j�����A��|
������li헑�JZGG����,=J��8�p(A9��С��J��n�6�Er��æ2Q�����P$�̒� ��12��<3m�,������$�Pʉnng�g���]]��wĵ����f�tCYH�Y6����ĥi<w;'�𲛶�y'�:�5O�"Evc�9�.󰫗��,mc�A��[�@�Z�`�(s||�����T%�Iw�3=�$��O��~�d���H�}N�"}sISSȕ� �����mF�x#��ig>
]:���A<V�Ofɓ`��E�B���1qV�b�V���3L�x�J�CƟu�� *�dY�1�_C�0����)�c̭;]�`�+�j���#t��)�儺~!�8W��[qmG��n����௙�!�\�W V1-j�rm�9�T�"c�1�!E��z~<d*��\f,��*f�>
$2���B�
3	:vv[����ztG$#W�J�!avt!��]�bDmX?�}�����R�/=�̑�Z�PPk"v_��9�]P�Ԛ���ԹՄ���W^�6�r0r���ۦ�6�$��ZC8��u����K�>zߦ� ;*,s""�7�h��yS��2R��~&�S�#� ��_���#�b�6Z���U�9G⻉\O�$�c�	�o@�=��A�� �kD: F��%p�/{FB� �)�S,��0c�V�%�'/M�g��Nbߑ C������>R�*& �Y*W�̵0&�#�N��K�=�Ͻ�3�/�l��ت���a�E;��yD(����>��R�)v�V���;¦M�"�^�>�
���j':�u8=X�Q3�GK��Џ��R�"�G�g$T��+�n�����j[���~�r�>��FՊ�W�!y���[����M>	�^��Ur{h-@�`?I6���P��]�Uy@-�b	��E�P��Tm�H:�@�p��<ZW=J��(HN",��g�w@�h@��b�"��ӱ�HߩW����y q�/�����y�*��R�Zh13�����#	 ׿mC�n��Op��VOW1��]F���
��6�86��7����[~�g�L���ꔓ�l�FB��'8�9��*aQ�'"�ZgE�t����0vk�l��Gq��<f!��T���j��ɒ���H#�s���8!���*lO:Ș���e��6n�S��`:ܰ�:%�ԋ��"1�����p)h������lS2:����2����f�|�&�v�J�f�,c�j4,�7��Ogk�=�K��ӊ� ��!���gB��H��@O��#~ S�o����vE��PL��M��~H�P��M�"�m����g�e�3J�1���و�M&ѭ;����3Ҡ[��Z���\� ��g��o	��c����єa�JL�޼ҭ������Jc�b�Hb�p9!������r�&�m�1B6��~M�yk���w}�\��������<j��E=��2��,�!���S#�&a�g8�H���r����a<� I�|�>YԌ��v�~�Ѹ���/��n&���]4-�r�3��V�ECoT��zY���d��Z�z�Wb�s;��7��C;B��	�{�2�b�up�ppd��G:���`�We�/���1�Ԃ��ښ�R}J1$�etaCۖ�I��t270É��=>'(�\�=_ÿ�>l6A7���d���`���0nw�y�B���Bm�!j ��*��=�2A/��Lî"�w��F� D�*	��: ܣI2��3]m�@ك3T�gQ�����{4��~,ZrH��U]����i�*`���V�ׄ�/��c�;�)�8h�Bގ�� 0��E�a/������ocPP�8�3mS$������	=�Ax�Ggu&;�Ƿ�����Qus4�����2T�)A�5t�������8Jg�k";�*TD=�!ܦko���<M;H�`� b��]�k����EQ�*�����pa �[@��E��"�]�2��w��YM�B7"w�H���p��݌�$w-b	�Xg�್�Xjw<#V���kc�}�\�]��1`��n�j^N��|?E.h�\�JQ<t�� �dј�^���&Mp�f���[heӆ����$K�/�Ծ3�������r��z���ۨ��y(����qFE��'}9����Dg/���D9 ����L0)�D������kvNd�t�x��_V(6Mc}wտB��8g��R�XR��&�h�v5A�Y?����t�ˉ���>��}�-奥�'�՘��Z�]�}���fx?~/�/�5޷�̷B�8�?�@ҟW���]]�pc��K�� �� ײ��<��o�b���a态��J���L�[2��l��Sض�W7�U�/F���Qv���嚇<��ׇ�o�<j"�Npe���Xy�p}բ�j�n���E��z
��!J���[��.���"����� ݊��w��y0��ݑ���>�a&�D5�ߗ'�h�����n'��[9TA��^v݇����}���$��ϩFf��Q�y�lȋ��T��"�uņ���3L%L�rt��*Ҥ�����|��ɭ[Q�
7�Uu�cb'M���U��8��Q9r�Ul�#�<o��a�1��7�EN�D#{O�Ct=%Ǡ��ж�a�GYȭ͊��}s{�*k]|�0e.�8T��m/�JG׳�	u�ѹ0�е��A��)<%��L*��%��-ݸu�d�;�s��I�����IWaX��aA@I�2te}*-����o�k�7� ��:��c0^a�]��b�z����VVG&��\��>���U��:C��6a:��W�ڙ��Y���V�|ǹ��1;�HC���
��Og�y4�'΀�f�V1	C4��E��R�)��p�@�Ƀ�Ԑ���`m�y�
=ћ@����h����#�u�к>��!����B��rJ8��L����:����,��RW �P���!k=S[b�d��XM̆H~��iM�^a�1V����jC++d���1'�#I�kH�3���M��J���kO4�
":]���Tg��:a�;^m�bs<,���	4��b><���j����'�B5�+-гCׯɞS�����q�~��D��Z&��:�_p�;9	��ҵ�²捎��C��q��C�U�������& >��짤��^뭺���U�pʊ�F+ ��7m�=��J\�Y��Q���1l�.zlt��`�ݦz�cx���B�tp�E�@��b�@ �����~ I�FT��M�E�v2�4"b�:e�$X��n�������M^����4/:�P��A�A��ePwo2����Ä<=�E&,��}���ȏ�>qi2�Iٰ������P�Iv3��dq��I-�F¢MS�8�4����S��s�a�����|t�&*�E�3�E^5]�����4
; ��Q��< ���w��	��Ps.��@C��^$G�-%�Xp2p9B��N�o����AS0����ϓ�b����]
W��=P6s3�*�)��c���x,�0+F˶&*	4����O�����(��O;aKQ���Ks�J��E����1\����̘��gx�|�)("�k4pluޢ=,TW|f����Uo�k�7�׽�5���9Nr�¦mlUU�t�3L���xV�&�����^&�!ȿ��%���D���S��\,/9+�Yee3�1e6.#����n��aɹog�_�=Ex�+	7�ۡ:d�-I{%��LxH`{������(�1�Z�
+���8�%榳.��ƨ˦��q�r�C,�j�v/6��|#���Ұ�����Íڡ�UK-����[Ƌ��zA�6Ù�GZ�N9.K��l��v���%Z'L+�ª �O�r�C!%���vr����ͥV��B��Y`��q�W�����<l�'�>>W��=@қmJ#���~�^��LJG]'�rF�l|�~u<W���-݊0���3��v߃�{�&i3�PO݉ܭ�d�Ɇ�����{Q�`���u�׸Ҳh�h�T�S��>��K��h�|1�ڨ��f
�o|����~�bsdN�(Z���;�ƈCe������}@ܰ4���׷����AU8��ϹK����3�b���7��\���I�ɁJ�,�V��A}�tָ +A�A'��"�������o��;H2/	,���R��^cRJtO�F��Q�Q���7<��U���y���u�����"dv�Xlh��t���1���@��'0�ᑦ�V�fy<h���;n�����W>����'�#�����[qY�ˣ�VhD�,��(X�t��q��w�'e��߯��V otLqR�oF{_b�_ؗ|Y�v"�z��xӇ�h]��	�M�@�X�y&��5��xU��lή��T������Of�~���,�$T~��a��k�,zs	���5��\��I
�^��B��薎�B�	�߬%2"�!f�����p���X������5,�O����U�jk鰪!���O #��yP��Cɠ�k
�NJ���e>�9��G1��D����tk�����":XH�\Ԡ��W�D���:<g�7-���x�Oc%��
%�xm:�P��{�Z�+�Ҡ�L>IGK����k���:d.z�"'M���y&O���R����pk	�i7�Vt�(H3���i-� 4=�s�2�.��T�-�#�x��,E��v~��T��$�+��ȍ3~(� ��Hl�����1��=���[�&LJ�V��7+%2u�VC���I�v��I��tT�+�.�j�T�Ŋ{�+�̏��sr����T���C�TL�]d���4�ˑ�1K�5�L�kmL^#�i%f$��w�-����M�ѤR�<A�'2��l�u�@�A3K�7sa�%x�Y�jU�4�D~��5"��^*�o��G,�W��vs��R�r�F6��;���`�uMx�\δ���|�x���:��7ż=.-�j�-����=��%k�"�n&������,pa���H�J=�8�&�rϵ�)�=���}<f����(�v(��-~ ��SK�/p���%�k�X��T�ڂ`_ܴ*��cH�m��<6�|� ������q�G�M�G�(4s��-.!"$|�٠ ���t3��!z��m�|E� I�Q�p�[��#����������>+Hj(�xg�*t����>���d������TL{ vqz��:h=�>�¡R��@]=�8Ѓ��\���"�e��w�z�^�:MRJ�J������L�v�\�.6	YSLc�׵��?�$,��o�#�=���c�f�����Ģ1�j\�$nǏl��ԋ���y��>��Ɂ�3�[hG�A���)��90�>�}� ���꜠�����?�&+����&����A���͵(^�*���u�Yt�Q:�pU��׉��h3H�s@Ĉ����l01oN��]AnR����$��4��η)�qg�	�A�VX'�LA� �S4��e���)�޼��mRCm!u���fkP3�E*#| K#���VV>0��#.O$( P!�a�젮�[��7�rA 7�聽 �R�eIk�"T��k���~���$P�.�3�"�����K�X��E�qLf��U�J�'Q�8� �sp�<%�ė����Ě?�f�ߌrb�`��~O���U���e�#�FS�!��*b^a'y�\�H)�AnBM�;d4Wv�Ƌ�&�ך����krY�ϟ?�^͜Vb�9����`QTbuX]�;0�p8�����aW�����I��v�P��  ��|� &o$���&$��ܦ��%��H��%9lX:U+� �)�� �抒g�׋�1�M�㴃�F��W�`Ɔ?�(*F�;H�#G�ˠ����o�~��xb��+z���,��r3Ѱ�Bl��}Yȭ��"H�� !�ћ����_$���3�8Q�� �J��t��Y�L��dub�y�d ���=fT���o
��Ft����6s�d��7�әj0~��F`������y���=<����.�T�?�ѶQ�B�v� �1�ļ����Jq��u9�z�C8���,��'C-E�р{
�7k�hZ�X=�P��j?U������j<��O8t��*k�sbw3���E��<"�D�7)o�VW-�1���6gk�L7|�����妖�7U������n+fu'f6ѱ�Ùz�^�֬��{F�F���6շ�\��;K�9�0���s	��K��^�P�q�p�R����[��e�;�1u������(�kRT~��qߡ���)l�=J����~���W��z��M�ً�����X6��٪z�w�+avt21��(�g�ۍ{Gq��	TJH�/�ft;q���ǜ��@�Ra����b:�u~,�=9XI46x6%����c�<гl9Pdˡ ���+�M��������[ ѡ��Jn^����n][�̖�w���ٔwBO�Q����F��c헔�o+�����*z�ѳ��3S��6�����w�|� �񟕇> ]>��ʘ �G�|��:�����Y7��& =<�T�q	�[8ę�����QR��k�!�J��Ƣ�W��n̊`JZDK9Gѵˋ:��K�Ou[5_`�$V(@AKت������{*��c�	���i�������^5YuY�a֬��XW��Pjl_}4����tQ��"�}���Q��Z�����5�]P�Q!|@���΂�����#�pʛo���T�e���Q���������k��Ȥ�,�����n�+�G���g�→o��4�.�� �����Z�_%<����Cn��*%��<'6n8��i3X�)�)�>������9��g�E��:SI
�%�Y���$����� �@����;�D��.��(��Z��&�J�߭�ӄ�ؖARQu��f]v�Ɗ��T�W(%}�׫�΅��aV|0���]@��%XU����/Z��N���g�?�Ɍt�i���\�S$�M��ʥM�p�fg�7�S����s^Mb3�Ku.���Q?oD�$U�{b˻�ߥe��¡&��UA�A�U�s��D��W�Z���3� �L^&�� ,=B��>�Z�x]��M��p
�Ꞇč+\�<�ﺪ�"f,)�حf��5�@u��4)nۈL���*:���Uqm��ׇ��MX
�{C��y�P��1��>��myF;�l��:"[�d��^�[�`yӛ�҅�J4{e�p�&�_��˛���R��CE����k�i����
��H5�#0p�ߺR����a�zb�������F���H�U �5�cvW.b����4�L��M�\�-$aÕ������u��C3���g�!WV����d/_�ۊ�5���YJ�}����"%{$#�'�M������\��P٠�vԪ�5Q �`�$�@��-)���n��d�����-Ȅ��a�:Ѣ��mWI�D�֝���6��ȱ!-&ܽ���ZS��5��4Q��*�T���^` �q4}
�˹%;v/�;_�#���C��F�����6��W�%4��F	џ�Y��C�yW�ݹU�:�%�̓��Xx~��ޮ�`����:1�I(�ϸ�uM�����l^�m�%P��ht9G�Q��0�����+(}�xWD�AF�H��K�[���N?���MRh���~�����{��
U���2�C_����C�#`:(��ܗAH�)tD�4t�pi��{28��l�W�%,;[v�?RӮR0	�5���L�~���<��T.�L�O
�[���+��+�ϳ�	� ���_�/�7����'�	N@�˲����x�
jK#I� z��L���΢B����k��f��$�sG�� ��"�f�t���FU��hA�.œ8�4���WS���Y�>�p�iv ����t/�",���D�����w.�=)�����r��&TӁg�N�D�/��{ͱ�u����@���ګ�Y'8X�Rw��]@���Av�KqL�Ϡ���R4d�c��,��y�X��eDe@�>��-4��ub��uAà�v�I-�k��5.6�X����A��z�Rl�"G(/��HM���Y\����7T)�@O�P˵�iOYV?%CO��x�lOz�D)�V{	��TQ\�|�T}R\���v/0���w���FE쀐{�@��w�������$�?޵�'�m?�����ϴ�g���7K|]�[�#�x>�$�~`�H�}�F�Әk皈��F���P߰W�K��o�L�Zj5�7`P�y�N�|3�^vY%}z��ϰ!�>_+�,�u ���򦽗_�ǌ�]��45��z��̤�6���K�b�ah~���9]����wH{ݞ��SLu@��Z���lqs=�-������@�u��+�LqN5�r���;QQQ4Y�����Ko�Fni]�����燪�V�*�	�/%Q�eҒ�VzJ~�e������9=�R�
V��l"�(�R7h�Q�bҧ鷓��� ���Uo�^�0Cv4�4�<�2�����"	��e�M�|�d�C�}���6��H��K�1Xc,4~0��(�i23���5�̆��5��=Ԕ:,Z�QxL�8��fXVU��N �ğmfm�r9��j��/�>�)Ca��ڃ���ص�l�i�!� �ÖF+���&r5��7���������<fO�g�g@5�T�y�~�����Bt�ݍenbϝ�M�jI8*��vfKF�N��?�C#��F1F�ĕ��2I�A�R݁��G
Kh~{]$u�u��G[��D���>�"Տ���:�pAy�l������5%�{+K�����ꊼ�Q6�sm^颇��&�G��d���J�i��6�E�V����Ѷ�(Jǂ�qa�q�q8Qk��V�s<1 �e��B]��<Mr�;k��8:/�{��[*^@9��P+۝�ZZ���$�Ls-�dݛ���	�%�[~J͋I��%q��Ƒ�I���fa!fd����0�e�J�z�{�0��ZG�`sJ�G2�&&e����%�7S�yW�SStXaV�	�a�Ի\_���OR������Y9��Kc�C���>E]�$���qc]3t�#X�ξ")*�S�~��H�c�^WAu証�n�ژ� a���|V>|�"Q��xԷ��/�h�J��R��_���>�H�[I��Ŷ5�WX��c�S{��*���}x�I=�W�c��<����f.�DA+�B
�Hw�ݫ��f!_�j�2�,B[����jtRb�K�Y�΅�!�__34�䀭 W����ΞZQ� ��Ҫ{�Z��X�o�� �|V޲]�6Lw`�Q�{��!H��KqSM����]f�1��!ըT�?U�C��<ؔ�J�*��	��^����]%��� �6��G�"D
���3�Umk�( �O� �}�;"�6��L����Q���,g�����Ζr�U[5	�>xI���$�_�X��o�I> �6�s�&Ξ�Ė�[��O .�9?ζ�[a��[�-�
�?��v���I4皅��TB�������=�G����uj\VK��UkG�\��Z|��;����+��U��""�.+,2���*������2��.�֫��T?��9%o$��=|WR�
3��`������m`�̯����M`zT0��6���M�04eD�A�'�}K�:p|
�1�d���ayMve��v�������~��-�>�^b�i�W�}مJ�֍�f�1V�� ��`5�
�+� ��ko8Һswr������@���^/�����#1�0]5�6��S�~�S���V!��5	;+b[�W��j��c���z��F�LM*��*>��*?r؉ ꊪ�1��������Q �=��n��l��H��ٶ��`�+�D�GHg~}ٻ��� ��/8�9�t��즽u1y�)e��Bz�G��7�0p�^�� �^L�_�+�$p�t�E�#���G���6��j��1 'cen��)�Fס�@,��z��
��^qU1�SOF��K���Y�N���9C?r�1l׀� l=K����|nm�����rw~.���q����۱�?��\���?�B��|���!ͨ[����%��<��9_��T��N\yU��1i|�ʘM����2a�	.vl�癇N��N�(3�Ĝ�Qf��#D�"i�@��K]��B�+�c�0R�����ߒ1|J�&3X ��h�<��<�������d/y�������4��g���ϙ��<��Nm��e�v������h��׭�
$���#�n�Z	�ļs���X_<�oe�d���EY��W�#IN�f��IȲh=�y�������a�3�Ԋ�H��S�֠/��"��.��n3�%�6�@�i�sN�����kZ�ɝ����,�ej�f2pT2<�|^,�8�Sؚ����e�PD7�!�K�V�٤��#}ܖ�H���휣��
^�i�N*`k��-�˚^u���/V��M�{*į&�(v(e��-j�ʤ2j�E���v;_��۸�)2�vmT�$ެd�����{���		���2�5`��g���fjƔ'����0�Hw����Ucl�����g��}w�o�B�D��t�\ؕ�V�~(#������K�-z+4�A�SLg�Δ��/��ϲ�k��U��Q}5�z8�ۆ�8�'�s�:N4�.�"=�g��e�������U<nI1���U4�����	����9*6�{�hL��;!E��Y�=�]X@\U��\���8@\|�?F�?H��o����@�}Ixz_T�#�9��{���#ѐ|��1q�ؾ�7�g��4:�~-`�@Z��
�!�A+.�H+;0�7��Ef�4�8^�~@��X��t��޴���l��*T.wY��
7_qvD��<2D�WR��}������Y���\����4�����<+����O�����ڰ��S9��F�v�M:��q�"ˠG`�؈�u��x�,��+�W�yIe0��K�~p7<�R�B[y�#J���o3~�(EO�ilW
�d��Rqjܭ��S������!�	��b���=O�G����k!��~��,��2k�r:v�S���f�x6W���Z�|�Oҩq�.$��"�}HRRC9��������X^�:����&ts$:ne�<�V�h/UG��~��@C� �{�NUZVB��A�5+&�m���q�Ȱi<�:WZj����C��I`E���b��FE\� ��o����4��:�C/Ɯ���f�'��[O��b�������:��h�?&܈���7�Q����d��ł@d���3����3w���k����_��P 0|L�Ԕ�$�#&M�P�����AD�	�*�[��S(���i
/[��G���+�����Pf�29��R[jOƌ-��@e�����o?��ҽ���o���s
)�d]���f���T�h=�L=毻�M�HOa0Nd��U��@(���eny����P��q�4r^�Z��{���oc����n���|<�~�Ԣ����@b��s�9U���a�$�;rd�]�� ܈�o��?�0'�ad����e���Û#�Fc���н�C/E��*��eK4;�=q��3ƹwb��EV_#��&�� ���H�\͚�Z?Ŷ}��Wj6&|����'���.��H�H�t�@�?��S3��1�ǀ��
��i���\C�H�j ��axeK-��e��H�5��M\#)��U�H�ɰ��<���h�J�OV*�I!��#��YF��Xqvr�k��;�मձ n���û�%�ab�5�����f�>*f�}���6�bmZ�rΖ��h0��F���Twv~�����R��|�`#oa��j�����늏��ƞ�X�o��d����)L��X9T��I�g�K#_ΣG2{��Dp���N؂W�VN��J&K���*��X�벿	
NMh�a�F#x�mD<H=���;̽����A����8�#�ث'y|ΆӸ��%����Z�g��+ы[�H�|�g�tgV����fH��Y�Sꭻ�M���mf��:Pv���S'��R�U:wS��b����a�H�(إ���lӔ�(�o��Z��\**�ҜȪ<1�~����π���N��znd�d��)!�iqC�ǈ�>V�W�b�;��;m`�V�m&�����ޮ�59��~�p=��N�:�b�L�Ӥ�R�'�?�W�8�*�d\���oF~����o�kJEl@��yi,�ILL]Go�D<�3v;	�Mzb���)�2��J럊��"�Gw����	k�>M���7|��6+�E�y�ԚBYLE�x���D+^��V���mp٪��E/��c�id3:l��\BZd�y[�L嫞�w�������X-�F�H��s�+���ҭL��x@�F�c�zp�/�w�q`���l��9�I�{�
���~�w>ػ����E��h	�z%�
M��X��*h��th���\��u}��hD:A�br�N�����9L�Y[싔���`�JEn	dEUǼ�X3�R����o(R�{@����I"G�,�h����	f%����l�P��c�^�n�	O&�B�I��/����"{)t\8qF��L8��R�v8u	��o���_n��b毝ivݡ-]͝��?z��)��z�����z`��`��S��ط�"ܒuU֫b����n�s�>e����!�8NHIS���(���D*-�	�j��^��Y��F������n?a�M	+�A��ew�	�<���*9C�o�,{����]��d^�HՍz�����s��|���o�=^lt�O��XGӶo�;��Id�1�'�`^		̺����r��!Ap;R鄬�(������$sn��[��*�x�s���5F �/%ہ濥�jA�<
3����J%zꀒ��l�]X��R���/^_o㮝n�:���;�qZ�VN��Q�g�u��c�I�=σ�DM�~��6r@��O�	uX9}GP��qlCx�\��Esr@g����0�J��S�Xoz����H(򹻫�����D�F���c���`z�	�� Q�p�RC�����ISQ���3��]c�O�M�+s4S���;	u�䇝�����ԑ��sf�x��ihe����tҜ@$;��u|�2�v�	!�uM�].ac��о6�G�[������C��7X��
�t�v�,�6�y�����N_랷a�g���F�f��{^���ǩh���d�`��n0'gd�ƫ��P6�0�t���:�D.�)Q��x(N(�%�_���L}ѩt�#H�P�T)(H��3_�b1�4�;�E�	Y��:�k%�-ըR��(���w���x(T�nVj]�s��bb��/"â�T�=�=�լC�U� $TD�{.�H�D��2��4��c1B*�w�Yb��C�������}���ͧ�7��[:�� �U�Mh{�R���__��-�bٞxg��1g(ͼ��8��W���#�Zx�����A�r�/�9rg���~���/�7t�MZ�c$��R�q��|����Ҥ	ZY1�S�Qݮ�x�����K��q���OY>}�ێ�a�.��7�eۜ�<��;�Ӽ{A1���t���1HX���>m$[ͺ��{/�.T�{��L�6�~J��Y��i�7���k8'�����TR����B�< ������_S��2�
ʘA)0W�
�5�>!����ކ��s_R�#�%b�Y������{�i�,�=n/6>w>ݘ9X�O���T���8Zf ثc�QT������X��s$�{�f������p��T��u��5}���(�u܏�6�W�(Ġ~�c�Dt:L�٭��t�
�E�� ���Ô�qM�-N��]���&m�5���Ԟ��o�m��3�m���+���_|M���'M��
í	�'l�|�Zz~�
i�t����L�Om��|xjt#��}ĪoQYH��vA��Jօ�j����(N7^����!��H �&�ȧH���J��Y~��E�-����(��!v�9[qGH(J�}'�!D`��l�t`�"�
BZ,{"�u��a/7�F�`�9�����=R�"��*u�?%X޹Z�wj]��^��'3�e t���5w��X�*�]���\��T���DH�[��LE���|���3#�S�WW�6�� ��G`,�hu�W|1���)Yꚬ�.Ýi�2~��!s��y��q�cHhGK��/(pUO<���:���p�V�9�K�����z�rQE����gvA+3\�Vk� .T���Ob`��0o'�����b��GNcg/A��/��r-�+l�@_k5����ZŚ���Q0�/Ih��F������wT���?PQ���Hd���	W�k�h���:~H���3A��`�eZ�a���>j1t艰��M<�=�.t�zYH�L��H\B�y��㌁��2��B;����%?�������c�`V%f��l=�r�5'����P���;ڸY��23���I��|A̺������$ynE�����^�L ��R�XF�SF�M#��9�gF�A���'Hew߻�jx��5�B;t�z�!0��ܛ����~�,���_`�W��2G��-�����Ȑ~��Z:������ 8��EGvX>��x�l]*�uU����Jf�+����}�	ܨp���w�aL:�D�l�#iDHm���N����}���H���+u��a$�!���{l�D�P"��y5`;{ u�@B~�� �sy���u��oQ=>lm� �ґ?�4�~pS2�[�Ku�k���3
d�Gs�;N���ʕJ�`;�a��1�Ǒ)}��L���PR�A ������;�T�&��X"Z��}�����.�U�JG�p���
�;�$,����{}�l��3	)�;wc��=�e�ˊ���ԫ�['�;����h����*Έ����[;�s�OI٢���˟i�c���L��t�����|�R���7�l�v�nzrC�:�)�?2L�ի��%��� P��*V�8�%.$ �� Ph��G����f�{�9���XlI�ʴ�hyA��~˫�h��W���=��Cm�� ��$�s�>�Uڿqz����bU�$w�!̓ͅ�-�9�d.n1?�C�]],�h�N�y�0@�cLeG��y���ެn��x��q��| -PB�]����ɻ3���e�.΁��0�kM�,�+��X�_�>2�����0�d/��4Y��Y.��j/�)��o&�������$��8-BǼ�+m���e{\�SS*��I�-$V�:��B��Zx�}��&����7#��'��(Y�������Szq*���Ԃ�����b�
���G~<g��@���ͬ�۪9��Q,k���T7K�\Òp0��'�qΪ���\Pzov@�sS���rX�D�ǽ�5�E�K�����f��v�#@4�uO�Q��U1?�X��}GCN]6L���o�U��.(tx�31	���b�6r�X�B֌4Rn�Ũ;�<��s�b�Q�b���b-���YnK3��7�	M����_�Ϧ�j[*���("@dX�����<�;�7��T�!��C@�~�rj 3+��(>�86u?lXU�G[&�I�����qzb�8P񙈯V�TY��BW��,�PEŮ�e�o���D�.C7�W����M]1z�G��l�J�s~$���cW������6[��Th�Bs�donP�o5��O��Y9�AUS9�L�<=n���C�J~X�:�$�(��f_���d;���eѥ��x���rz<�q�2&�`��j�����j��:ś�С�n-�9rY�?�5c�@v�P��N�k�--Z�,ܣ�|��a���?sڔ�Y\�e�x�+5SƋ�o����g��!�Sd��
rsHѽ"J�����C��T�ۀ�}	4�Sx}�����U��dKM�5K	��{^�g�]DwZ�Ih�S��iSL�mt��8N#1���}�1���3�w[2�i-����e��7�u>&� >�s���$Ĝ~���hE^u^�s8��P��>]x3Tγ�N����'������}D�o�l)1F:�_Ue��Z� J�y�KԚH���?�t�ܛ7�����ՔW	עޅ�]�TAL�����E���I�d�#��6���C{�\#w&�tU�Mnc,�V�G��>���f[zF�yl�\�5��}�#�;%�vys}cfot'#��n-i� ӿ(��V�VP�j��1�J)ߵ�4����X���Zv�m�"�jq�z_�zLL%���]!��If:��Y^��}��ԝ�ቒ7�f����ml4���L������s�&+4��㷟U�7�D�m�sݽ+�T9��`8�A���F�-Y:R��+P�;�+���˃Ek�����v*�7���0(�Q#�(���f)
���?��P(�4'i�ϣ2�L/J�;���i#?��Q�W��Я�A�V�'����+I�t%>��2ث��v�|Jɼ5�?��(��{cɂ��
?��N�rK9M���q=Μp�Omv�ː���;�f��o�v���Y�:���9~��$�B�<#[�~j�_j7�� -���˝a���1�w��^�Zt�1�L���{%6_h���ˣ��݅g0=)�p?��q��E�X��[&��K�Ul�[���0�.��ai��%%�����7҇�V,W��x�����w����1����8���)�72�=G8�v���o/���pE$3\hf���Hv$�%�z^t��i��T�)dC��N���~��=�x�G#�#M4.!u�Wb��S��#�I��3"[j�l�m���r��;>��GA[��X�B�Zje��Ud(���X��6!�5r�� �*5ӊ0�x���͍}u�����W���#	 ��xc�Z�O�~�A��3[���))Z�j����vm?^�WE�� �u��8�<vpM�{KU�I�Z7J �{�&��<���n`�L
9;��w�����q���� Y�cs`$���P��S��pMD}�Z�	,zy��L��IbH�I��BH���4#��2�[�.\��]^Y�#H��t�N_�"���\���\��O�� ���W�2�����zU�mB�`q��z��N�����������y���n�1�I����x����iw0G�|S%Ճ_�O��&<v�dTsݯp}�0�|)�*⹹��|���ה?8�t�G��ԙ��?*'�ώ�~�h���I&^��Ww}�Ւ�"bMW��z���E4vqBu��=_<��=��q�-Y3Oȟ�^fT F 6�8=�Zm9��z"q�tY�iT����X̷d�n؉]_#k�P��t]H� �����WAC�R`�jC����u�k?z�1|�R{.8+��T�#'����*%���,U�y�y�i����v�֨�f�8�ZR��`�U�'���G�J�]~�� =vs<�q) �#L�j".�����p�6�*՘���(���l���t?���i���W�K�G-?��X ���EUFW�|�7�^ M��k=�	����!7 ��	�s}C;�MV���4B�oDDˮH��<h@bjn}�4|�_
�8�n���'8sc8�u�Ֆ��<��GN�Y� �O�~'<a�ɂЏ%�̔��%W���X)5[o��0��+�^u��-�]���>�ؾ ���K�Ji�?%@*�#�n?!WW�O��F#�Ӏ�U����;R���3�Ɇ�l��;q44�SҪ\����з��`������V�r芝
*�&Yhb��\+�f '��vO�
A����7Z��u��~���A�Z{aS�|`��V�0�~%Y`�@О���+`f���@�0%�Bk���x
�IY��O�25�Mt ;k��J���j7.T�'�dۄ�A@�h⬀�0���ne�jDuQ�έ�w�Η�C�@=S�PH��au��P�Sub��ZN֓C:�^��.�?������D8_�ļiY���ق$�'��]w����|���R��xƹs6L�����P^"���Eo,DWG>���l	{��.�Ƿd�AXߘ�����O,�s��-���$p5����:�oYvj{?q
�q+��uHe���֧A�|3�Gt��J�8$:Rs��f_����������>9;nS��3S�SrN4�96���a��+�H�jb��L��J:��5T01&W�!Lc���"a�皂���>*`
�!��M���K^�H��ɜ�$�s�:(���b/���c�ۥH$@rb!)�Hv���X���mq��J'6��4R.�vg��f�� ����L	g�E|`N-Ɖ�@�vN?}��[s���u�C�{��f���M�Yb8�g�j9�h9�/шցB���2넝�@]jڼtTGIF��z@����E��F�@�����9�,��t���8\N]ӧ�8\r�t]�O��LʸS�:�P�pY�Gu����pn�:L��f�_�R7�$��m����W�X��1O-�g��ϿЕ�X�`��py��UB-���@�Vy�#�=:�(G�x�+�v��~6�v�[=�ב�ᖨ� w�bi�:����r���q-օ�b
��d8z��,�S`,�+ͧi-4^�u��٘�C�M�W��l?&q��4WW�"����(*���]���X�&��Ι�݉Q�P��1�{A��Jd������(f��qĪ��CY�z��dm�!nk������&�mC5��f�D����s�=�� �z4lˋ�.H�Q��b�S�K0��'��C�U]kl�.�F�E�[5I%��cD�����WIy�<���zGʴ.�|�E^��kB�����C&#a??��������2]R�G-����@���&Go{H�ANBq��h%�����
#���{+�N���0zF;c�/�v5#��5�g�g��c�P�K�H}}�
�;dRW� �u� �4�ͪ����aQ6��~@��{?K����X���SJGj:��d#�\[c�e� g1G�4���j���`�B�l�f��w�v[ ��Qu]4��������g܌ơ�ߧ�і�`�� �w�*SkKC�)���'�.�X�|����T9xba����\���_~���?��ȮX��G�S	���߹ڞ���i1��j:eB�qI4C{{<�DGj|��}��J����)�Fo]�9�3՝�2�1Bz�f�Iɡ��� �A��~Za	�����a����_�`yQd�
�uW��(��
��M%�H�2�#�֕��XRY��fi�]����Jb��M�[�2��/ &�Y``�� �gO�������n^MAp��`�O�L�y�Wߋ��`Na�G"�2i��jW@�����P����6��lu0��s���,��>nJT��t���a�F�t�Qt���P���EZV�T0]��/s�b�����음3��C�ΜG[x�Z�h��?�U _�r�;y��ye�S��ӳ[z�L��jBe�ج�'6�Q��t��2R��b��h຤���"��"����
/[�7��r�A���7\��.�7���� ���b�2S�p�V���3���=��=^�P��՚R!e^���5Cȋ�oh�S,�O<�ߥ��,����;�������&��iF��@��Jޭ�q����Ln�ƭ�@�留��}
���dN�AAb�����V/3�#O�-E^.�4�t��H\�3��
q��~�LD	li��V�%�i�����0��ʩE�_�L�pTNȿuk�*5�r͓���鰣��O8C���3�'T�'EA���p����tQ{���̩tY�Q��H��+�^zXL�,$}&,�+J����Ƈ ������$���;4
�Y4&wͱ�?pl��mLc�G��)yB�ւ�-"�#EO��*���A='lB1�C��G�k��&Z�$�?��:~�&�r�{y79v|�|w��d^i�$�0�=��T�A�	�9�p)tH�ip:D�;�	J_��̾8.�QQH�r��� ��R���2�j��(���J��.�E��f<�)�,��~����^D�P7���*l�ۻ�ڣ	/{x�<�mj�+uv��i��!�Z9y6�H00^�0"Daoe�L]"��$�I���Y����M���rm2Hu�-�Xh��QE-A�-kh��9Z�ðe2�?q��GJ���Q�SroA.��8o%x���:��;�����t����*;�B-�v{��c{�ӓ\�؃�:0�D�>�}(��m�z'HS�B�B�27�� �Cg�w L�s(&� p�m�-F�F��qG�TL+�zv ��)�֏#X��� lW��֞�����,o_�T�}�����G��x_\�gH�5��8��+�l�_}r�=ؠ����,��ɦZ���4���C��[y>�ڞr6�u�h��zVwb���e�|=h�3�b+�fK(nF���N|����Z�@��ҿS�I�~�w���Y'S�9؆,9�7�<�/���.�� ������W�U�!]��,|o���f#m!ǫI��F�{F�i�Iu���^0�e��{,�M���ƪ@�:��$�5(d0_3đ_Ο�[N�T$��,���i�ĶK�+W��7O��C�|V^��5���"Rg�{- +�zC��]Ǿ^�8���$�  �x�1�R6B
KRUCi xN�a̐�lgM<넵��ٔ�g	6L�$V�*��/I�4�4�� ����[GJ��}�/�v����	�0̖浏�h.��Y�,W����.c0R�߯c/o������*|�7_���7�L�b���N��/�g<�a�jmO�������y�(FU���k:����"�#�w��D���I�%���\�]ƚ��kXN�����;J��XaeXO���I��)x���1��V���XԐ=�{�`��_��D؇�>d���� 9����5E�k�����x�C�+����0���̕q2B���Z��+��:�^�� 7���=-��[�N�|j4��'Fo-�:q	JPth�С;LU�?��] b���e��Y>V��b����P����vZR2r}S0��?���6���7~7T�g�ZY�=�a���O
6f�8b�9z_�r��'!���K�fO��7����e�#!�+5��Q����� ��E�b�[�p�{�1�YR"�+��b�� *X�"��IT��XI�"�4o�8���;��%�(oɴ�p�(�cK��V��B�>�v>^o�;��vOg���6�&�&H
\U�rs1i�d
d^��T%�jw͏�ď'���j�0�!��b�YA(�!.)n��L�����N�ݡ2��(��LQt�m��l�Lm1$��2�g3�_�Vߕ/��86<���ۦ\R��}�u+)����-WW�u�2v�lgۡgj`^pϱ=�X�]TB��B���Pw3)�����	p�ĸD�������Y�ڟ[m����Z
s2�=���*?v��В0��*-�V9�2�C�׉=R��cA�M��V�mYhŻ�mۑZ�Iȗm���`j���(Bc7jy� �x�[�{����1��۞�'���C;�*�uSn.�A�8d��D��K�~��A�*��LO��?�vF�r�~z�+�'=o��l��o7���"P�E6��FQY%�9�id ؟�wׯGь�p"�Hy�[�9l1F��N���^.��~�c�����aS�nF#A��D��^��%Y.� K�@���R-�eh�Tɣ:H�!i %#�蛱p 0���bi�"C�rܝ�U[D
������8�� ��Vͼ#F欮���	�'�V]�9�Ϊ_F�$鐱Y�ۡ���Gd,��VOqB�����.�*�`�r~@:-G���[��&n~=
�U��Dym���n?��cv������W�&��2={"x�R	'���ڳz�+�� ���/��q~�Q��EGH�U���eQ%�� E����_��Ӭ����O:|�ڳ�@�ِ���[!1/ ��T^��q��iI�V��B�A��G��4��K�5�']�\���.��F�^R�OsU-���Z��=�.��q��)�G�C>�f����Q�㟩��r ��V��)��J�2�˸����2sa�S���<�uD�׭������Ɖ��ܬ
�LN��-�W�p1"+1�P/|�6c�M+X΅���\�r0��̃'}�k���yT�d��n��aR�{�B��'HM��]��Ȇ�g�$#IK>e�͕�[m�i��U,+n.�?[U�ZJ5Q��I�9��{���I�qY�т�d�T�D"�t����:�����!� c\�{���j�����0Ԟ�U�x)ȯ�(ߔZ�i���l����5lE�Q�]�5`�:��~b����߱95�a.���y��̰;��'�Wt_�]հ�lR{D\��5��o|@�R���N�FQ%Y�X���o�C��p��7�^eT�������K,8�� EN7���W����5�C#2���Ǧ�y����+�J��>�`�{a�̣�ŭ|�m�}~�75��9��
E���x���R�J肰�F�n�6���5F����U�Q�Ư�{]�VϨ��4{aM���ȬPJ��x����o!�a��?��%���)ct|ʜJoBMS5X�������s��L� 5��B�+2zk��5BM���� +;*�;�j72�$]�B�s+$J�[	����2W/��OT\��u�Y���'>�6��/-�K��m�	((�P�)?�%�^"����*zz��e��*��Vg�f������wt!]l��)@7X����c�r���K�د5�^)��B�h�2jJL�W����ey���uP�+�C��pt��FC�t�_t$���#CP���Ѭ
o�3	O�u����꘿�#VH�詩dǂ���&�X��o(�L�w0#�V�G�>&9��J�H�CU']Nva����.>#�z�}b
7r�]�^������d��-�@YZ�����f�:j��|����B(��/%����#*)�����8A�1]� ��9��@m��h�%Z�:�DB��<���F��F^�QHR������������"D�&&��H��Q��a����.T�r[�6:Q�h�\�YM �PF�ަ��m��J���&�!�'�@SC=�H+P@�b���p�_:�C��>��Y~̍kܻr:/���,P�8A��~zeʊvׁ��:Xc74�f'��]Z�����Kfe%	�c �ŭG��p:	#)FU_X�5`�U���q��U�z]�ğ���xU��R6L_��<q ������\Wĉ�af�F*��Sc�y;��ld�m�(�2Em�8��Gng��W��Jx]�q�X��b29������_5�(����c�j�-eY���@��w����N.c �qUڴ@��n�1=}|�q�j��y+0u]P��AQ���+��]�U�i��x���4��+����%�)'�H�1�@�4��L�(�׮� :9E��-ѰF-�,ŌҴ"0S����:��bB�s;�oɨ?�����\�9ǻt�a҇%Y���Ef����f�j���D?P���IηVU�)����^�q]���)���3��;�AH�\��m�%e�{
����/_a�ɧ����f�΅3o�2�ϒQ%$q��jǹ��5��/[u|�H����i�P��x+R�U�L�3?��G�r���=.��!���?����/���"h39Z־氟0�t��<f�	GG�t��L�XY]��o����� O�����[�Ry��A� a
�|��~ܘ�d�����=G�#{*p�`Ŝ���8����1���ߋ.wj�/Ja��F�*"�6O�f�h<f�,l�[
�� t�
9��xA���m���L��o!-n/Sآ��E=�5f�ْ�j�����ƪ��4ʬ��8ge��P!��x-F�[��H�K(�:|����Xp�@Ҕ���fcF�է^��i��!��z�KC����w�kb(�q�r�5R6f�D���Ӵ�gUh�vb�d���o��s�N�/��G�ݰK��F~�]X6��Y	?��ޑ�FFS^�/Bm����},qQF�cs�qbd+_�g)]�������( KK�[n{���6�;����os�(�c�sM{j�L� ����#�=M��Pa�"r�>��w�п��P�1�y�.1@W=�$���X������AnP'�P�ٳ(/N<?�散.L�2Jt������;��dM)M��x���AW*�i�	.���vz��C7�R�0�'Hf��gӘ��K���vF����K���Wϙh��Ph���x��7���*G��X�W��x
|>�t��}��M |q_R:�|W�F	�O=jR� �!����Q�v���Vf���`�S�dt�	?�����!��-ŵ�@�J�u�h��������%gf��?M��>H��x��*�(+�vbA�&3�T�eQY#��$պ��@�E�n�(��?�ƨ���h�k�[���?�+D��è�@� 0�oÏ�$� �N3I�g���O��]-κd2�����u#~/gw �`��I�[y��N��w��X��-��<�i�o�GN�_
w6�.�Ǟ��Xh�\r����ebn�$8R*��eR�6�����J�F3W5�g�M>H��F#�I��B�;0��YI�x��P!-v�2�6f釾�P�ؽqYF괥�@����>����(�?�n=����ozd! ^]�mv?�S3<�ێwc�R��:�g�;�B��,�ږ�2��{�mF�<qbh�]��#��@mE?�QFX�f���z�
\8C��.)��5#}����-���u��
����Ww3e���6��J:P��@�?����?�&���>�D���1�N�˯�n��t���"_"#�b/����7So���1>��J1�y`B�F������:��tD,Z��j�3�F�n7̤��#E�rM	Jj�|E�A2�Xb�<��CD�����S]�U|*v�
�v~�ʱf;�����ɛ�����xACZ�S�1p�&��b�[,��!Ji�T��VFf5q�b#b��Bh9�{��J1�9�@�����'� �w�D���T�>WC.9���py�������Z������r�&/��*?Nj����i鯬���-�w�35�f[c����m�����t����1Hh�1N��Q+�tϦ�*d��91�/�$7������$���z���ǹrs0ͬ�dշJ��-q���A��қ,����tf�gN�KK?(#�^fM������y��]?z~��2O�o���"��;3�J:��
`�����W�d>(�G��U@���6���}i�����̔�� ��gJzn��TAD}�c���(v����ː��11=^��l�n4����{Q	�������-R\��N �-K�j a�$�s'�W��N���S�2'ZwB=c��v;2)�4e^+?�<^��9��<ɨ8Iʓ
�Mk�<Ӈ��2�I�G�D�6��l���zC����2�|�狵��Ͷ�I��!ݮ�֝!}8�r-λ)�;�܅u))+'��@fU7��.��߳y<|���֤��L����>���"=t��
$�i��ėڃ@�I9!���'���9�6z��뛨��`�ݕ���_�g�/�VU<��I��ef2~����Ү��B�d�? z���}�ذ�k&��7�Ar�������cH�=OQntVGǥ>�{�BKgczcUrVX�����9�= ��E��Nʓ7̎��o#~�6�ZVl�x�7P-�EG��e!`
��[�����೙>5-�q.;������	a��f83J<6QH�FG<<�#У-;C�oH/�Q��,�{D6�>���u[��Y��fKuG����ўLf\y��̅�����E�v�ЯO����; ���Z�	���ڷ����s�S<�/�)ɷ���3Wxa� T���B']i���u`�o�^2Α1���"�O!Z�m�o6=��n����}u�!؊ϫ�3��8k�
z� ��1U�1ӄ���U��M�u��C_�"Z�V`�t'��
�(]D>�AK��I��Y?E�0�C f���YJ��;���-���ՈeT�GBvk�)5K�+���h"SR8k�}�S14a�4AM]�Q
K�M�>�9�:@��/AچC�Q�$�[_�U�⸗\���,1�Pm���V� *5�]���jQ��% b�x�+i��~^ ��<8���w�a���m9�e~����U��T�#���2��5�9m4�Q���Ϊ�ۛL���*�+c�b�τ�ӣ��'�f�}�e�+qR�.�Ŭ��0�5��eka{k�L3<l����z.��7s%��%o��V�}*?8+8�ԟ$a-��B����Χ�O)���6"p^ږ1�+,��pϫ[%ϻ�L�y�������g&�˴�3�g���)�;}j+�[���7c��������_�Wa�*.P\<tBz��-\y`tDr��s���F��R")���z9w��)�r��f�t�VN���*�t%��|�v��s�T�t`����t�Z4��ke[�5\LRս�<��Y��M6�b�ʖϖ�B�1`Hπ���0 X�{�k4���[R����h�9��C)�{b��lU�y]�*v���&��YKAė�)z���#�_��f���QO/Fi��%�Io�'�t"5v&B�0��*�O�t(^
-'���n9���D������C��0K���I�����U��P�
����1.H��1�#K�G���Q��>�zK�ļ:��>�y�p���x�0I���$�[��k��+%�T�M�~�Xd�N�	��1*}>Iɤp	O��a��(aY
:��j��ɎR���a4���K��Lی:g�z��r�_��<լ(1�(�B`3C��4Q���-d{g���]��=$��~:[#�'=��vD�%�~b����k �H�y	��c.��7��0�"�s���@����2.	���;�3E�>����� ��@4����l���	hq����v[��A�˞?�ɚI���!8сx��̏�sN�ȑax��)�F�`i�*~�Ϥ�#G1=���$�s�G�]������g��F��Q�7�S������=�D�(7�f���)K��Ƽ��i�Oh�7Mk�� -b|��$$���@��,�	��1���$��Eu"y�.�k$�$�{�� ^�X(H�!<��� 4`�-VӍ2m@)t��/�쌿��o��F����kw� F��v�Iめp�I[���
�]Ăaw��3�
�X5�,�]DZ�>F�Wt���"��'��aɬ�)T��{���B!����iQ���%-���AC�C��9#�����eL`�4��u�!�Ban�Zv^ݍ�,�3���eLv��H�G��m��GI�-uAb�#��� +>������v��s��:EWMS�}�e�Kn� q�Z��}a��5
 �׮8W�nᜫo6�ƹ	>�YƐ�4�X#��j���9�V����\����2]]�)h|w�r0-�D�zq-)��o�r������{IG��koB8���,��Fs	Ò�����os�O�%KH�T�m7��}󰳀�������F��"�R�|)�U$
L�'Ki|�u�4g��U6���D*��,���歗�%�s�Y�1H�?,j�̲������Я�B�wr��H����%���V�񝦰���J�V:�T`ju�����b�<��o�,�O��M)�qH��@��s1и�g����;�d���:o>�d����O��l^�&�X�Ԡv �-7��f_��B	#�6S@9$��ȢB�ڜ���Ry�\O�¼_��K�fBt� �N���Ĉ<n�5 as��@�+��j�L0�K۹�O1`/�a;�~�'�����yz���rv�� �W��`>�8S�c�kE���/�T!B����p�z�� jh�3���K��HH��(��|��q$3_6$��cA��g����J�NS������t��nx'��8����e	+����P��	��ʑ�Zz_�BO&A�",��H��3�V/QW{�H�q��6�bv��L���d%�u��R\F?G��Diő~�<毷��42Dx��W�$=����e����5]%l�-�g	U�8������j"��2�V��K���?GI�m���97ǏL!K��|1��z@�yɋqU@||�/���^��������K�z�\0{k㚆��#ls��*e`��+*$�����P�n���Uؓ�5��"Ԫt���:�b��T��>U'������0��
��w�E�W�r�Vy%���}��!�gj&6���rP�T��y^a02��ԅ�y'���������g(h�;�����t.���e	�:A�9h/��6%�v��b���ِ��(L����i��pÆ��osj9Z�/	�! �
- e�{�;	�@2f��ε$�}�.��T�����R�[s��B�K
�}e���`p�4������#�3�����X��`��P�V����/2�+%��[�6�TW�J#zɶ���'�
ݸ���Ե��V}�H]�L�5ۘ#`B�VE�9�?��9��t�
��}'��;�e��Z"L��@J�f x]�P�HQp��o�]�1ue�Kw�I��=� C5F�m:3���
2a�x؁Nc�	#�{�O����(���C�FV�!C�( ��QN�b�y��N�-���S���%(ıi ���Ls��x�h�^�9�w�;�YݵP�-Z��ц��9��o�[����)�?A����7�����J�Z�v�Ot��m5��iP��+��'x!�V�ES:�'�wx�+�9�Zi!b@V����5�ƓE?��ʯ�/L�r�j�y>x�2M�ގQ�g�ֽ��l�x�}�8�:}YC��Al��Y��y�����i�|�J}�^�pLh�W��T2S�;�wv*���٤�$����~)"�I�bXCI��z�TǊ�]4�6yuW�\H�Y�R����j�����+���U�jWT~᫅"eq?r۸2Ze���&�B�*�d���öLP����6Y芾b� �k��U��Nq7������@e�p۸�$�均��}F<���߅ڛ�]�eF'ӫp�v�e	Y�q�rH ')��U�S���(��å�x��h}��	>�v�}�-�$ډ�l~7d,0�n$���<�4a��������Ԕ�"Qض}بR2+8�_i�
�Ӫ�H=[pm���}��X���7H�H��Nu�bEɸ����� �����B��:�[��0\5M&t����M��,y>q).}s�ѝ�����0/��yX����C�^L!\��(M9� ,yg�k9���3�����}۳�Y '�G����$f��mb��ŝ�G^=�7(���[I� 7����J�#�|��pf6�<Z:#��ĘP�ru)���q�K����}S\�����-s����¸wXq"��WZI�����޷�f.,Ku�#c��2��g����)r}���Q��4�ľ��L�D�y�
�,ٖ������1�R��^���$ /��e1�CO�������`��߀���q��8���������Å8UϤH�%���&*�+*�z��M�G+�f톡�o��;��ϙ�����`Ϲ53��rBӌ��|���v����s�ɧ����!��g�'n1����z��i7,��fR�� ���<+l�p���I�[��B��Ô�Ad�bӰj7�>pN
z�Ᏸ�m�A�,x�N�.>���IJ6K�d�>�_,�F8�S��ǫoC��?:��]�}���X��޵X�gy�,����,;�FQ�|^x)3fEiU\�#rf�/�-����ő���Q��ӹ%h�Bh���h1�o>N�h���&h��a�Me\Բ�	��(�^E��ɇsqD& �>�Ä����E���Ãnّ�/��f���6Q�5����i��`�H�K�F�3��Y�8(w�����}��r�	(��Zww�/�ub-�no(�J���L����ҧ��G"�ã(O�J� �=+)BA�7T��ԓ�\r@{)�[�.(��vX�&��»a�Oޙ?������ar��aT�ꡊ:�X�*�Yza.h�
�ݦ��`�	W�f�9���$j(�o�G(�+@z�����k�0�3EW��c[�]�۱i����X�S=����fL�4��>q�0��?�қ��$Į/L-ayI`�O���V�[�q�l��d����t���1t�e��/�w�wE�8ø���:y%FbOZrn�H�k(q�O�f��M3��!7�&mQͲ�T�Q2{:v�k�:6- �`�JX��B��ԅ;s(�1���	�Ub+��߳aBV	,xK��6Gϖf�X���oΠռ�\��3@ˤ�l�Y*4�$�����|�Z����>�/6s�'�i1_�*C?V͊��d��@ʹ��Μ�����㣤
��.�?��2� ?bg-=!��'m���Z��Y5�!���9깣/X�5+�8��ݔ��94EO����@�>��^C�+Qu�2����8q�d��Fʴm�@<��E�m���AY9$[�)j��"�� ݆�$�*L�c�z���b4���e�T��ɍ�Q�`X{����Ӵ�+6��߈i#oެI�k�W;0P�W�w<��F��F!-�%�[�D���a���]3d����S<ϣ�wo,1�{�|R.�[8 n��ۨ�K�M�_^�a�_V�5�妓��)S�V�U1��g�+���$����BD|з��*1��S:�i��Np�o�����?'	X>���S�b$�?7�ņ 0���IqK­����Y"�{�˔eT��z^;�l�Q�O���W��?APR�_[���tSe�o$4�\'�_�J���C��K�!7M_�n������)OC�	��]��.W� *�q/d�ZQ�T��5��@3t�C�~\�����2۹4����D��5;��Rz�1��7�|�_,�X�y���U�sE�/ct8�:r}��*�}���+�O��a��2⠂ V!L1�K$���E�K�c9�������7� 8�9_�9��������#֪����?�:s�C��B�s|���/��%N����iwQgmU��`��^3��QP)r��&⑸Ɏ̜��9�� �VEa|
�O5x����:�h���sQU��o����-2�,I�>r��n�n�ڝѺ+� ��NL�KD��k�o�UDBu�� d�g0~�/���0� ��H)T�HEA{*����O=�{bw]��%�fUyw�XJ�P�����jJ��B��5�WFa\�K*՝���B�&܌��4��/���8xO�\��.E����јV���R��>��#h�&����<&�F?������z���5ۜE��H���D� �#1�K!����.)-�pteGf?���.�X�Ů�F�������
M��x\�Ůi��8��٘%���ϱ������ 4=�������:��8F(�ǌ}��^N�v^�Z,JEΪ��oc�tͧ�� ��EEI���S����U�>�
�El�M.�\sA
/��$�ۻ�/RƝ3뉭[arr3V���w9\����aT�M��'%l������>��ҍ���?��smӖ��i����
Y�:H�+��(f� {�p��mقpy!���Q2̛Cϥ`#�L��x�j!l�1��*h�3caS6	�kO;��j��$��rP���VO�m"�|8�&V@�m�ڣ*�4]_�GT���=�A��G3�vA�C��-��r�g�X�{�1�S8����Y�] ��=�,T���u��Uoг�l�\�Dd���#����p�yJ�C��y��)D�5��>T-�^�ҍ��F�+C���`��ϒ��Y�2�����D�ߴ5�����a� 탗Z��-�̷�=��5���!H9���	\G1�|����4��,����4�T��Oɛ�\��apa��ٻ�늦0�\|�MT�G�!��\���E�A�w��p 6�d��\Է �	��u���Zk��� ���-~�����p�*��K��B�$�d
��h�^�˞��u8 ܞĆ�$O�26�"�`r�W��M��٫�$"*��+���QXo�~B�D�߯:z��8X@![�eYI+@��ӁMK�{�\S|�'���3c3����z�F�լG���y�ϸq�D� ������q��|���"<�aJhf�Ĉ��n�%I�A�HQ6:���č���|��a�AmI:]���b<��8���"6�����[u��0�X/U�;���m��^G��ZN%7�=���Ќy�w���+q�yZ-	!϶�4��WΗSl@x���F�LPv.U��$��ϣ�ix�'�����3v>,�H:�r�ݡ�G�s&6��w#���P��o5n�{'��x&��iQW#@�ڦ�/��&���}�vo��r�yP���94�,��M~%�9u6��20�Xk�gNK��nX��A/�=�څ��~��a��$�zWb�x����k�8Y�G(�v�=��ӛ3w���"� j��G��D�O�/�5$Wݡv?��tv=B)x,F/t�Ҋi����E��X�Z\��9��*�1ѻr���ʣ�<�|#��1�|
�w.���V�?Xس 0���!�k���#����a��ڬ_N� vV(��/-���3�с,�G&d���ۆ��_g&��;:gx	6�p �z�&���M�x{�0�8'�Qx4���31H_�aR��7K_D�x:�,�J.�WM���J%~	�R`�5KU��1�tnE�"��=������w��<AG�d�V����<��.�����,�Y�8�w$;�ZU9��-�o�o�\~\��[���{Ζr����p�8X�W��q. k���ο�!g�ɩZ��ea6�J���Q�M��a�Wߞ|%�[��>�gpoK�C伐�ߜ�HO�����im�	������L�:s:dܦ�U	J��ґ[UAY�=WJi!�
#E��?��OHI�LD�Џ�ꕗ1�m��qo�@��4DP���"sP���J�#�]���o��A��5IH0�P?�xz���h�b=`�T��<w�M\!�Ea�?����S�Ҫ]�Ԃ"��p�g£K~iz����.Se_]L�{��-hXz�oߑ��!3�whԃ��?�l\ �Yj�E ��?����~�p����@��=oL���t?�@�i���-m��e��R���>��3\n��l����!��Umze�F�tY�P�G���o"ޤ]���(=��l~,�^�2�.M-�3'[~�2�U���}%�}(C*R��5���9�dF���N����T0��㬔���V�~��8�H��m�I&���罭�XE"IO��1Lo[�Z��^6��s�!S�%{��C&p0�r���h	[11J�a	�	2j��4�k�&��9!��*�,xn�$.V߇p�qg����ր�}��un�T~���)���)R�9z��:{��hм��Az���@ǻB�� �ZHV?��G��)��^×��O�ή>f��b١�Z�$G��
��jq��0�cF,Ϧ����qz��ñc<gm�l��6�K�����	�3F�a��3�yKa�"c4��Fj�
pO���i|���,@��U��	��= ����<o������5J<>`�hh���jL��%l�W�l�T�s�hy͢�D���au~���v@*��){�Y��4��'������v/��A+����+�wÜ��tYe�ز8��J$[(�׈ ?��nr��`p�:�-�W�I�9W!6+U�1�̷M��v2ϟY��F�R�����ޔX8�L��9}H^5wr����ӟ��^�zh�)��bG�f�b��3:m���ə�N���k��5	qr�둀�� 鼛yg��8ӡ������,q�|�YcJ >�r_�a����R��gց��iU%#s�t��	�:8�CS9wl��H�D|����������3�L� ��������U.*�a�({�-�;�m0)�c�~�EBN������Y&�C*�b�}�rV���4�l���_��t��SÈ�%��i��%`Kv %�\�pď ���y�xH��s�_N°"�Χ۰g�S'��7W�pKCm�	U5#�#D@#��S�W��3l��Dk��\x�=$��~<��q��|J�MQs�����*�k�U���<೔��9���@�)�_���%���|��()�?
�kx
��-� vV:Q�lPMkU)R�yMz���L($!��Z��v�1a�{Y�=`m�Z�X X�F��x(ov�oDO���x�xaǷ��{A��ҥ=,�C��h�|rH��`���f�p�G���3�D+�z��M��g&$a�sc��X��[T��9�	�����Q�<�W~�5cϖͻ��웙g�N�&�����`�ئdy0L�H�B�2$�~ϕ��q���c�S1�%*�l$�߁���&�	������>�N�xu�	@�ș|[����<t9���>U8��n���zE:�&+R�{����<I�~�b�U�p`O��U��@Iz�LaVw5C����n�;���Pݿ��
�?�n��+LJ��o���j(�1P���DA�>0�΍�u=u�����R��9q��8\BE/�4Z�n�����:���n�:[\����=$M#f�|��b�b�<�h�1�um�I�`���4�Jc���W�\
H>��}��Ф��^�e)��N��d�)�K5�>`�?7���L8d�uɇ h�$m|C�C�4��8/���s@ж�9?���ga�*�� �4�ת�@�$�G��<��`�GU�����gP���0��K$X����g5,I*	�BԹIS@D�[������a�����oԠX@�ǀ_�t�k��Bt�� ��P�Fg���v�N��H�'��� goA[�n �$<a=��'^��H=��ҳ���Q���0��"��.���Lى		0I'>޹Y	O��A�{Rj���ώo,*�&�;��N�Pi�H���U�ďp��Z�ۥmY��u��"F�ѮtQ����v�;CBɡ ^��bKZ�-Gt��u�������2q'�Hպ�^n�o�˭�S#N��5xO��з�RgT�H���^��U���*�2�\yj�4���נ>�k���۫��%�UE�	#J8����;�M��nH�Vs�m��_�x�����h�T�Kd�n]D���+�u���Gi<�I�ԍq����X�O�%�ԋ�2P����m3j����v�U�}�\��H�j['�1�W( :�q��H/"��_���d�h�/�S�ŉ�D��z��-�M.c��}��B���χzfƼ�>�S�S�K��8���VU�q����i�8��L����`��V��k�{���a�0|��z���I�L�y!{��^��܈@��yi`t�$���о;I0M`�m�
���*׀oON\�B�f}k!f"�J�����K��"����7��9�l�:�� �w��F���x�~e�G��I�)i6�5r��,EPH���+�'!���0���@`x�z[��"����µ`Z'�4].ы��h.����͐���U�^2����=`S�t�@ȴ%�Tm�M�;8�y�w������H��tӐ��o�{ה�f�Ye]���乂���qk�{� ����T�L[�>�����Zƞ�v��ȿ9V��~�U3'���z-�Ȋ>��w� �l��&+kY�{��3f��'l%�u0�+A����88��r�Bo�!ّT,��@w��mX�y��x�����VY��f����	V0��pp=H����3n���	A�:+d�E�xD[���(�G6}E
%Ci�����zO�HI,��DX�h�]C���?T���Q]7՞��5� H/��9�����J����$���אIR-�����i�hob��O��#o�y1�-��G�L���#d�w.͏�r��1�J2	!C�V;X�q~\�vPf�ҳ��]P�N��P��T`k�U��5Ԍ�bN�AG.k���T��Q�V\|Krf�m���ꤒ�݋�e���A����~�5��C�3O��|榄P�X�¤~,%��auVL�	-*��r�8�ʮǓS��Uj�=�
����;��4/�{!�P<>*�,���ݲH
��Vv�k"�H����*h���uN�誵y�l&^y��I��X��v;~p�fo�t%��&��*dޭm��0�h��m�ccxܯ�US��[x�oh���y�Z`3%�q����� ��%2��8��dJ�<��樳;ʕ��7U��6�H}���R�i���C�v��q�[�%?2�t��G��K����o=&Q��Zn�"�>��R�ގ���7�� v�cp����<P�$�6|���/j����A%����`ȠJ*���P�7�Cq�<���	a��+x�U��鍹Z�������lh ;���E#�K�)��Vw}�5Xwk�-��笡�X0	�_P� y^��10P;*�d+�X9���Ń*?}G6����Ǡj<1}�.��J��n�}�OV��	��c�ջ�<H�"Sgt>���G�̺�h���R�"�B��.��@�m�)��CXm�Kʈf��`��eq=���)��pX^4�x�`)ΰjk��?�* ���x�D����O�6�Qʰ����_���ǈ�&
oj n��n�..	�
���/�KW��@r��;�/��Ëq�������qk)�JJ'�����[��5;��%?��#c& �1��!?L�;���! �*��sA���+�������s���P[��P���Q�n�y�Hju��]Ԗ#�Hf�gz+ޤy�|4A:�"��1zRB�ػ����Ҧ_.�x����ʂ�R��p��PExyl���C G{����/.4��gwe�|U�U����P^�dǢ+62��H༏.����tH�M���e7�?>͕·�H�a����p��lY|�t$Nh5/��R��	�+�0���Ba`������xdL������������(\6�|o[��%G���~��b��}�״����ס����l�����ݹ���XM��D̘}Q���U���cJ�	F��� :,ox�,mN^�ڪ�g���K<	'��#�9����-��+m��������?���-'F�.��<������f� >T�Q��p11W�3.F,���%^H#v��L�&?��r(,���k�2��D0�sH�F�w*O��N g=8��a�Vnq����n��
��j������r�c�L�����a�:��>?k�	\Go�O|-��� �o,�y�b#�8<8�q��否Os�}�S�2�XB|#�{7�o}���z�E�n�bW��(��LeV�V&梽��W2�Qt�A5��Pq��S�*�'����8�� �l�a1%���D�N�"�
�s?�������������sq�*��kW�tW���Q���'������{�+- ���
9qs�*ᛟ[�Ѫ�����Q >
z�Nb���*Qg{2g�|�`��@�Z��)�F%B}2�)6'�N֧X��GnuH �`&�(���p��{��7vD�W��H
�m,�������f|����V>�9]�խ��I��$�Bx9;僧՘�5�S�� ��?��كA�ˊ���dx>-	�<���X<8���g
E�5��sh�xފ>\!ْ�G�*No!چX��������Pp�zci�wr�6�r۝��2��)���(����\W�ݧ�+nCA�EC�b'^@��JˠC��!�,�ām�������7�e��RC�}E�<��򋦻f��m~��~����Q�1�Y�\8Q�"�$R�TIu��6�����mN ���@�H���qb��T���#@��}���`4��8y)h���B+S�D���,['�_}z��W�~��F��.��������n�"�
+�Lӳ3�Xxq�9Ncc�����A�����Gɰ�W���u&T�ǈ6ƽ�c{�,f���J����~];]Q��frCa�� |��
#J+��mf4/,*%T�Ìk�
�ނ���p[-W�D�u�����Gb��<j-F�G���	E�X���K-T�]�mA(��&m i96�{�"a��n���Ŗ�����&[pÒ]���|ɷ�&H.�H�l�]��3���%��X�s���dDu����5�|���M��36���aXI�
*���Y��U�:�4	�aK`�O�����z��9�g����z>M2�b�}����CN_����7)��9�gd3��d���v��zF� JQz�����W�&1���C�z�����cn�|����$a�#i�D�R�2�U���8h���_?b4�;��Y�D��t��AW)j�l/�.7�0��S荪�S.�}ߞP �`�+���W.;�)��ae�!w������π�ᾰ��,��V�(�f�M�	������!2�^v��1�%�S��忨���3�8��c��{K�w�W ��G�r�N39�6�ص٭#�0���T�5�g�������#��nG8���6�Q��Y�\g4�-!bH��Ro�)Q{Qt�H5Z�6�g{�Ru��}[�\
,~Lg)�%D�Ρ����j�E� -q�BY�Z7Yx�fP�*�O\;j	U�vy	.����[`dU��7@����P��՘� ��b��J��;�y��d�"��V�pq���ʵ秩�wMz����m6��EH�(�Eh����ߎ�4<͎�h	T)b����@�K/�h�7g�>��dtGR\����,���T�m�k<���6�n�M(��F��dN�\}�@�ڜ���Ky�k�@�&IWK�Q�e���dret_�^b	��K�V:���a!��!�ba�\�M���c��Y��	�|Md�����"����s@N�ܰt�.�a]M
H�}�~��?t��H�GX �ܔ�m�:��)D�,lR�S����ko���#Wg1���b��6�S���k�#
=m���"^��a�7~�j/�"sb��	kKP�.f;��i�F�(�}���U4�8��:��ɡ�a5Da� �O:1m�(�H-��Q�F�)�ˮ�o���ך�4��h�` �st�}�=46�⍟.�c��j�W�:����]���:�VB*������"����}���%��>9%�{��Z�E[r&r<O"[��W*Y�r�3+���C�I3��tN��ldTy��˱v3`���u�Z���Ɨ6gd�7�GT6� ����B�V�&Tң�*�r8QEF�IZE�F(����kw�r6קp>�jWŁ+>��N>��T7���#�n�x�d~���T8�⧦x�"�!߱����A�c<��Z&�#rFxE�~Q��4����z��n��(mg�*
<Z*b�y���������"���9FP��`IM�p��&y�,�I�Q�
i�A-��;[�,�CZbx��ϡ�6��,Nz^���ո�|s;��Z �}�QT:�i ���*��6\��7V��eN�DB�V��w�s�{k��D�k<\������s����7��~�ۛx�����F����]b��wI*iwD:l;�>%�7�3�nw՛J���h�֗N[J���ѻ�a�]I��o�"W�	�q(k⸍��!{�7Q	�	1����Õ}����D����! �蜃d�}�y�V�x��!5XY��YE
�ư����;'cb�y0�ڈ@bA�[�1#_V�XR�q�.�B%Qܷv"�����U4��
�(_��pڋ�'OI�7�$;��l�{����{F�(,��ϫ'��`��@�#1S]Rn2�wKe��^~,S���#�&>�Twm�9��k��a��d�&�mЍ#��ms�2��p)0E�W1��M�|�󪥎b�YDH����f�좰��
��JZ��Å ¢�H��m���Mp��6��_�x��?��p��d� ����d��htt9�?	m}��(�������!���6!6�yWD��ez�}��*g��렶�Q�N}%�_��m`E��- 42�D|PW��"��+�O/%;�E=�A����.�|�v��8  {!�g�[�v�!��ɜ{��9�7G�:��uޅ���o06� [�onb'HZ���Af��*�K�+� �s�p#�-�:���#�Y���?w@� ��X�:Q�����Z��f1w��7� a�鶰��[���'���,y_�(����wN�턎��f����A_�gfլ��Y|�@������"��jJO��c���rwE�R��U9q�*�x)V� ��_ni�ȷ���,fS)��
�^E��� ²7}������H�������H�j��"ڧ>�.��J��k~�f��ZE��\a7>�	wg���KBa� �+4,����o��]t�� ���b_�!�n<KF�\1��)$��a����MEk���]��Ԩ�?�#2fLg��!˱��#� [��c����ҋ;�x%a8S-��]aa�?���m �����ĵ bDu��:b)'z[?4j���d���ë�(�������
[���t�������$�[#�V�7�sI�P:���|k#��T@J�O����6�A^�"�	��%#:	s�Nӛ�l6˵U�rs�@ ��@����^ıj�=��� �+�Q-��{\<� q)w@�C�Da[�*D���J�:�T�؞Z &�ҍm������9(��U��9��8� �K1�f}t}�b&�JP@x�[�d�㴖�^�(:џL���]l��,(32�5��&���獨��f�@�;h崈;݈b�]�%\�0	}��@�\����ZE����N�}ۤ�H���,��#(�V��ٗ�"�#t2u�Nhc�Ύ���Y[�<��NKj����C`n]�W��5t�ЌC���Й��)�i�\v�;�ѓ���e���N����x�@�A��?�ʾC.���t�I͈�jw��KO�X'�������ڹХ�'|&YN��o�b3W~k����JC#`Z[���67v��^7�wRcƲ���R�\���(Yb��,}��:����n�N�D��Н���!�"Jm�����F��p���[� ��/q�p���LJچ�uw}��3��I�km��KpFz�	l��x�\�d�CP3�z��J�� F�I��-]�r#z59��DHz,3��<~�0۩�;㗎�ZRn���ʋ��P�t�s�|8�l����/r�b�,{�
�o`���ʖ��y�W�M�7uP�\�KJb|����-�|�s·Ta��~��w�<0�O굴`����v�V`ۆ;?I��qlZ�<��8<�)N�Fl�R��_�O�M\^�َk���7#��X������=���h�V�/�]�U텄���f�b��c���",G���V���
m��?��C8�*sֻ��O��SU s>���(֜�T�|�h�{������V��4��.�p��b��72���������2]�˛>ȅ�͎���~BB�9Eq�a�d�blH0r�:k9K����Sc��ƴ��j=��lh��;u�����^P�Y��.M侑T�B�O+uD�P�Ll)�T�xF=����s`ED%�u��1�R_a��n�+�c$�>�){P�b���5��S��;�IWQ���S�wZ���z.�*����ԍ|T�j�>z{��Nv1��$�%�e�l%��@@dP���'xĊ^ڶ���28�2*��i�d���!���ě �l�YT��>�q®��sS��%p�8����b�$
�pI�Yp��b�S�`̘�x�
��v��z=��1I��Q��&�nP�[��� �#I8_�&���&6���Ǐ�:���?��ǾX�GN���%ӵ�i�6��j��r���(낅ȥ��K���;�8Gr[
f���_��Fn�n=&}��2�`�Id��]��
\���1��\�V�t*���r�JCa|਄G�8.�\�6�^@���VS9,D�pA|$R0�i6�{�;��� �3߉t{ɧ�7��!;�?�hpp�g}��n'�j6���B�@n�U/~"��ڨ:�-�Y*�/�� ��16���-J����^Qf�;�V;��8ŢfHBt�v��`lcl���sT3_��Z0U�g��n���m��VdQx�L��*�ʃ�6"�0��Q�y�Ш��sWBC.���J:���w��$���=R�P�Ņ���"c9�E6�<�e��s,~M����<L�H�r��оwۿ�&�	tT�?4<��gQ�u=_�Y��۶�]��0�ݽ8���G�#�j&��g�ʃ!��]cy�~���s
����e����I��s]��M�)gO�`�@��<�V�Iq �6���LQQ��C��7I�6Ԓ��E�Ez��!m.|�dr� �$2��Gy��!�6?W�@C��H�X���lߟ�W��:{9�@l�(w����O�_����گ�r�)���[��p�?p$�=`/����H��z1�?�ݎ�ұ��ۘ��t9)�C�k� �����¢���d��K��8[��=�\���@!Ǜ��'�^���ݜ���M��VRsv��S�m>��;��[mz�����h7{���5�0a�;O�꜍;���rl����5��gV ��}J�����&�DLO�޿3���$u(�^j�:��6ѣ-��ti�6�:�l��!3�+���B��ԛ?���sgԎ8��P�EO�O����[l�[�a�K=����i�)g����ĄL�f9fQ=�}��HIl����N�ӓ�:���{3޾�wW�ZN�9�#*��\�����`�r]�C�U�@�d���8C���P�?���V�����+���u��teHC.ғ��VN��~Q�Ps_�nE�lcP��M�0!��o����p��]�Q#=X�����"Z��޾��?U�*�[����g[��Ө���j|��P|�7�^�U�����!�j��e ���R��f�Z���eL���OK(a3���[�������CQM�G�~��>f�7�@�h��$�d��ޞ��^��LeQ�6R����^I�EB;���%+i�
�q�lS�^v>�
�t*޵�b����1�kB�KD-}�@�(z��K������G�'��{EC�0�ůR�V�&x��^o��.���;��8��R��՚����MK�,D|�լLh-|c(����d������]`�?L��<?��)`F)��@��e��w?N;ϱ�Vgp =p�rб�����	D�G��V������&�x)1*��R��y+1i�%y��)[�D �b�װt^«��\�ÎL�JC�r�]���,�G����E�a���Z'.���җd����s]i����!�J�}�Fv+��5*�ʗ�V���/j|h\$� �4.��v^����?F!���sW��_v�:k�H����t�{����q:�h�����a�����|����e	)�a�j�D�O�����|�q�R� L�gh$Zr�q�2odXP�γ�^L��ȁ@pYM<�?q{���a����޷����h�FA�O����"5sB��;5�~K����:�~q��q�Y��/BV�m���c$�����]���/��t�o"��U��{�����ה��ƍ�X�{}:�D�/�dc`��������=0o�Gk���;KS-a��J�0r�)-z�>, ��n�/��[�Z�.sE�EHld�R}q�>��-�$�,��|[�_�+@\�G���\�}��NdA�V��`��Y�#e��hG!���:������P�5�s�pC3�a�� ����%�o��&��c>��9uRN�.l�M��V��Plɐ����A��W�H�]��0������u��Ƀ�_3I�*���-�n�xZ��zߖ�ޮ�h�dǁ�,ʝx�i<��yyq��'�K�R,oԛ%ܞ��_�yc<�S��c�֘�G����q�Cd�!���ش;I{�Ŵ�
0)�|b���P췼g���E^���J�ecH˷8�.����s`�ө��m����}G�A+.��B3��<�%s����\U#H�Cm�1��=�Vt�X�ķ�4^��d���|̗��R��O7��-�䉓c긃W�	�c#lc�7^E����PD� ��kj��R0�}C�@��6�\=�}��s4���:6ѣ���'&I�o��A�(s��}5_�Lj-��݂�,�����3f4���>�L�A\���!c�;f�	���$z�T�(I"`isx�7J�3�L����D}:j��x6F�icWS���?������Wq�]=����|����[�;�y���	�.�})!��D�GC���mEk��>s,ԟ/=|>�b.>f���m�ӽ¦���+ue��!T��x{��T&�Q��>�7�0�(P>'�Т�����@�3-�2w햴0����� o��T��{�����<yy�$��!%�_���@hPr��+��H?������xk=�/C���k���L�?&b��L�A��Tr��Od��;]�j<�D�Y�L'ƻ?�]���o'�������Cy�2}��~V�{�L�<x8�z�U`��<F�%w+u����yrh�E}���|Ƀ-��I\Kc�����!O��h�76pn
͒�4�7�D=p��!%�.����_2vl���A#4�e�h���*�M�� ��	�4<�ȵ�z*j������V�џ�m�L/���� Oq�T��"��ZW�
e{p@���v�ⳙ�����Ǣ������*���q���ҽ��P�墺��sju���G����4d�<@�W�U(c�&��E��7�6]����	b�8��مA��9ʈ��ֆ�G �^l�o=8uI�`s��4��H>I]�=K-e��_bŪ�}�4ҷ�)^+��x=���a���Ϗ���Lė�K���Ή*�ٶ/'73OOCX�ۙ���ǻ$AQ���J��O���d\Q/H��ܴ��L���̝�"m@t���]�q^,�q��78{�!w�p�BZ����?�˟���!{�2,�tV }kj��Q�]��r~�y:$z��7$2�,�:K`]�ﾛ2i��O8�XԽT�!�&�=�~��J߷�t�T�i���)�z���,��FdG|��O�rl5��2�Ww�M�~oY�u���
u[��,��?��k�&<}Z�o<����tHRv����8�� K��V�6�2pB1�rd��-��������,��[�ڴ<�N�k ҞRI�.��C`�`f	hY*�X��5p{�Q��D�p���nsT�}�&��-Xgr�FP�A���º�b���>/�J���w�0S�/�,v u�) �s���s�6 �i������-Q�H7�ҳO������p��Mk��S�+��{�idWf-������U?5`�p�-���� �/��<)��m�<-WJ��T����bpD��ߐ��څk�f��	`�x'&ǋ�׎Z�7ק�FD���f�����g��8)���b����Q�D�&�rHA���Nu2(�ʜ���w�#�Y�A�X����0��q-�p^���d�ħJ0f��gK�j�l�^ܾ�
	!-�Fm�~�^311x`��y�'I/j)�wcp�ȸC�N�_�R�b��ɏ��^ؒ����p^-����%�����m%�]a�~n�y�L%�6�a�a��M�Mz��R٣�\��� ��bF�Ƣ�PD�M��4O"?���
�6��k�u��x�*]�R(K�TO���:H92�-Y��oʁB0zGJ���d58��5�[õhO?�Ю_Ľ	k���l+�`��~z�	��{*��1<ʆ|���#5�Q�V��7�>�W���^v�kۼ
y����扥�M!�,)4�Ċ	��6�L�R��C��;�Ŋ
n��4��|�V��S-!s^�����tVLg�L}͵�Sg �Y�݃9jO��ù)͖��?d�K['�JaQ�>�/}����a���X�˂'���Q�w��4��-�ÇN��<�.�k�����ܝ;��4�RYn�ǉ��P��q�����1$���l�
Lʍ�c��~�e3$�X]�E?��G["�.����e��V��ԫ�wiN�'�Ď;��С/_��B٠n�)�����h1���xM���O�s��`oL��4�T��
���)(����������U��Tj@��n��>P�����4��Ҏka�ǵMs4��A\[��i��K��F�Zl	x>�ⴉ����_쁩.��{5Z�>w���~�s�[����K=o�p�v�֭}V����l��k��V�����9m��jI�5^��*�W8m\H�}��+���%���H]T
����~u�H��8;H��M5D��-�YcY��8h�olx�I�hW\���B4�Z�آ,z��.X�)��HSWs�3)��PY���a�?��fF�ܬ��.?Pb�[��R�����$xk�}kZ�� ����lnr��M6A��Y@�/t�_괞XZ`�q6.��F(��j�'z�G���8�t��Rs��{�e�1$X�S���|�vq�~y	����+�`�����!h �=���©�d�:��G�K��_G!F�(v���C�zB�v�`�,}<Lr�&A������ ���?���(��w��� X�OI+*z7��K�BQ�F8'ɪt>���v��>\�Ǐ�m���Z���\���͝ t�%�i����P��̡�o��T�D�W5���u	��ثFUn������Q1�Fu�
�ڀ�����܂��."W�әM:�Y<S�VC'X3s�a�00�=];�!M��)r(�ަ]0��X����#>�e����͏΃*��v�W�#<r���� �d�|�dS�Q�����σ/�aM[��K�A�^��(�����_��M/S�$R�/,�s��Ə�t/��M�����`�n0�Uřl{�S�_,�%��Ip@0 ���?q[L �r�V��z�<kik*����Y��tj�����cD� >��N�D�æd��X��vؽ<V0{k��,�ѹ���T`��f�L뀳|���<��|�Z�įn+!L���QX�Ħ߄W��xReQ�{�LvR�������5�0�k�u ���R�#��#�Ê��i�|Eΐ8�XO�}���P	���R�p#:S��8W��O؃M�DEP�
$�t��g�U�0���	��:E��)���Ho}���1�N����w��װo��	?Na͆���%K�[I/Ov�
���T;��S'<�XW,�
<��j�+MĴI;��X��C��1�z?O���q�߬*x�R�x�m����R�)SiƄ�D���괙�bg��a��Q��0��Ԫ��>�#n��x���0Y20��W�[�I�/%���^`#ϯ�a� �XIR�q�=��v�8r7:��H�X3�$�֋u���d����VA"-(H�#�[�J31���L`ߜ�j���w${[���zfz2-��97�Z�$1�S�ɞ�V"G��Y�\��6(�U�_�I)��4D�s�%�,ql\�ݢ�>�>σ2݀Մ�j]9�팏��q���!H�j�7��)�Y��n�\ �ŭu��пܟ��e���>5~&�&9n?T�Eg4�-!�y<����hF<�=�E���9��(l\�(�#�S�_.+0��z/�6*���O��Լ]���m����ŧ�0՚�������j���y�c$�a^�֯�h�1�D5�7	o
!�m1�^�����;0�3�U�,bB��>������!��۶��<[�ᤉ����,)�Wj�����b�	�tBp�c��F�%�����ۜ�_�
q?L��W�2�mxǭ�E_�6�#�q��pÃ����M�r�k��6��3e���e�%A�!�W�l��U�޴$���;�X\i��5���V�f�^-����m<ި����i�j]#fY���`e��)�� #d���ϕ�Py�tצ/B������o�%�dz��
g�%�H��}�R��CQ�1K_`�pƆ��ۤE���U��K��M�Q�'�&�������$s5a�4D�����e���h�|K��з
�ZJ����q�	;����C���Zh�W�wڹl��f���A	�\s8�\s���%r��0�G��-b?��`����L�i��sBL�&�z���f�ŧ���wңh�?S�s�i��t�T�FN�&V���"R������_K�*�g��b����y�2x�!�C�RZ��B
�9������	}A�FV�������!�z�P�R͑����_���Yh�^4��#���Ys �u(�I�1�*P�`�7/��f�Tl���L^E�o��,a�h�!B\���[�
���d��H��@FQY�"�~ie.����HHZŌ="�G*bX���k�H7῵lHI� m��Sa��+��QG��\>�G&��'fz�<MW	��0�TP���q�.��6�T����#�%CS�XV�f��h������/l���$=����%�M���[&�2V�gr^\�?U����/��!�>�繳R#^*� lh<�1�j���[�o)藐��ЏNIH��0M@{#@<��ɺ���t��ֿÛ�!���7��E�精�]�Pe[�T��Mwؙ,��7&;��k�>�+���QN���a�4��nR��:w\'>#7�W�U4�u�(�5v��� ��d��=z�x�	�'�^g��%pY'*2��>�=7�_�H��i*�0�8��
;�����NTx�)h9�x����<�bD�0����oi���5���,��h ����T`�\�!��e�A����V��ռr��f��=/��8�����&Z�4�\I�U!�
Z��>j��>������\�#�{�C
�Yj�i��ւ덎���Rt/
,\D�=K��}Φ)�0���� �n��R%0�ʌq���r,C�!����s��/K$���̤^�Xh�)�t{�"���5��z��%Gg�q^;UR���f��-�¥ۛh#=
�RWr����wc��$�ܪ��!9Q��^�|0���s�ˬi��)�IF|�Q�U�rK%�7fjY�M�Ę�m������c�1���x���`�����8����2v���?��t��@�K�����p���O6R�6��~G�d�����Ӳ���e�Z^^jP�V�Q�Fuі$�vn$�G�bH��|������L�N�j���ӗ00	A��P����~�L��CN:�T=���	td��7��,X Д_�p��Qŝ@�k����T����e��j��aYO�� ���T2lV��I�]z����%�I�Ԍ�ݲ�J͐����[�R>�?B��@���e��G#p��F��5���Z����I%�Ǉ���|�l��2�*��J8"a$KJ�>* 4����{�􄩪�d=Š���Ȇ�0�%NoM'\��f�
5��웞��z
ԗ�ˈ��HLM��`��!&��Y=Y��ISE��E�I������Y�&.^�Cm���)dxRc�K|oD5W(nh��������y+ &'1�93�q�:'�F15��e3������)��t4� ��r�Bߺ����������"���13�+:i����9�Ptb����:�"��u�����nv�� ~��X|b��i��&�´��fN)�{=����h��2�_�=W�3JhMҦ����ؽ��s�fA�el��r\3�c[�0)A����@͝ �xmFF�أYBWĎ� �y��Z#�3��P�,\�#��� �qD[�lх�F4�M|����`T`�-�'Gɜ�|��<�f�|X���uS'H�,�1׺X 2w�-"�a�O(AY���M헜\�_=zݝˑ���q��s�0�ǔT�r���2�C	��e3������/1}�n�~�J���������&�+<����_�y����Rz��j���?`	�J��В��`I>�ٹl�"D�����c^�	�x�teؙ9��}��`�;�X��o��������DF������'�)9��L�!&/�����\�~��/�\�v��H	�,,�pn��^�Xө
Q�aO~#e^�L�A����Y��[���=W��ILx��ttF�t:��K+Q �ۿ�L�hE�Q�;����7��!O�k��P�ٷt��!X�5�Hb�ƺ�u1���ʥj���,,�/���G�f�S(}���c�����P8}2>��F6h"H�%����
��sMz�䤹���@��]�ӕ@4�`L�(@?�h��:�?�&�T}'=��8l��#��$A'�wW ��$��)<��AM�ȉ�@(��ݕKb�z/s����d>3
}�� ��S{t�w7T_#��f��ћ[��x	�����&���E���QЙ�$͟%g�w�0��n!l��������>���8�	�0�� ��\���s_g�Q�8�a���4��=Tq�+��x��L{3�Z-�\���Rx�VP��rR�מ0���t!�(�3q�����HFY�AN�-����^�4퇃RTq����ng}���d9�Zҩ�g��[�c(غ���裏�a�(�ֱ$�FP<Vq]��au�����@���G}���3�ث�2�z�%���A?�#�Ln&6�`�Зo&����IR{�L��5V 
%���_U8^����"��B��B��0_�`\���}�I���dv��s��  C�v �m��\���E�#F���EC�id�z?�����:��/��&,�%�ʳ��~:XI:�`��H���s�α�rg�!�f�de��i��\�0V_�>�},�b�ʜ�Yԃ�"C���t���2V>���K��WI/�y�t�M��<�i��������k�W�U�����v���䤐�r�ދ�c���UP���YGM��8����Qam^�Q���:X�80�<�Q����g�,9�����Oĵ�ȜKn4�E�g��˷�/�Ĳ;�.\X�V��S�8��^}6�
��(W.˚1��rE<����K�/�������mt�g�:��5�q�uG/��c��j�֬��K?
��[��M��Tr����*~@��q!_̯��������?� �O�.RY�"��L�o4L+��HWe��3��1�i�'H�5Ϙ��^�4�1d���P�5>�4�]��9��1P�&P��k���H�vi�O��@Xߞ
[tҗ�N"��%orM��%�'_�v�1�;b�N�����1�0k5��*W9Be�|�hl$Y��;��x%�a
�c�� ���ڱ&a��L��S;y�X�J_4��E$�F6�����c�ţӐ�p�����Ȩ�؅�lab�2�7sM窈Χ�pL�1{��4�{_�A��韎�9(�.��]R
�Z;�ţ��v_k ��]f���ȜG��ҭ�@Wtڄ`Q7&�����-����k�N��D�%��y	����$�,�忢J>��79��'A���_?�xjy����3p��E<�I�$��Jȫ����0��jtAcc�THH�_��F�y��
�Ei�����"���Z��𵗬!�P�K9���S9��矁>��A�w��E@�j��|C�G����C��$Ds}W���M�R�m�Ӂ��y?S�&�=�Σ�9��n'�1=���j'd�i�"GL��U��>��53��6k��63��us�zZʫ������9�Ҫ�8彣!�(#W�zY�kGQ�;6�O��.zX�f��6�HC��fM#o��[P��}���?�n`��TZ��,�|״�1���&b�Ԇ~ѩ��֢=���kv2-y�,[�լ�t玹m�s�/∆�x�s.b�fyƣ�4PV��g�E¸�
E���E�f?��Fџu��o�*	�6cn��^�&��$;��utv���0�L��lŚ�3�x�"�0�vZ�h+���1I��T�����r��(j�'eJ�9�۞$�֣�.�v�RUɮrW!�9)�B���)�}�^����]�S�տu�rt#��g��ԛE%S~&O�W��[��:)��ʺyò[��o���ʸ�X'��a��:����bV�T��l�Yo**��]�����[��χ�;ٕٞt]�C~y*�����φ��TTD���F�s"��4��_�@��]�<8������O8�o�t�8�n�>��G"4�1��8��p��F�E�+�u^�'����Lds�M���q��謏U�A�X�*��?*����qg
3�y�5S�ׄx4ct����>��[�j��a�ƸpAx#��9�v� �����a0�A~^(g?5�F���)��Qm$r�G��&Ѹ�s"�ӮU�ȅJ�t ���G��/ԕ������P�����f�B�.�2�ذd&�� �݄�n��dm	�;HY��ӧXW��OQB'�:6�V��W��
����B�ٍ�[g�xjDK��w���n�9o�B��W�9�)C�)�>��ݫT
�}hb|*n<"�q�F,"�f����c[���D���]j����+�����"8	!����OX��GU�n�����c��8�p�.���%�}c��
�y�Nߝ����ZaY�'K�JP�C/�P�eB{$դX�ǽU�9n8/ա��v@Z3��fecͲ�������Z)�Z^V)���n�yN� �]���th[��%��T�����A&�F�Y��*	WZ;�E�.�U�%�
��Ѕ��0�Ό�[��qR��_�3�WE8[/ǚ�&�����eN���L���kOC�u|�(1�q~�B,@��?��[�;�E����Ow�!���Tn��Q��հ�IE,Қ�z*�BEsAdQ�G$��������ˌm����?d�t����5���f���{���4��"���2�ȓ���Q�Mg&+���G�3�-ae��k�Ƃ����{�V��<	���"h��6yn`oZv�?�Dg[��Px7�7��k�Q�=1�5ᦿ���.^�2����^ޢڗ	��l���D'G����s1p��H� ��.h_%�dM���m@�Auq�s:�kKy���A34��}}1��p����Ꚏ���T�6TW"Π���4���;�n�z���;����������A3���S7�7���Z'&~2��{+l7(VJ˓-[aH�+m@�B�5Υ�gȬ���-!7�N�)L��|��cR�����¢d����Ƕ�x��KI/�~�2C��D�ڝc�����`e��� �N1ǀ��^L����11�9�kj4)	T�^�=�o}���a%+�o�~�h-i��dV�ބJZ�����I-{?��_m�S��^M�Z3�
{H,}O�AG�#Cq��.����ć��qPn�t=�x0��Q8�����\ژc�;�YXX���R<�
};.2>�9�U���5��o��8sc���d�°���V��ů���i�{�(zcH�>G4��ĝ�ǉ�I�@@��=��*�C��oS�?�����3�(:�������k���#-���J�>tB�X����A2k���b�J��ԇ�ɴ��(X�9�5]CS�*���SN$���2���Wk_�{j��n'���57�U���gt/&�
{  ��U.n�IY�ErD�ؽ�7�.��X(�ܩ�(���5yN��y	�@Z/���|Z�ֲf'�E�ݚ
��}kˊ8�M�E.��Q�1SJ��ZT���V�m�W�~X��@Ɣ��!̥�ȳ�g��c��H����~�$�}儧�d�DZY��4�w��;Q���Z�0,���<?��)K�� �s�Όۥ�4I#���o�y�D�%	�>T�&��Y-h@�t^ef���'\�bZ�����`�'����D���H���CC�ʳ�;2l��'��1>��rn ��������C�J�qV��F
��
}F��"�K��`_@:&xs�-O�� l*�R��hΉk����S�3=�}	S޸�ܠ��
�mj�\Y�Î���s���O�ŝvb� ��s����1*����3˝�
�,$С� �1�ژ��þ�t�t<>eY�=��d�>Ċ� 0�G��b�0�	��Ms���&�0�
͇��w�r-���X1�S1r��Ohֽ���`���(6Q�b��u����>C��#
׿M����˥�>$���� p��n�K��w2p_o�b�?�}�6�zj�*�ݖ�o'�;�qC�*t���tͪS(Bi��ɴ�h����i�t'N��r�v~����-��넽���v��N�N6'0X����x��~�!k�/�s���4���r�q�\N��4Ԏ&E)��7�JW@r?^��a�g�i͋�O�Юh��t� ������B�\�b��(��:(�|�֧�+U����X���,J0b��lyz)5!��5�ev���˃�,uM7��	:��Y�+��߽Va|���h0�Ƹg)���"G�&�����C�ƹ8%�w�
�����<��N;z��먱��G� <�![�jt8�ʈ8$d)�׀Ϩi�o�?����:��;�!��R �y�^��&X3l�j�Q݅�J���t׭ �l%�{a(��N��L16�V3��V��b��?V�h�N��x���T9A��E�ѤE:ە9�
c������s�݊�qkN�����o�Q����Nc\S��f��!�*`��A4���W��a��[1��Q|���E�<myen�b4������dÉ���!{ף�g~��SJ^C�TdU�-zd�v-�䅔�%^�/��0��#�>��O+9Rj���X�Ӥ̾��)����"q,�Ct���@��F9g��$08Jh�h��v��8�����5Wv\���>/)�L����b����k���N�K�{\��FpC�6eկ��y7{��y&�W�r����`9>�>{��wK�X�B���%�_��$�,R�@p>6��ɥu�͜R��:�gT����!� ����/^;��D�$��5��}n�5�I�!�CZ��'�r���c�VO�C�b��؆�hrT��c�FF͇���!�qѳi\���?7]�t��q����3��-M! ":�/3m@�8��5�U�I�\�7���t�$)4��{�X4tַ�p��Io���|�~gg�1|�A�1\4i53�KS�~�!_����S�����G)��c��%F�L�J�X#��З������#���i3�i�/dϊ*���d�R�H�"[��-��HΠ�'$��A��!g/��=�nx�LK5-�JkE���+���

�
�����i�X����FB� g@����:3�9H��P��R�6idF���Q�oh|��R��(�[I�gڂ<���T�����Sp�b��@{�@��Rl���򁹺�z��K����B�.B�I �	�NRO&N~\�ˡ2�����Xئ��;O��")�'C��L�u#>���K���tY=���ϝ���s�`��;�>luӏ�2�ŉ Ͼq������`yKc^�� &m�߫�Q��\�#N'X�'2}��E��
�"a��fj:*��^���{f�E|s� ]�2����v�Sc��!� `����pU��5<�R�ئ$F�ŗ��!N�}��>�}q�H�*��8Hx����Z"BL�F"y/��cg̶�C|Ҕ[�6���w����Qˇ�Yr�n���xKP����U�UU.��ɜ.,���2���"��r����T�co᢯&����6㕂&���90�$G��:��ht�"���^�����g����6�	�Zr����79����A�$`i粋g���n`����roD�/?�Q���`���6N���ݹs�99Y�sΒ0z�=קtaqh�`�,�I`������$��i������0�_��?6f�,����g����lD�q���#*���"�/���P��ҳP�����8ef��,谶兦�i�;�}����A7�� �����Rf��^:Z��Y�Du8V[�ϯ�E��& �G��fp܏���u�؀�Q��~(���y�����
ly����5^ @�-�3�<�w�ʺ�M!��]���q�)~R)��Bwc6ʱ�˷�,#�A������K����M��y�w2��*�I*�%Ɂ����ع
��=6n\��a����k%����e�t���EH+D>�^T0�f�ȞH�M���rӜ������(J)���w��%�H�v��D���\� �S���s"]cs�ɭw;)�A�4�%`;W�m�~q:]ֲ�AU�V����!�X���o�������S0ԟMٽj�k_'o�_�fw��+;Y/l6�Z����6�k��H(��a���D�^a�5M{X�<>�a:t��E�2~흌�Ȍ��ǑdM�uq)�wG#"�O�Ӛ?R+�����,��u�G���/�@�h?��f���-﮶���q��Iu�a�y�֍ISg��ʹd���%b)��|�U_����� Qx�i>��N�#�$0�btiLqԃ{ k�]Y���;��X}�c�/�l��eG�C�tգ?�2K®[y&zZg#����z�
���VUh�y�La���D&�$���f�(�U.���������(y�Q�Ѭ]m�����(}+F�����FX;^4��Ӹ��>�L�\5�f:�Up��D\�41�0! �O�L�ȚT7��r-c��@� ��£ݧ`��Dk���p� ��v=�D�ˡ�̡��,y�DN!ݸ��T��A��꿧s����ez_P�ճ��/O��Pq&7"Dg��"_~������Ks�mY��	�xFԳO���T�Ou��|�}�k��;ù�6�
e3o�D��e��5�8���0FG�9N��&��>�u��ۼX3���Ƕ�Q��D����4[I;<e�_Z���V�z��`x�V�M�DFkU2�������TCt�P���ٿV����F`�ƝJ�R~�Z�3X��<Р2�m�O>(�>65zK�#2e�TMq˪�5� �+ %�m��!�Xu<�A(�U�gN4W�<�y������K��m�l(a�� ��(c��j�f����C��e�}r�ӣ^-J�g�p�bx��6)�/&<�. S���XB�V�$kx�ޥ;M��9�y���%��/J��m��J���A�fE K���I�ؓM���� -b'3�2��t,��[$y������Q�XvmB�g�5I܏Ԡ�~����+�lk����2z)��5���o�h��Ŭ��;�,3~T���o�p�gwz�P]�M��u�_vX|�����Yit���H52�{��,"���u���!��'"8Q�G�����b&_�YA�,R�����y:�P�:�)�f&B���gA�?��p�t�[z�~���@c#�'��||`"�Q�^,�%Z)�"�H%�9�g����@��N-�<�5�X{�R���:�~W��Pw=��VU�}��p1N��[V��N�$	�c�j��s��N NWP�yt���8I�UqMN�[C����3�b�&�"a��$g'��B"vI�1nB���5 5ĪB�Q��V�>���C9�~0)�	�2`���c+��ߩ|ۅQ�BZ���������1�֢(Ԛ!�d^n�~n��643�,� �ov�C0�+�(2�� v� c�H�i�-�� ����%��	�+��Q��8���6�N��3����F��5Y��ٹR��p��͉� V��|�>]�W�O��8eS�8�Uz~�c�wQ�o�9�)�$m׽|�xR�$qR�����'�Q/n�d% W(O�İ�~��X�b`y����X�Wx����5����G��$񈃩�1!�L�8�R>1\}N/��M@n95R�~�p~���S�H������-c���JTlC��.o�+��&��m�b��$X\t�M�4h!I;l8cb�$��3���T�^}9�V5��uj,:_ʆ�4���q�k��������K�d)ԋ��b�n�d�([X�щ���>'��'�,����	KP~�L>���e��Xt��"8����7���<#�.�R����M�=��G֋�߷q؍����8g1��T���v��µ���T.2y#E֨E�1,Q'y��<Zv�w]�����x� }����j�(������8G��z�פ�u�d12�9?Sƫ'��F�c�vyb��A���+���Iͮ���H$PX:��O�-7�+��4����M�Ϲ\�Cb�wЫ�H��r����0����,M��;��4=�X�L��O<9�";���13��Fq�%�4����fD�X����N��-��S�����ծ�����t�rC��_?�q��>��˘�����A����엽��;zC�)�(�xoGq�jZ�^�b�C����`��fK�t�2mT�b���5z��OS2�����Nq�*d�x5G�`c_���;R��T���{܎��:��Ir�ٴ��ਸ਼U��7s�7�P���w��x�cq��̲�uQo�W��?8T�%�u�F��ET%�˕�<ga`�����,M}�0d��V	:UW"��"�S��{���t%��)��C�^":��-�;�'�r�~��)K��;CG}?M�NN��H1e���I#�0`ֵ*���\J���=�G)6����O>��Z�׮��84�|S=�q+��:���l0���C��B������,r��!�u�{m�D~c��Z&oG`�鲼]kp+%a)�j���"#i��E�r��I�(�$��©v�|�'�oٵ�Ԉ�,����Y�����܁�����~�VL�E#�"��cգ�?a�j�b΍/u��Ŧ�����W�siI�P��Ec����*GQ�v1絬�}�t[`ޑM�hp�!�$�ɯ�H�t���k�Ƹ��1;X����t.�]�ɾ��z�û�¥����z����h�\����j�K���](��-�]��Q��8r̪R��x���f���N�9-fpM7#@7�d�Ϗ���!;r��oa7������k�!�&F�0���Oo*�V�>]�V	7=��u?7��V���f.6�B�>�|T�}Y<�}��ʣ]#�@&g��f�_��!"�51�{��5*�:�	-��d4����������m`��㾃v�r�S�1�����iB4��H�i��_�U�lA&�#��g����9T����>�G;e:�c�\�)�K1��f̓��S}��vW!
����1�ݵ^�iew�����T���y͛K���rms�!�~���4�M�'�sMf�
��5a�W��8�R3��}H��D�1���A�9$���T��(�擎a�3�1\�۶�ԏ^2��ٛ��#/c���C��N�=(_���!<>���u�_��hT�t��!S�����M7�܍yV2<!1��WO��F�U����!�@�|?*�K-[*^��p�ީd>���9���QȟV(,��}5lm���י|��p0���*���D_�v�Ѷ��H�]/����a}��guT6��2�*'�h�/ˇ�J�PZ�3�$��������b.ۆ�	��0޳;Oճ
KQ,��u��i���:'�CpsH,Щ-�qy�����c�VFtTٍ�(}��O�W��
ܒ��bm��ޞ�d~�4��e��x��l���[��Q�SM��u�c�u�kQ�<��r���jnͷFA2�X�#B�k��i(S��DB��)�<u
�?-|��צ���	q$�)���u6����%"�%^k�
��O5.�LG8k�=�)"Z�% Y�/�]����	�Ԩ1����i����M>r����)F��������9�ڲ��	��r�I� ݍ��{�E�簌�;G�,+�i���I1&��Y��Y�ҩ��L���W�@��T��w��Ktf�%vf����ѵ~��/��Ǌ2տo�D�N)/	�G}�U��zs�~��	��v41�6b?:��>[�������6�m2�Vg0/���#B�Mq]����v��8���	���Y�޹%&����j~ztr�����[�Dyثψ}CR ���#"�G�=@{�G�Y��O�i.��'t?�ŏ�+�������HR?�,�P��Pp�i�:�I[�TGm_X,����<L�!�{IT�SqN�ј斟��>����I[}Կ=6s+46jD�k�C|&�S<�򶇩_I-��E��l��\�Y��/�C�k/��qB�m���d�t��	F�c�)����ݩ��#�(�LY�$,5�U��π��]����p�س2���W�>9�
o+�D%,J�9� _S)�?)iI���è_�/��1�叶���U:��n`v3���)�R��
E�~pn�"#>@�D�����׵a�I���dl��M����$E��[��k��͚�HD�H�<O�ϱ��}6��Y>�A��/؄����v�̖6h�^b���@{���;�ы������:eb��R��P�c;��F	߀���X��-N��i
�2|q�ʬ�������6��9�I#2�g��]h��|�BZ�^fe�l;�c�6wܷ�g�Nx�7�?#OX ib�h�b6�t���"b	n�gZF+{�R`9"��p��q��*��(v`����;Ζ8P��9��c,qZ�{xc.��b89�,{�p�C�"��y�����z�Qd:g�!�����IE�+Y�A*sR^4����{o�����xW�r�����71S!�j�h�c�tB�V�~�7Ty
&f���_z�rd���������C'e(��5Z���T��|� ߢ��bdQ%z��+�Y���m4 ��
�K�(��7�iZs��s"���؞�8d!A@�(X������mk1�����:咗��h�|*��3%[1�c�<�vC�w�zi`��
7�:M}�@�mP��k��/ؿ���� ��1����@�u���8+):�.��9w�C����#!���{a�����Hz̎��;��|�Լq K q5�֜ �ӢvzfX�r�=�z�ơ�:��;���oH�S&��!%-|8�u0�UG���Y�(������FwF�)�������T;�}�ݿ=�Xa�#f��tZ�y����6zI$2
���� E T������D�ͭ MK	�?��^����Pq���ȅ�%���=uwu�k���ͧ���F
K(�v5VVb�+y����hC��K�����G����7�lj�;I��	Ԋ��� K?��f�$��m�LKq�3�D�3p�1��Ϊw��׌NJ�Cq���.E�辎��#�>�u�_*�eRAP�k��Oᯞ�p����ey/����(:�Nyu[�t�4��%��' >p��c�q��O%���W�o������	�HG~k�uzy�VRٴ��)�R�ʗ��q��ʐ��tgJ[�OZ俁�ᖻUUβ(ҥ�A�+(�szXn��i���/���L��FP[�V7����8@T�R�SC�������;T�5%��X��&�L �^�/#�q)�-�C�|���w�QB>\b^�$�D_"����}�(�®�7��b6� @ҙ�1��e�σ� L�៮���0J�q*u��/Ա��l���d���ў�cS�
�Z4��okp1!1^����err^��m��/N����M���V��A�Q`�g\���e�Z���g�"�&[�v
���E)�^;�P��Z�7mO䇟(�J]��)_�b�sgU:˾߫�^��^�{����#���3m�lr�r�\����OSIt��0,�6�5m��Q�C9*RB^p���`f��*ۈ��t�8�cV~���[.l��mTq���|��Ɠ����:��G�_nuS�V���d����O
�H�m&1��U+��ZE��%��&���5�C ����w�F���c�=�l���v�H�إ�%Wu٭ZmR�u;x����i���M%������FƼ57Y���_$Os�uI�����	fDV���̣|�^{Q�\���դВ:��W�nñ�^�'�Y����O�{ͻ���$�
�$W4\�7K˜���]�(�1p�"��ϱ�S� ?#�y@4	�匩]
p�o���z�góy�&��l�b�?�YlW<ޖU����-��qy�qAfw8�C�y|�35c�������Zxz�[��~+L��P�7nU1+� -
������
;|���Cq���#.R��p<�o��w��_y  �zx���L�d6Q�)c�ۆ�[m�Yr�\��69΃Hjc��3�vq���6Ɯ�P\<7<O4�~x)�A�e� ��F/~%do� xO�5�X���w�ZHO�5F�e`��N�~xߙ 9� +Izd�Ӣaa��MI訤�L�d�M�&��5h��ǣ�wBU��}i+*���.��B�ƞ��_t���
t���x'��-���y�R~V���-.=�: �g�/�,3i8³'mև����Q�#��<ƿݭ
H���3oz(wSgX/���5S�Y���i����:���z�U�xJ\�/��t�1n���'�������<n���ڸ�x3-�Y�JkK�CU�l�'��d�'Eϝ_����c�띑D����C}H�ɏL���g��\��#6�G�w��w#�	k�V'/��F�f��):8�:M3���'n=h��(}����jO/S���fXyO�r�&y=�`�9ѢL��,��H��aͬ�+F9�f���F��L��xI���B;�$h�G6�~=S)s �9�G��M�3��gɡ���Lw�*�j<��'6�Dn�����ﮡ�ʅ�"Ҳ�A���T \ó7���� m7{.�\4:��e>+.)#�D��?�x��O�T��J�}��5�0S�yK�r2ŀ�x{3 ���0v_Y�w�
+��T��l�W%a�������Ö�U��(NU�#�	��m��V��LmQV��o��ύ�re��*�-?U��z�)����.`��u@���k<�K��c�mu�E`��1�I�)U��z_� �98��V��#��?��;4�ˡ�.���BD|�f3���'�A���9�'�T��(��?��g�� "��*2*����(����n=l�����|`ǽ ?L?�@���ţ�{}��	�P�m� �h��'�$l�jO��!��UxU�[�K>�oYI�l|��ސ��'q�$	����(�f��]�/����#��I��3��PTړ���,l$��U0�Â���?��X��Q���d���
7��
߸)�j�D+��&���e<�ڎ�9����(���B����qH.�U#p@��q��	dJ��{9��{�ya�c�8[��G(1�L��w�s(�
��4�@�,���F��0����}7���Rg���t�w��S&�<��ZE ����׳Tb���=KJˢ�h��P�/G��ʜ�?�h��Z؄�#L��ё�I|���PF3M�C\ϲ*d�Z~V*ԩJ)�䳳�-k�ig�}������Jnf�3暦���=���W������ɘ��'�-���mr�=����d�jۮ���F�L�S��'�n*������*&�Ϊ����b�2/m���`�Q�?��D!��s���wo�R�ʞ^˪�>-�DUD��q��ZNԗ�R�����چo!q�"~��p���a�1Y����/�	�kg�[ �(�H;��x���~�5Xe�)��b��M�ڶR�?�<�v�����*%�>*B�m����톜K$8����Ȝ����[���(K���������{��zo��[ZI[7ޛ$��#cȘS�"��b�XH&)���N�c���o8��k*`�B�g17H�1���j�8
�S���}��6����PD��l��v#C��w`^̉ ����<O�����B�/X�$b� 4�H�Mv�����2��Vl��mlN�BKyb�
j�w'��\�4���߮ �.��x��zw��v���c��|QM��Z ���� h���F�Ex[�faPj�#���݃g�"��Fcj���6H����U�ε�4��jM�d����]�\-�H�?Q8v1��\��D	�Κm��1�����$}�1L�}��{�%���P�6s-k�ʲ%�>�0��7?�f����y����E�.�7�d��\�X=|���M���V��L���>�6�g�8:C��V!�uZj��0� G7�Q�MO�w��4za�I�j�6J�i_)J5���݇{,iA��"��j5������ӌ�,�M«7,�������M�S_Y����6��Fޖr�.�s=�L�����LN���Վ�TuΤ�X�l�佑�[���2� 𴦖̝�l<o��iuF�`�'G�1@}�KDm��k�ga��Ѡ�W��R#�]˝�
��NL�oH���$�O�U�g!K�o��1KM�Ж�u�~���pd��A��K������͞oU��ᔉ8��#�E��vC��Iu�v�pnc�TS*��Y\"Zľ"�w�״�*0�n�D�5�2�+���T�垷-Yc�JB���̨ԫ:�M��T�F�y���tr�e��'�4Kn�U!�ȗ:��~��r�뼎��-�Gf$���@�#Ͳ'o�%��~�l�}���=䣝�e)���;~�㴥|��:�4�����g3�٥��v��m�����[����v���|ݗ�&�������]Z��f1����,�~��%	c�8��8��c/��J c�"�$�ԏ�x�?�(|�Gפ;���~:2ç:褷���M߭H�"y��C����%+5�6'v/� )�r&�S�V`�ʖ����.�o��=Z�Xls��ҫ���͢�TO7Y5�Ν�CH�g��a����wEy[o)A��笈�k��w��v�EMN���@u	(oW��z����Tr��mr��7\9�u-=�;θ��~N"Q���-�J	����5�V�=��8��(�C�Ŕ��~��>���^rgP��za��"ǹ�e��[X0iv�?�����ϋ;��
ë�������2/�q��鰅��ͨ�$�J�S�ʪz��1��#]\Ӗ��yCs/V����pBo<�b���D4�j-�,�ԆQ��ݘ�����0���B{d9��Yh��į�j�R�Z�xSaf��JW}Nu�9����bob�D�@=�W,2���eX�zC5��������# �Y�N���e�۸��"��"f�k�H��V��c<��%wS4�J)'��:6��q\`�T�V���ς��P�9���O*^�Ñ`r����a�_�l��Eǈ�'D	<�M8�7��~^[��2�˄���N E��	�_�  ���++��Q�G��kӺ��b�����y-�����1���HYD������!�7W��6�Q���m��Ý���ik	֨�ai(;��eT�0�W1(��X����:4��n���;�Hp��QmG&�tf���b����:���e���+W�������v�T� )׭6:[>yt�1��(�n�����Hݵ���#r��:�5'��(�I���dd�?��*z]C�j��X0r��̰ �T���r-]�gH���k���k�C#&�����н��̤_3�P�*4b�@Gq�ep؈�I'�|mkk�Dc�+��=����	�S1l���Y�RSX�"ud@��*�WW�5L�Mɸn�&��i����ݳ�Z@�_��r����Y#��|��'Nz�s��wf׌����N�^|wz��6�X�KyfY�䶷��d�(nk�,��X��G��,ĭ��Y�f�9�r��2{�׹��;s�N�ܕF�O[l.���c�/{�������n#�f�(w��H�hj��	/�%�ԣn5���`���q@���eX�$���P}���I6jR��w�L��Ϙ�D�����uM�WK�`�?�%����W�Z����/�!챏���,��@��0�s�@�:B�����Ǻ�*��]��a]�L�@�}\|p���`�b#�8��F�rRU���`���;�U�J��8O�.�H�Q���R��`�\A-4\�]��/G��ڻ��~sf�J?���W���g��(|�E��g�^�s�5'��(��6��
���;��������풢l��~��"!y��72��1�ކ�}ӚL����*K����j�7��q��F���� z�H����ٴ���T@�����F�O��?P4-��}ː��%�%H%TС��*&%���J*o�t�W���P�=��4&/�$ۊ��ADpr�� ����<�3�5XS���u��}V���.�X#!�6G�V��抇�}�~���t���y����=;C����F醙�p����!~�X��'J1�'�p.��3i{s�F��ܐ��D0�'����g��z�C̲�N!f���$��f���4ʈ�Q���X��y�����ٻ|��'t���>:ژ_]�z��<�V�������I^��a����YZ���*��j�Y��m���A�J8�O����\��H�VF�����B�v̿c0LQz�M�lf���8!�qĺ���)Y���g�=�� I�~��u�C$�&�h��p�|�B:��Q��;ν�|�6~�^{�[6A[(협�;,�?�D���!��Z��2��� �U~��x�a�0��,�zt�KR�#�+���jZ��b�oos̊�����u��QbV��}�8���?2&��T�E2&���!T^L�x��Z�7�ض}*�-�].�A�Sc�X��t�UsW����i|s#��*BO-dzДc��S,������-��Q-��̌8�� ~+To҉H�W��_���i�l���vk�~m��G����=|�V*�����n�F֖�X�{i�}k^��?y6��v�տhL�@D�2	�oo�2�K1�+��=}�� ��ͥ��vB
o�v��"%��`�z����4 �$I����W�'/�7��+���/�BB$�<�k�:$�F4�XTU�.��hO#`�$���K �o;J:H�
���n9�- ��>�*�KE��?l_�v:l��2�nP�g^*m[,�Or� �����K�_� ��<C������,��W ���!>�v6	G��?SD����9q��o�C����<������d���� m��H�P�����X0;)��ܭf�w��746ې��8Bp��)O��G���#xǰD���s�B�rDpQq+���.Ej��D��sa�0��NB?I�u�a�T���u�jEoU'���
clg��e_C���_M_��վ�w&7r�wl���2�����?���,��Wԡ0�c�_L�*�U$ ��>��bH��NΠ0_�)�O73#5jV5�MW�<��5[�����"I���a�=�-�I�83�ܩ>���b>��'D}3s���ڥ���rj{�'��uKnd�Z�˩T���|�����2h�9{��K��/,���l)c;�5o$�T3��x�5��I'�s_�Kn��6��f1*���H��m�w��8����N{E�3�W��x��>��ba��?�P������w�C5]�bJWPث+~s��������I�CN��n����f,�����x�o�%~R�ꓵ�z�Hk��a�{c<�~�d�vq|+𢆾3Qwқ�Ej��dW��Ý;T�L/qY.���g*�7<Z���	b�f@�^� i� t|�3:]��&|��Arf}_�ˊ�/�������N�4������3|<t����w̿��
7�<(H?���Q���~,WB��F��b	N���0�>��@�h�
��B=�D)5!&�5���M�t$���}B������/mC�2qH1Y��ں�l��EB�[����9��i�nMU����/
F�C�g*���\7����ڿg���ӹ���R��<�P¶��I�6taŏ\��Nq�V�/�o�P�_2���p��kA���.h���bˀ4��̴���!���,5P�Ə����[�+�C�0W���J��G�-����sY��qT����q�I~8$�����;q�EᵴTn���!=S�A4 �b��0�r�wM_1n��|�_�!�,1,ڨ\�c<��N��\��U������J-��^L�W��E�fL3��oR�2�c	}w�-��6�h5	�\*H5H�ި�z9�?��M��q�<����_5e'UĜU����Y�k�r�ߒ+6*����w��ȎX�m��PO��n��v�wk5i�h�4֥��`y�����>��O��5н<lCW��ﰆ��������(����?46I ��G���֧��4��ќ��1��VH�z��T ��I"��)���U;y0�|�\~�J��b�-��[)*}su���	��j+�6���������n�w�u�~�6߼6�+n	�k����6���q�16��yUP�M��}"��\|�C���NK\f��S0ǎ>��_�Q��V�n��:�ӆ`�A�΋3��2�rE�W3��x���.�('��x�A��:ʧ�%eߢrf8f�,��1±?��X|�)�O�T�� d僪�0m;r�*�´*��č6;vH@-���6�'���9��U�>.�)�F<x��Gp��>� [5-���LF|M�7ś���p�J�h �m�-���S	'�(������.ɤy���g�Ȟ��D�A�sb���2,IƅC>]fu蛴Zr���H��O}��A
G��ݹ�����2��v����1���m�_�����c�ɰ!���ev���@`�;�)�)Q��Y��i����hE<��ܔ}���v�����i��jk�5w3�)w�B7<����ۍ�[�!��{Ize��o�	��
,�a`W��S�C���T�

L�ĳ���)�sZ�m?���a���97}`O��5��B���{C���/&��������@5��\}#lS% l�����E`L��O-��O\�@��
ࢎ{N�|Jj�@��W#���0	����̋�*�:��ɫ6^�xk���F��᛻]P���h����V�����/E =/�/R+t�����u�a�K��uO|ّ�:7��E7.��S������u���U���X�jk�*v8���Q8rk0	�	�	��N��>���&bR�c��[�,�G4��p��h��p��lf`n�3��<���>��L{}ׄ��Wl�6$.S����~x�?#I�Q���� �m��l�r�4��.b��$��9��*�Acv&BO)_ӹXAq�.�u�;�v�}�� A;��A��z�<�6w��샻�T2S
����`H�	�Lr~���o�>8������T(�w)O�h�2����۬�;�9U���7�6%��҂l���W�,��F|/i���ǧu1�uä�bA�o[����j*�]!\H�ͱ_��&q��#H���fe>S:q�G�~����v;j����"t���ȣW�!g����=`�;Y��҉Uy�6q�m�E�W�Ufk7��R ��	�^���\���pC���+�}����vX��b@ ];��Ǒ�^kO�&��!�V��Q��Rw��.�Y�T��B� ���XQ��s�1(��T����CSA�L-�J�>!>��r����6Q;�c�ˌz��PBCY�F&�����+���`�AL��Q�dN���b�E����A�xėM�AY�y�Kė��Ķ4&�:�s��������Q�Te���&��3)�bă
Y����(�c^)��лP�����S|�x��	;�����K&V���d����c�yHB�E�ݴ��H�[�N�E�܋S�ԍ�>�9�#6����b!Q������x�2��J�W�����!�eߺ��t�	;������K�Z�����l�,����7!��i��PD��a^��%�� ��@F[ll�эs���Á��W<>ɒ�	�yټ@ �YSG����] �lYI#�pӖ�Hq�.pi��ɏ��z��+��MۤC��
u�43�2^p�Ҟ�ޯ�����f�:M#";� 4�}�x�1��	����^��Mu��$��[��@�Շ���K�����6��)��üxb���-(��6�����3��yC�ۘ�K��RxU���@A���5T�_�א��Ɲ��+Az���7S�Y�tі5+�M�7�,�F]�s�+z�y�՝��o��>[&#�<�*0�Q��j#��P��٭%�9��Q��2�q�Ŭ�dޢ�E�ɩ��O�^��K��9�G�<��&�y�x��:�+(YPJ��j̿Yp�����ʦ���솾�ܢ����P��'\��0}�����:i6�}Q��w6���������ѢU�0V�&��_?/9���}ӨDK����L��P����~UX�q�Eѐ(Z4��[�S)��5jS�ي��ړ��<[[6��U�/����˝��<Q�,�d&T�ВJƦj������0C8HPh��9|��ƕTdG������LЋ R>�c;_}�%+b �v1��)�}´�X�~������J�^����^��m�gMլ_��8�IaB4�e}�X(U�*m#e�Ԃ�SM��yRr��n?�&�۫���V�V;�@�f]�މ� ��.�J���`V�mNQ'��8dlx� W�+��
��������R -�#�B�6���ׅN��-2�����Δ��S8�J?�n4{�ߘ�^��|U��h��JO����������&���I,�?���bG"�m!�� ß>��Si��Γ��P'8Q+Q�,pӤ��>�+H�W󐠵��������}k��o�a�;1)�:	PLU��	io��=D�ѯsD:~+r��4~��`�WT�OX��xYZ��!h�@�O��\�,C�p���10�QQ
�c���odN�o��cmqR����(�?u�$G%�l��?V��x��@۴�迕//)_�L�p��}n���tZjq!gq}����vn��O���VĠJKΩ��������gs%U�H��f��I	jR���¾o��H0����B�/	��l��W1�a����xc�e�a7��4��H���u��v�r��������㼴����Uh����^p�.��:k�m�g<��Ғ�Y�.�d�*1މ�US���`�z� ����)O05P@��\����9&����9K�Z}��<��%����oE�h��x}sċ�D*8z��Y4P��^ۘ�f�4o��9%������rmȱ���������L�[� 
��|�	PG|�){^)1���	�!o�_�Y'���i*����w�K=�?ի&�(UG��z/+_��PҬC�_-C׬w���ű�Ǹ�V��>]Ň�r�}��{h�Gf�,��V��|,붑C��
��AɕL��)�b�S�I��j�乀�7k)ļb�&���~5�����I�9K��a�P�>��r���RT�G�9ru�`r�G1�Sg�R�n���[������'�B�ZZ�p*���3����\Y��U��My������ Z�mk�r�I"M"��t5vH������(E��:&��ײF,X;�}HA��V���$ �c�]p�1{<�j�Ǯ�f�؜�q;ԏ�"kU���Oz�v]�]h����+��� ZPl��є�+�Tlw!�����=��J,A�(\^��ADe� ��LoQ����a�:a3���FX��m���W��Ε���/�N����N�g3tyAl���"y�<�"Y�}j
-w���30�iDc>Ҵ!Ѥ�;dW@�n+�o{D.��d:��h��u��Z���O�D�v�M��t�1�J8�v(�r�%��Ӟ\-y��zU���(�R��t,��)+��X�T$V���e&�~*J��{�C3CIr�8���}fP2y�M7nM1�(9J�/wF�x{�O���`��y���YG'�������[y��:5i���ɳ���vߠat8�C�Cύ2�2&W}�J_�A.�]��]�ǝ��|�����p���)���K}����k[�&*c�x]@Z�3�v�y�����lv~��Z/���%<�\�O�g�6ȹ�+"&H@N9��A��E{�������X8�(}oT*~�+r#@Xm��O���M"� �v:���np#Ŀ8覈#�ℓ��,f ���w�����0�B(�bW�����0]���&L8n�XZ8�b��s�L��#�`,3�,�W�(]� ��<�F$R���Z@�b�S�ZC8�O��q&�H>��Yg��r�V�3-�
�O��C<���O�#�/����ƈ��Zs?��["O��������Z��*�fP�B�{) �e��#� �l�7��[�>V��Ӄu����I�E�����o��>u4g�f;�VR߷�dg�u�b��
~.��^�1o�����_�27I��WÀv�Պ���#˽�}/�&o�ݓ�PY���FڑN�n��Ɵ �[G(x�m�x���
������ ��
�g���<��..0�<"�]1Z��Y�d1����a$@�0�?�n)ß��F�8�S�[�dg���D��y����˵�;��`h.�<k$Y�� �%|��\���$d�}#[a��f�B"ʁ�����x�D���y�3ٱ��xe�.(��Y�Z��U��ʎ�`\{�죺KT�f�PAl]���s���~�Q-�f�f�E<���7� 1���(z���;ĕ'��GɥH���~`�[5l>�w��c�0����Gy���򅹨��j������d���T u��8��叠`H%j��_oo({�y��Zc�VlE�76~kcq@��-e���B��E��7.�L�td�Ng (r�2ƥ���D�.��J��'wl��t�`��#v5�=���+@J��o���3�ު��R����\���
���w��F2��x��r�2�|U���}�pob�,Y',$�C-��������:d�i�
ެC�A�P��V���oh�'Dp�T���?y��\~W�O�VR�N�B|a�ч[��n���y�1v�a��Ss,Ж�K��ZJϢ9�{���w�� ��M�CR���3ל��*�A��f{j�H�
*Q�1�(�	vB������?aU���,85WA_�YRG/���e�ߞ���qk"*��qyL�=�4���B� �%�D��T����t<�ɀp��y��O�(�h�3`ٙ��%�M2�i�~��cf��/!˿������072���Us돭06��h75�2Ұ�A�I����3����2�1���2�Xm���<��:�M#X���]����'Q�E���O/�rP�9�|4�11Rd�J��΢b���w]*ب���w���rҽ�㰽��=zcV���	�[{
��ġ/����F8����Z�#�ٞ�rւ͵87y�~��ґ�o���U�)�v�;�w�E��`ē%�ZV����G�V38���w@��L�uj�8����܅����ȝ<$Y��V�=1X���P�+~\�0	'�0,h*W����x٣Z�dYO�{C�X���-���u�at0e�h��+{����L��.9���4����:ۇ�ֵq�n���\dǈH	�(�BI�̟�s*\^lD��3���4(��Wc���?��1��_�J˘R���GY��yP9��(��w@&�p�*��Q	���>�e %�S8`���a[^�k�%A�����ޕ}x=���I��B/�X@jpU].m+��9m�~�A���O�ʏ.ۈy����j�S�xT_O/7W��f��n(9��,�{�9������
��.�4+�Շ��I��Z��z*J���~�i�^yQ�Ĩ�ݒ�倖�J]�Q�$�7}S����k)�$����\k__�`9����u��7$�v�結c�Gs_Ұ�<g�JkM�+˶
A��ȋ���p[��ԕX��C@H���)����<g��P8Qz���YyX�2d�X@�uN	t%Ue�󆔍*�j���'8��A�)��M�eg~H;Sv��>P�ħy 3m�����QМ�nÞ�$�K醙X*R҈�>H���=�[61����z�[�
\�_��$W����q�Q�p�����#�R6��â��� ���G/� ���{�`��W��"��Vo�KKM�j��1�������3�^�����r���]^Ğv·�Y�|/ڠ���O��ŴXٯ�����8�[(�+��&g����D�F�X{��JF���x�(�B������d��D�MSmx;��Lȧ80:`������F��H�@7�Z>Ѽ}����[����R3>�+N3y)03Bs�Nu�G�E�`�̼�V8�6x�T-��H{3y��������/B0�k)���c)AvX=���0��H�u�� yſ���0�L��5g�A��o����jr��pJcDX��{��*���a:��eG��fZwN���90:)��.��U�w�
����y���ni'`D�Z��ׄ|�9.C�j��fg�!Sʊ�TTyiϜ8��{�5��]t�U4�d�&;��,vN���Pj�qXR�%����Syi��>��nN�^r��$�d"�� ���=
 ���5ܘ̨:2sfzmvDĘĩ�bC��I"rU��4�6d�գE���kTPI;�v�о魨4N�=�Y!�e]B`�5/���W�Zl|	&��[����:��ts�J�>��潿�a�չ���nQ	��e������ڀ����~d�3�(�U�V\MQʫM}Wk��Q�nt�E�p��ރ1�rE��NI�"�W� &�L��u��
�zF����w�5�RP1��SI��w�4��/�#Ύ9�YFz=V7��Q�0g��K��8���.���^��F��m��S���Ha�i�>\I,U6�R�hC.	[bx���e��I�ߙ�bJ��6�����+
5��q�tAt�7
���Ϝ9W} �:�ڻ��ґ�S ̣���g����$=�3>�U�ժE�-Ͷ�C���q'�u�Q*���f��/n&���3c�W"��D�_\#���r@@��/����D�JPzw��-�V,��S[�/�W�p�W6QG(�e	�!��>������q�u;�u�ҺzR��{W�6����v螂�������=3���=bX������%��-ܔv�B|K�wK�Y?�Tm�SY�;^��.���qR8��Un/�{��2��� �N3�txN?�WO���!Xj/�چ��*��[��85(v��`��4�V�rd�=@^�ɐТ��Ĳ�	��2E����D`�.�؋�T,I�Z�Ā�7�xҋ=��Nܰ���"�H�Iү��,���Y	0j��x�;���.oW� �6VG���1�ٞ�=''n9s�o���J���2~�]��=�$b�0��S��,���Ґ�R��)Z��J�����趆�����n�`` �F����|��6�m�R'�Fύ�gㄾ}��q��v`q��F�b���M�?a��66�Ѣ�L���r����]�9�#t��#��F0���"�X�=�ap6�a�����G�O�͚[nZ��h�Ġ3�lӓ��/�����6̬@x`M^EʳZ�'��\`�94����Qx�B��l��d�w���K����J��r^��� �y[�Ե	������@��=�6�*(��K��4K$��&���pGJ�g��"ɧO��*��/�C!��E�rd>}��	��u�,>Df"�NIpz1i���� 8*3�Yr���!��9���E��z�|3F،���&�Ӈ�(�m��0�nC�U��,~�@��;h�Kb��Nӣ��
{�̱�k��k/�<I�B+$��V�����&�8w�2uX�Vӗ��%�$db���{��6��`P^i\4/p�\��HL���!w|�]�	�;SX�7�~�}s��r���]h�ْ�;h��m`��a�$��ϊ�G��qh7���/�o�O�W:�L�
���i��t̟G`�íR
��t�*���mʱ�T��yT�|Þ�U��eTfѣ&C�\-���>�|�E� ��s%��>0cT,2�}$�
4a�
�'���I48�@�WD\�"�m�;/R8���>�lfR�M���9��uX(� ���'#Yd��eA���l���vX�0_|/ޫב�b���K���{�=��x/���$��ɼb���Fá�a�M�[A�n�= �)��� ��s��{��<�A�
����	�{��a`?1;���sO���{[� �{B����Y�s�������N�nd�0�g`�ݩ��=���>��[wW&�K�Q�k�~+���]8q�<�����I �c�y�� ���8��w��ʺmSh�s��\_O��8��,�`j��!�����UZȡ\9Ҋ@Ke�2��: ��& Б�|~.��Θ�2H�'��d�F��s
�E�r%D�1�r�Kc_�j��s�P�v�(%�+����.uC�q���<cӽ̿�_��`t����cͪ������{�`Ff��=ӣ|���o��Z��z�R0��A��>qACCұ9�jlH�~ ŧ�o�i>���x�KJ(���r>���v�>z�=lw�h���ͻa�,o(���O�H1�1e�%���Pbq�ܦ��
��(Ƚ*���19�f	���Oc�fc�� �n0���k��嶶�R�pu�.��e����q���\	;�m�&�5c��z~:6h-��
$V����~�.a�F��rm��#���?<=��%�t��
%ƾEa���� 6��0?b���3�L�\18h�!�6vm�E~He �\�t�s~/d�	����V�>���C�j��޳j,fL�nS����jv�Z�z�3��ylR�T��FQx���k����]�.�ʜ�����wS�֙ ~��lQ�n%n�ެ��˺\�eK�H{�5>\�h�l�{�9�Z��,_���	�{0bG��pTF�T�1��Fz>Mح!�2��O-�H6��e���s@"�8!D��]�d��y�V��6�gf�Aʂ���yAV��3R�>��z���ē�����GCP\��0Z�����Ĺs����%�2M�������?T/:���{9�\�ҋ����q�W'"S���ǒF�03��߽���8k��"����V�R*A	c�e��R��P��L܎��ӓ
�����l]�Р胊(��dĢ�NTz5�i�Mw>?���5��.)�;X0I�h�:̠#�W�W�N�鶨~����ŁP���r����ƌ�xp��i�ǡ��������B�O_��&���Þ�|i�pRf`ۻ�s�F��R�<�$�_8z�m�b��f���Ƨ�]����Q�fap���H�ϭ�Я�����A��X����C�1��D���� ;���;N��M�Օ��B��#�#����ji��I�\5g �߀��Я$���yQ3�.�1,�X=�ΒeǴ��!���DM��0��؁�	�(���������]����Xo����Ms��!�U4)���	�wԝ���Ȉ�kjs2)y��,X�ȥ����c�3������>��]4},���h��D�=�4���.�N�I���_'Y�IF��2%[K;���RezΥOc��Hr�����^&%���J�oh#ݒC�%�[f��3dW�n��9����5\��=fK�_1��ƣR��J
��+P�Ҳ��H����b��R>��%�??D��Co����L�k�S;��v�e��oVu�
��z�3����&�Ҹ,�Ť�|�%Ra�t/��_�亩4
��.���*�ϭ�&�=�#Nc�̈́}�Ț�`X|0ԍ� ����p�~}*�� �T"���@��C��uN3Q�W'��F�
�$Q!`���aVSd���0C�ɌR ?���Y�L�#�Qӄo��n>G�b�n\�q��ө�0Gv�*�m-�K��Q?��:;�_��� ����6
�-('b������/b�
�%G"��%)GOu��G�\���Y@v�4��n�3|�I���WI�|�t�=EW�qU���B�~�4�5�><�w�O���jq�����=s�uۄ9*�T���ΫZ=J��~:��GC��`0®� q�z!�J�d�p��Adl�T4��z��%m5�'V�]��50k��O���a��x`�Zÿk�z������FME���X�V���B��F	�7.�#ȉr�nYէ%VC@�� c�%\���K�J��i/���r`Vm���Y�5�}�砂���F�*k�!�k�4hs�-�Q4D��������^L�U��<����N'�;@��=���U��X"r����Pz9���N>!b����_Xг/~vkn\}.�:T}�JW�jW��5��x�GaN�ݷ&�T���C9��|U�,�J����t�O��{���t�]��O���M>Q�ME�A��~����3���z0��@K�Z,�ZF�l��d~z	�"qj��=�\ϴv�$��Gԯ3L4�R1v�œ}��:돝�]�-���?}��(o��P��źg��h@ms=Ga*��.+!��  �Z2��OJfn���XY�?:������r1Uf����'k���e4-^��!�q��F#`�%g�J�\���v��]�|4P�5H����-���*ϯ)]KA�5��V�T �lr6	����}{p��t�Dy^�iG���?!�0@���!�A3�!r�|~75V��t�{�7 �Yy��C,�ؕ+[W����.+}h�6dp}3��ӊ�����)VR�,C��WљD�t5�+p��ʣ�\J�q��Oiğ�d8����>}8����/�hY��g�ԃs0r6�Y}+C�n�x�]��.Έ��X43�S�v��"�����ލ�~+X��%+�B�N��(1V�~���=s1a�>1�E-^��z,y��!���
��['G|7�Y�e���,l���Wx����(||��n��;�8�w^�F�=,�e/�9����lK��&2��	��k�u�E2�y@�Y,�]u�,��n;�O7��ʄ�����N����(U�,_Ÿ��-�<�O�����F�K���.���HT��7�Կ��!'M�D>y��@�Z0�C?|eJ�R��\Y/e�|l�	�K�NZm�l�����T�=�^�w���`oO�|��is;|?`����\�f�{/OO��4 S,�9%����4�m&�|m������Sh�Z/���+��+$$�UU�@��٩�8�+����!��Q�?�N�NK�D�0lF�}�����]��P����ÁF?��c@0B���a=I��#9���؈��4B2myoN&@�C�X<�>�嚜4�)�]���]X�N�$��!�r~,`�0i�H��*�����j(6�@-���ʚ>�!�O.>�do�|y�E���o$''٧(�t��{"�����(LW�[�I���(c
�5�c-��y����VI>&�┧xJ��e�Q.g;��=���<x�A%z�̗�)Gۆ"�B�K���u�����E�g�E�� �k��h��I$c�;�[}��M@n��[�
(��v����1�����u|��0��t �ٖ)Iv���)E&�HQU�=�٨g�'�nw��h�R��$dl��w���/o]�Z׸ꮥr}����v��hyDɃ�p7����M��X`��ֻO�TҢ*�]�3�UR�t�@+)� �69+�b>���塙CX\Z�:;
t+ώx�$����S��C��������pk�ZZ�4�@^i� �_���O�t�%&�y�&J2�ѥ�{�t��K��o=���Fp�i���^FӚ�)��ř/�jkVgϭ�%���>t����KZ����X�4�^2��G���AƢF�}�w%(��Eg#�w{?�d�i�~�{�����g��7���i��U����p�߇�`�|���m��,U�/}��,n��;��<�v(l��>r�X̄�)�_F[���&�~l�F�/a�,av�`�&D�����#�h�����w	�7R�eF'�������e�e�f�9,���;X���8��Vl�L~%bV�ӽ[͏❙�%"^�AS(�{і���ؽ1.�,��.Jx��}oj�C��#�ơ9�ǝD%˔�����`h��K%�gf�"Ы�d�[��<O��D( G�n�,�|���O�����"�#�ș&�'>=쒴wF$v�9,<o�p���-��F@��Jjm' �\��nPp��>�G�� Rh3�X!v�.3�]�n��C����E?^j�"��)Q�Kik����yU��6�!x�\x~���'P���Lm��*�D<��c˶�D% 0g�Z{uK�J�h��/od�P#u�l�7��(3�Ջ����Q������B��eeB�Nv�7v�A �/���Q����|ؘd�Mn���v�T,����/`>��f�KR���/Օ��r9דy���{�TFyn�����l	p�)�~]�߰_�H�&���j�Y���bh��W� ���{�2cL>���o�FDl�(���F�T1���|�&��D��=ͽ�!��}�θ��L����HR�dYu���vI�_�@n�� ���I淵f�}�x.W�����t�AtW��p�m���|͆˃1щMsω(�O�[J�`�H�dB��U��@�ҥdUԣ���E�S��������1'�-�ߗx�$��ڨ�3F���S�;�é9���b�o�j�s�m��A���=���3RZ�EQ��~�i����"���=)_����V洃H��Ə�e����XO�{iJ�� ���e��@��HO��VH��o���:�kHq�j�� �����~�2��M�*)���p��� `�� ���P��Ue����@w%�<)��1�����M�f�4^���C�\��Ԭ�?���E]�)�v:��Rol��,r���	��$��o}+�G��җ�0&�^��Z?�N3h���,�{H��._5��Ôm([I����D7�{VuQ�(���N����6;6SAW)��CV��LݽlY'PIQA�_4�?
<0&8�Ɛ�`1:����C���rT,uP�EO&�s��~�kD󧸹�`� ����|s3Atz���4۫O0��V����K��9�ſ߇�Q�cc��q�x۩�U���W�A��,ͨ����۠�U�#"1Ԫ���LgN��7�m�TA-N'�h�J:��� 4m!��ҙц)o�H�V�u���y�DՖ��4̭l��io�+��p�d
t����cM���Ὧ����@�Z�v�,�d�������b��Ճ++�h|F��&�Y4Df�Z�mo�ٌ0���,�&2��_�'g�F�s�]3���,�y7��-�{��p�����������j�L=;޳���}�r��s�+ 8>���� �Z�To�;�K�-XL�@y�-_VN�F::I�n����W�aC����\���8�'O�:_�>6$m�}H�iRuP����/b��?�t�1� �"9�����1h �U��o�[�W�뗉4)�A�=m�����,%C+�p��8U��?â���+\h�(q�pޚ*�J�`��|RK4f���_�����yN���J��u�M.lI�#6 �%Z'A�k5���s�=�>�5��Q��v��s�<���tcܨD�-��x�f�1G�_v7=�`*f�%�L̱ȱHtc�K��[蹔�SE$$fk��&��4Q�_G(�w������穥'�p���o8* :�L/j��`�&�$�m�x.���)��%�q[bh2ԓ�J������~�J�kn�� ��ɫ���m�"������R�����]�oF!�n�!v�N�A��W�M3�%R���ٷ%/���p �`Hӎ�1����cë�F�[�_��%��s����&'�b���V|�C�hc�����K5HAZ� /(y�L*����r��c��F�t�����T�c������}g�WX`Ұ�@^�T�����6�ף��*��(�E����VX��^&s�R�i�"ħ���՗�
7E\��4X"-	�gd��>7M����S�e�|��(d�8U0��S����x�QX��w�H�P?1sE w|ٶ%h�DG�Fa�	�l2�Ě�,�������e�ƕ��(�x���x�Ws&2����!���mQ�yKl��^�^�s������? �a1!��%�����kU�96�G�K�8LcXl_��/��i_k� �% m�:8_�b���lډa�B�����)��Є���vL9<���=xZ2u�2W�
>ʈM���$� h��0�p�.�Zc�"X�*[МN���[R�'�#�|�^`ye��+��;>2�,�H�!P�׫����|WP`�Y�چ���9.)�����,���2fo�Ѧ�+��I�����9��e{}H��"�h�hȥ-�8�T3�Q���+.�ā&���'�W U��f��_P��O5KF�h���A�sV�{�R�uxO�D�S�����+��DR_�㍖%��N�u��-�����|���~4������ܓ���B�|X`1\�ߝ�
ТMp�F�:�DFX�nzZ�C�"����y��#T{.�C[�ܣ�2�6��1�k��fV'�5�c�us��A�2�*���t��斋`�g��طu�Pz,�Wϝ+�8�>��a�4�\g�E��J�g�{��r�ێ��t�����m~�NhI����Ip~�X%j�~�|9dD��[��(T˗��tJ�\�m������0�˒�)Y�!(
�gf)?����H�K�E��=�����g� ���X�����w�1�5B ���qq8̊odd;ԩg p�I2oe�e�zԐS�t#�w�yA���|�թ ��0��S�R�:QΧ3��������`��}eܴ��$�x�WZ��K��O����	u b��yR`�Թ+����?�h{�r�n�6$���%�'�' �}m�@I浔X����M'G����4[fe7Y��e)o.ӬP�KR�p�¸]��J��1���C��=�@�j��>�M�U��k��.w��"����Ŕ\���!�0ʡ���/h�L|E��8myp]�@��;����f���=F�O�6��1~�Ϛ��s�`P�P��E�'ΤN��ـA��sf>{A�W��M@{1�9B%�6{���@^�D8��^W|9;���!�%�n٭ɆhCOQ�~_�N[�&/HR���d
�z��V����&QQ嫗��� �%��I�ӛ]]��v8���k\FHR��t���`��G��9�6
QT/�!����
�#�"�u4Z�p�T�;1�S�Yk �.q&KQ"�;��L����� ����u9G��J����9�� E�uv��ѯ��j��[�)~ܒ���{|P�X������(��{ZS`��J���y����T��(i_8J��BAnEY��J
�a��Q1Ǧ�"�Iz���l�]E�_�`����{YwH�/曪�*<�K�2���u�cڠ����4��P|z��/�%�d�XJ�h�>g+ �M�^��N��"w�M�8�n%U�C.F��3�,M�v�Z�����:�����Cϣ>U�c?Q�$��R�Yɹk����?����}�ؘ�_����:S�֌K�,��ۺ�̞��%7�B�_��Am�r�4�b�p���@�$���2,Ӄ.���D�l�QL�,���!�(J����u�m�=o��͔�\Q��|�goX#<���(��D�ȊIE��������v*|��޴����k�g�b/Ȑ�����] ���r:��=V	����H�3�R��֊6��uȴ���4���ꥥl�{E�<�	�ȋZK	D�������MB�Ŏ��u��>|,F���iI+����1�{��G_;���U#�,��g��32�s��l��I�Ml:�
�/��nk��ҧ�[B/^�0J�/g���~Lt�����6��"�Fo��\�B�U�b�8�#��i���[a%)IP�����/U��c.�#�5�{���/d��Ʃ�=i~xq�T�=�j������4BbAKs�v�E'��¨�)W@5��%⮺�A�S:x��!^��h�-j{o[hѱ����(��D��R�-��뀸�~G��XB~֖9�vl �"�D��V�	�S��U◙ǌ8y����7�[-Mң�	��6�����mK�����h�����Mֱ��,EWdm�$�B�m�v� Ϟ6�,iW{E�?D�F��%�hV�zCvQCX������cB��W��LP��Z\~�~Ǧ�zٻ�'��&t����5�8@y�4�o9����Sx���-��S���
�[Ԉ�ND�˓J�_M�ِ�Q�x~#���_�� �,P��qP�'���4���a<�Ȍ�/��S���!�ذ�=�=z�� jǗ�ּ�I]��Z{��y��y��l�	�~
�Q��:��1���QV��j���������S�'�#�l���L�d�Uفe���n�ٗ}K�v�nI��$����5��T�GΌI}3a�%��̻oA�g*w���܆��s�H�q�^���}#W�kR����]�4����4{/l�/�9�NXZ,����_))�qr�ׁ��5�k�:��fܖ���4�R;o5V/�
�'��'74�g޲���".H+��~?MaOE�v���c�s��F��!}�{�?>�N�{cG6��ң��QṚ�We�����7z.@&gy_0o��7�zϤH�{���)�z�����mV��Ǽ�[�k,5��V$E�P=�oz.`

������Anr���d����qp4؊P�f_6�R�i�=��I�l2g��1~j����k��M��`T�k�g���Kkn�JחsG�{w#�P(��K�K`�檏�l�5�������H�"���5����(񀓻��^�H�M��[f�e'�ϴ�$��/o��͐��!�&z���e�1A�?�{���A������D#w�X��mЮLIN9u+�q�hdFa����ݰ�1̐���~DVt�si���-~�0�S�u����,��P�_݉����mz?q��FvAa��u�{{��ߍ/H����+�����$��!���`�D�*�Enn�Ѷ�+kCvj�T�-Oe��I���ӟ�Blop� ���d0Ƥ�/�D�4�e�/Tr�ux��&���1B}����\��C<}�U�Nִ�g��e9� ��`B�����N*����R�~#J��㑯�k/\܂�Әb>D�����Ā����Q���EF��zc�}���Y���H[�H���Um���]���)k2o��.���K�2q�L�����o�5�Zu[�V@�,�z���&[#�%��y,�4@����n�����p�r�{�[F%���,T
�O�I>rPRQ,�|�=�z��p'��a��Sڋ S����!��z��}=�r�i�P���92Q� ��M?ʥ
a���Tj���-������AA*ΦLB'�a罖Jź��c"'81��h�Rnخ�9�%"��y�sv�&�W;�h\v}��C@Ea{?i�	;��^���
�Ł��ު�.[��ժ����a�1
0��r)䋗*�=�`?a���N41Qd�;ް�����������H	d`�l����$�ljo�C����f�I�����Q�)�0@�!��Ѹ������0�D#���<B�e���}�������X�����\qŘ!f�52K9�g��@��߁r�r ��!��1U�e��ĩ�ΎS�+c�����[���[��;^Ͳ˝��^��E�p�Y沄��)B��_��O����9�t��İ��Y|������s�c�Z�D-W2i�=M9�T>��ϟnU�6���Ɩ/�(��8���Y�D  �"%ۜƒ���W��G��/�G��#�P]���î�n�����\!2�D�Avk�-;�-��QĠ�Щ�s�c>�4�_!�I�*bN�
kD�B;C'��9*j���PR���E��a�/��y��ͳ��u�'��M���'���Ō������V�BL��s�U���
�V�d5x��0��%G]c�5�s�q�^T�}�HT\S�KC`��cO�p���+���&���{%^��0�<gZL�)�'��ډ��$��p ������Px��;�Cqce�����mD�i�>SJ"D[L�7���Z���fD��{��ᠼ��� �2���Xx��Ԇ��M]��9!Xch7Ud�noƓ4�S���]4��Ne�M��o��p��x�a��\6�sMh��i�Y2e���Я��J]ތ��3E��[W֌:;�>�iU����@�՞vhe����w�JT��;J�"�n�~6�w�4զ��zucN�^w��CP�C�	���$�����)��$(.�F?@�4�V;^��-;��4�7���A՝�;�{����f�Y$/�����;�1�$>�he���@>��4�gǇ8��a^��h�-}rEKwdGg,�u�nm����FQ���:��+�M<�id�]yob^�f���S���z9����En�e�p��S+��7g?�\- �{���V+��mu<��1�u1�"�{��w���u�wY���=�+��b?�l����E�h/n��O5��Z�	�c�N�V���o�h���죋� �Wӌ�qx��}��R�����E�B?ݍ\P,�&Ԡf���47�>^�k�Dҏ����[m@'�Cz{|���A����~>��ı~vf�:���.�۟����V���Kk�®�����W�Ҽ"���y�r��(MR�3��[����!U����u*����b�9 L�kq�t��vr�Y������I�\���խfR�]ÿK�U����{���L	��#Ҹ�B���Qn�Uj*Cf���]���ŀ�I�_@qE3�����<��'3-
��4�" ����Wf�'���?��<3���Z��f�Q&�K�>��p9��{{4�rK5�p��</s��{3+>��Ar�c˷7�S1͢ ��?~�	�O���QR<ܧ�魆�dzU D�u��=A�m��cE����?*]���AE#?pG�]��u[�傢-��ÕN�X(��q���qj=ߣm���:��̽��/����̾�Du���7���������U'A�����M0�����C_�B�t�P�@�}������aL�F��(?Y
0c39�m�f?�bc�'p ���U�F��j���I7�Om�^�v#A��}��l:�\׾+	(T��:�OU�Z�~�Q� Z(̀T��T$J����9��C���JM�R���9'�r�ҿ���	�R״���/C/�Dd���ZQ�I�Eԛ��)|���!k.�ɸ#�ԋ~M]�d���g�G!x�T'( �S������5�ו�x$wW��������3x�������(C,�XnvS��os�����Ìj�q�ã��s���S밮=9t'^ԚQ�`>K�b�p0�����u�h>��0V�¢ɿ��0>���;�0xO:�qS~9H���EK	�y��(%pˀև2�ce�T����E�<w����!	�msGGZY�4;=�e��z���0Z����l��/H�>��3�ͭ�K����{�Ʉ=��V��{a��[��q�'t`2O�<�e9`Q��Ϋ5l7�k�_��h� k�n<d�����J�c�
�j�۶=r.PZʦ�F��}�^��8��P���p�>ڝ�us�5y���d6�����~�z�����Jl�fd%X�.:Vn����ġ"e:x�uN��1m��6��鄬�b_�v=[W��6��F��M��ҡ7��cY38%�9��t�0|뾩E�o��I�3n�yu��Zu�V~�MV�'ԳV�����9��t�TK��0�4ɰ��8�����i����$��/�X�;F��xC{��Yi\�X� )��0�#�S%��E2 �q�R}'�	㾬��t���$����^���2�+%��O4�~fk6�$>�~l<�ۏ����_�G��~!����Fs��}��(0��vL//�@���!���l�48��
E����Ɵ;<�64�u�NǷ�\�7[��)��F��2�B�����+�`;$d�hLa8������%HR��aW�"8�&��cu�?��L��Ee(�H�� �Q�i*���x�]�fa��_3�S˹%q� JwY�8��ؘ�}=��Z)nҸh�׎���P�	�6���DƊ�ҕ��y��h#�/�6D���>J���@��M�*��X,��T�6�R/f�r��^��4�ԣN�~��	�y�^P,"ӟ�\oӆٞ��+��W�f�c�0��͐��2�7��;Q��3V��.^���d'��/�K�ۥi�d��)����s@������ _�>�*��#�. �d)�2i�;F`Z
�/IF�Ě�1����'y��n��Q��-��	��q�7�����I����|�/�=	!o������Z~8�woB�5=�]�B��,�2���]���bp���U� �h��HZ䲉�_���
��=%�9b_�`�3���ڥ'������.������I��:l:��d��?�Al!d��~��\?�Ac;k�Y?W&���Q��$n�@nd!�2�������F&x^ ��O��0�@¸Knϧ��1*�9��T�c\����&Z8@k�̺n�|��ȡ[cT����Z�HFT�:XQt�@@׏� }$:�Z�<����pC،{�uG�=�ǀ�`�?�B*�Y=�(fc �;���):�Ћ1Q<�İ\AQګAH��=*��Z�8�A�c~t�Ȑ�hh�%�P�IE��*w��ˇR��ma�S�-�MT��ʩ���>ۻ�Z����Ư�%5��#B;~n��dxS�>���:�o4,��|e�
`pZ��N�>�F��~�ܔ�3C�#H޺�X.�ꪁGW@^�NP����Y�$�k�����1����?b&Yd���1�3>=�5\��D->/������v��D�JCl��s"I�%�9ߜ�yL�D���ڲ>���o���t�sh�G�U�QM�Q����[v�פ�;�p�γ����!'m��Y.�mI��=F�����%�A�n��
Z܅�@�T ͊R˂�mP�6@q�ΐV�𩌄U��F؇{�f�RN�d�<�z����z�,�t�}��	dr9��UV�F,ü�"�����̓5��h׌���*oZ2�zF6��\���w�P�40�O��*۹�S�cH�A�M�c'��+���2~E���-4�:0p�L��U�0�2�
�<@�_�v]0	(�z_[�V����%6���{X&ѱk_��o2���{N�/��x�ϯ-F�|8��(�b�]���M!O�7J�Qͥ|!~Φ6GU.���Q�;=��)݌���D�}Ӷ���~X'*�0T2@ׅ���'�'�;��"���j�`�φJ*r��P���@�y֑A��z��N����~sc�zO0�IoJ�4q�n�Bb(��m�m'Q,��c��D=imT;���x�cO�3ǝ�O��3�TT������h7z��|��&��n��-D���.uF���(tL����,n��4������;����0�D	j �.�\�_~^Zv:jY�4�p�D�l���o�t:���S�$�0��K���9�< ����-J��������[����I�X|��gb���Jf'>3b����\@����1��[����]��*����c_���F4�J=��|n��11�?�'}=9��#+��b��h9�D�}T���L����~��;��
Ǯ�a\�8�xQ�縻�"�����%�dڗ�|'a-N߇s8�������b.%������7��~Sd^~�j�*@ۨ`�N�h
�f��P���@�߶O�Eim���>4�����G� ��Z�;����O��+�����ڼ�z	ڰz�G�����4������ek+Uv�À�5IϵWàĚd�f�G�(G�'��V( �����Ld��9��M�?��!��V����[]� �`�KNo�ڣ��"������XT��H{�μ��WjHƛx}^�K��<p����co���;r M�TE#�ėl�dt�e�ʹ8�/.�q-��<�s�	zbJ���j�cNbwZrY�+E�$΁����s3�txֳ�twǢ��^�>���톫ٵp���W�E�����%p\Wv �9� �4��P�x�[�'��@Y�� b�u|%|Ȳ̉�_'h�s����%��j��e?�:�u!��Upپ�dn6!ܴ�l��X�B��-��ӐI����PZI�|��:]Uf"*/�T+�$ZÓ�.���)pT�ܵg�#cX�5U>n�����>�Нnq�� rc
i[e�2�H8����p�R���K����\��O����T���"1ڍn��FGҙк5��F�-�:ǆ5�R���<����x�Xv� B��9�y��Ye�iۙ �&����N ��`o��:�Q��KH܋�P�&T��´���䘉�Z�P����C�f��K��54b��=��3�K_����A��n陌j�E�P����o�&���e��覉>�5��E�����K��9���A��S5}c��h-�a���͎p�~8Z��S�]�ԇ $Z=��/�R>G[X��R;�<�@��W�+i�����V��&T��fN��cs�B�8a���R5����x�o�l)��Rb2b��5���ᒜ����T=���@}���m��E �Jo�������=�_���Y^���E&�
�d�q78 ����^��kCo�����+�y5]f(���m���T=;-+'쥙]���]'+T֋��^��Gm�6M���_ݳ��D�V��h	Ґ���J<�V�c��"g�ren�-����7�S�R ��}��y�O���~҅O�	��D&ό��@b�`��R�lxu��i�E*�}! +�p{�v���ф*4b��b��̺�{�p�8����D�Ɓ�|cU(�;��>7'�ߖ
�\����A�.��)&���E��Rlwi�<�C���x�t�4(Q=�'�J����6j3��w��P,��+N4��Ȣ����ɷNa��5wץ��lRZ��#�	/����}����hTlC�%G+���])q
*�A��:�^�l�ߧ%� 3/A?C }�vz䡮�b�� ��EP"\'~�h�� ��VB��D-s��ny���ʼ�l>y/�f4��]D<���͇9�P�"�xɰ����~k��ʉ��71�kx��0���V���N^���E��y���> S.�%�"2�w�İk�����o�1���z֫���=��OЧ��zf'�^�SA,l"��͔2��,��ƀ�q�7�E����%7°/����X�+NFZnLqy.�Nב��RQ��U�s��t���d���Vl<���M`�<P�4rK1:�rf�K�a·�"'�e��'��#�%������M���(c�:�p�E�fp/�5�; �Vՠ������Fx�?�<e'��y�x�r�.���˒Z���$���E���ӹ�Ǧ�'c6�ae}�m����t��ue��_<���Pu��RD�s}�D�[^7O`u<h�S(za�C��kc#�o� �m�T� �0�V��Z��Pbv
%�g(y��[�bv�m����#C�n�SV,�� ;�?h~zϰy�����|�[��<2�k+)�ȣ>�����j6-%�4�����D�A޷��Q5_�P���k���֛����m�E�0��>��u}@���v��,��&�GFyLl3q���2��WS���Ԑ˛�I�צcuё�*��:Uh�W}��.�� W�'����Ű��㗸�y饠���ݍ�֚n���Y�Cǚ�?KJ��k�m:$E5e�����J:��	F[��~/�{
ҏ4��g�'O�]9�A����`m���ԏ=(Jٷ䲲�K¨d4A���s<�a�nZ��"^���v�^[�R�Z��D�w��A�B�.9Gy4!̖��γ����7I����u�Ɵ��((���FpZ�+Y��[��*6�{�ߴv���FM��t�kv���	i�אcL>C���!�1!*���a
��L�v%���|#�-��1�WvkB��OD7�
Qɒbc0v[ٹ�۸Y%����/:����fBN;�.q�3J��LF��������A������N	����ն�:�|�h��R9d]�����#>�WDA��<�3��iF>�vM*�� �0'R��f����T:��w�i�p	���v��Ws�����GN��\�� b�}��(IQ�G����Q��'���O�X�َ�_\��;�dx�e2?ṭi:z�h5��B��*�SٔK�_R���|����*�n��	y�+ �2f��´�US����ԗ��<֓����!��!��0�����|��d`J̄�� �6]GnUZt��y	�?� df ��l�ş�������o��Gi�K�ز�	%FV!]�B(�1�&ܽ"2}^�ղӴ���M�^j
���%�Uz��d|�|��m��w�џ{0�%�u�u��>�g�1�) vu���y[��`Y8%�Zk�p�!���U��mOo(}���Y-�L^�R\o�EA�Eqtjɣ!�x����3U1��i[=sT$H�!;��-k� ���5�ʬ�J�K̶I���9{�h38�S�f�X�-�ڋ�j�$�v���FAF�EIu��T��W���>O�9ꄠ�S�O�(�&�<9�w|O��\q1^�#`ݘ(,�4r�e�HHE�&ǌ�l��Z/�mծ9���/+�hg��M5?j����+Jy3�m	���k�h��W{ 
��L�0�����lZ� �Ժ$E�L�`�%�4.0�������bS@	�-[0gl���I�U�q��C��ڲ�����9�=B�z�!yr|��x&{&��}��7�ɡ��=Fq
4$Λ�B�& ����D��=���L묂���Y1�=B��44�r/��� C�I0(�?�v:�&���s��z�޵����o�A����Ӿ/�B��KA���<��`�������`fx�,)۾��q��_3��~����z����K�ņ8�n^�&�"�%����7��?��Nw��k�z.8岯s0�������:g|+���`Ռ
��'WoB����@�jO�|�M��cJ���,@#q�>JAU���jЖ:�.-�3�]J'��M�B�̓���4�Ղ�۪�/V����������t��3O�r�o� p@�Y�g��s%�蘎��cnB|�!vP�e5G=q+@x���9�	Y`J �S!���t��˭)��$|3�q$ �P٥Z���}S���moc�O:��� �CpcK���w�m����#"I���"z;`�x{�`AE�9#�O���\���eKED�1wE�
�2� ]R���
g�E�Z;�����ѩJ:�!�"��-3gB�\�B|�9�"&_�g�&�=A��G7wT��c
m����/q2t���ơA>��iwʛ��IxF�k �v��[7IC��r"���LxW�DD�}x��1�^�ϓ@�Q��1���&t'�C�IT���C��%����<������ŋ(p�"��j�Oq��dQ��aF����t_s�i@�����o�=6*}��ɘC�{*�Mtޗjf�
,rw�O+���첒�z��դ12� >�q�J�Ek9���F�Y�����/s���{�&y�
����&t�x���aBWz!����q`6�4O#�yKcE)��]����M�rf�����Ӹkh�`UT��N]�2�u�T	��������B�u(q�����}�+Y�
��	��~���E[�������o�-��;1�Q���������"W��oV�7�(?�|
���b�Z0���E�W.5���"V(��N6�M]޳g��,��0S�"_��!�����4KU[�<�H1��K,�.E_�5������XM?�@���@h��K
U؞_zp����UQ�e^9I�K��S�!�����))Xa�ͭ�kq,!�K�0����-�8L�ȋO�fj�P	?��w���k�N�1�[k���ߺyS�Vn*|�أ9��L�PP�а��[[.�����	�����7v��§�DFLۃ�i�7]]���O�ޮ��\���ۿ�$�r�k-}�{��c��]�/�Dѻ��:�A��C� (Ho��9��J� ��5M%aw�S�ğpW������/%�b�C�<r_F�ڙ*�r�:�X.�=Ƿ?����Y��"�����ָ�Z���m���ȇf@S���~]�~�LoL�H�R��^��y3����$<�҅1��I��s��g����R�aj��"fK���阽O�ju���d+�����ȕ[�k����1+7˻�uH��p	ݵnFAXD�'����I�9,>WB�_�n�t�<��ҟ���o/$F��^��F_G�z���A�j�U�9e���Ú�#�4��4)K�/�pJ�]vLu��UN�z��>���bP�NO�Wԃ��(g�t[������0?�#*]���˩ !��]��ʯ�\��A�~�%"yх���+I	!��G�ȫ�z��K�+,'�mۘgѭ�O����>/?�T�/����5�F4�L1���s���<��I~�g����?����~��M?&':/S��L��/Cao*���U�*���!�W����R�	�6���lb�4f�Ur�o>�5�ح°A��\RTcLUM�wս�l��[�5���
���+7ԥ]@AE�������Ği��+)�}n{=���6��>��Q'�;��{�L���)���jȁ�;<��z5�c5��$� �X�4{����D�;�y*6mg��T�(�ӉՒ�y�gS�VT!�ĵ���CM��R��o��zP$[��`M�*;��'b}.x�'��N�HU��d�A��B��LCk���@�@��������Qˤ�T��m�i�1y�d3�9��kk����J5z��@�^����B	XBڨ
a����?h�$�p� �q@t<u���6��1�tp�s�}��R��'�����_�P����9�&�;�N�P������W��
>��d�mjD<y\�Q.�!�!�����PqQX����ˤ�)��>cV��&�E�u-b����=`����֝_�F�诜a�s�S�ᇧ�V ��T_�d&��y�f��-�?p�]PC���w��3W�.�2P��l�9뎅9����q3�4^R��^�Q���d}�;2���kTY�\xK��5�<9%(/���CwH����B�Z?�h��o!be>1�~L��Ê�� b�dwkr�/H_�����:j9��W�)���fз}b4-+�2[�Eg1��� �ü����[�Į�- ����,˻�6�^�S����u-����+N�ɸ�"˺�Y+`��+q�z�@p1=����	I�[8A���̾J)�1���r�N1�5���L�mhCC.m��z��K��YG���M��)u�ѺVAӻ� ���}�f��G+/(�?�� ����
��qf2}��Mm�[�1���R�Bq�Ű`AQ�]6���<i�Ly����rH(�ppct�z��+��HH~Z ��Y��i钞^��F�!����Ғ�� ���p��?*�M���dYVA̚t{
c�>�0M&�˱e�\q�~��lxP��]�j_a����A�S׶A|����V��J�y>��w&k�Rm<]������F�Ɉ!Vq��=��u8jb\���X�i �6�W��[^�MvD�Z�W5�[����ah����k7x����J>&���=�����ل����D[�"��R�{-j�?Z��'w�W��"p9�瘑%�Q�i�|�.⭛}�aҤ�m`���FL�!#D��,y6i��@�{�Y:�$�4�HJ�D�jkoa�3��XIN��75�S]6Ee�9^a"8!�Z�����5�|Fұ ���Bt�"l��� ��R���>ml��h�#ۓvJ�)��S
��7��U�����v�~��q<�PJ�O��U�'��B~���}R@qt��J��δ^a.O�13�Cйҫx�3: �H�8{c��K�?�UH�m4Sn�a�R>ѹ��D��|#�Mh�v�_�5��6`�X�H�pGq 
Tɫ��2Q�&	��U�-� n�ۀ�(xي�\�|����b��4���Qx�����&�TQ"E����O�	���Լ=I��7؃�eנ_�v��Q��C&��1�����yJ�G���B�JQe?�%��͍D'��<�zy�C7���M�2LU,�:A�ii�����5�d7}��"3�ZP%�%���"Em�?�M�Ț	�R��*������b�'s����o���̐ G3�9A�poɲ�4Q�񆠜=�����}l�ӛ�?�=�oz�E��y&q�G�'K�&�� ���6�2��.�P�j?O9����a<���o�eƭ������$*$L'��1>����8��^&�1�~�br<�q��{V|�M����ֹ��3�y��z�#·8G��^RY�:�/]���g4��^ݚW�Zm�==ֳL��+��^�x�av76\
h�7��	b�Z��I�wf��r��Q�0��ë���U�W�S�k�]�]jp�vmy�_�Y8�`�o`�M���.W�Jw�2�g���΋��A�'�� ��t���5_��f-ʬ�Ѳ��Y������s݊���ƚ_�ǽ@�n���?��^��{�\�\y�೔o~S%�`�.=��f�cy�
6��>����t��؎h�"%�)=U�s;>���d�PBV��E�G^�U���0�LГ�_��̣�o�����@�%�a�Һm�	��wU���EkSm�8N8�3�w�&Ә���$~��:�Ս4_��0z�N3�
e)}�oz3HE�t�$��Ƈ�Կ���ɩ� ��p��A�U��/��(zK���� \m�B�n�z����2@��N�S���0�¥�W��S�TY}���]�U`}�t���npI����Z��샖����W"��A,uo�n0�����_���6fk�G_;�/HN_m�����^n�H�a
/�Ԃ"�註��s٠h�F�J��xE��p��L\�Ĩ�N�?A7�̔�Ʉ�������sq����d
�tĲ�E��}��ߒ/z�L��J�(Bꇂ*�Ȓ36�p�U�ON����qJCl�2B�{�5�*�w�h�#G��S�-���	v����t��&��>(s�%�<�CM�
ρ��x�8�a��ǲd�7\�˝�F�9�^_��?%>��'��=�X���3٩!��֝���d�f������W3rZc���Ylo��Z �i�sJ�NMC�"b���4�����Ơ���gJX��7�1��ėk�	�S�$.k��_$N�?Y�W� Nx��@�_�{c�(黉#2��5{����H��G�VSClb�^�N�0��ew��a���	�Ȱ`9^kd�{:��%�!�-�!�d.�X�������.#��<p�7�G�������M0�X���e>��h��IP4H'��0ͪX;0�֧畚h�,J� s���dc96����kRn�	�'�1}�0�'��Rt�:*�Ӡ�]�D�;�z��O�g���K9_�ߒ�?L�*�(D*!�y���E�/O�z_�ϝ�������(OpsW"��~�;�KB�T�µHF����r���a� ��|����.���w9�,��d�d��GI�h�~�D �Q�y�0q9�`�p	~�q�1���mk�ځ��q�yc��Y����G��)m��YG�������,6MTt,��y6ir��ܘ��ԗ�ʷ�߆S��aB�x�o�Iz	���'Nd�?������ס�1��Y��kٟ$�g!�o���w`1���H�����=M_�$Y�^����UA�a�ss��r���łB�iݱ�w�T������6������1�h4����qi҇�q��|R�1y�>��z&~D�rk���Wo,�[kkI9H���4��ɦ���\r:�n������fT�tH���4��w�jW�'nʍ#ܙ�ZIPcC>j���[�[Y{6&o�40�Bjt�$pG����V�Y�/���_
�K��p	�����(�jpW�7^Lf�%۔Y�����[����xRó,Hik:0�%����oS��G"�/^˔��Z�b�D������b ��6�}N*ٴ#��Cdm�Ya�j#Q����$�O�$�92ڏ�bP�E#m�ʓ]�FF��,8}K&��##�9@7Nhz7���7#��s�)�}`���B�ɋ��D[��!f�d�)��x�ۧ˒&�R<y�|�-~����S��#��H"7�]RE�?�Cn&$<��������Tq�4�y5�-�w��/9��U:�(��	�$���Y�u��~��<�� p+�ÅQ� q6�CZIn��E�$�Y�}�H��g"�J�pӎM+u �.��}5��s�ڄe�:��*P
��c��MzZ�:ѱ3(���Bx��0DI�:6A���8��:�L�+1	6�z6�{8����-�:�g%A)�C����̏K�B\n���{Rj�[(~�#��ALa -��]�>��~��.���d�)��?��E@�R=�e��Z��qoT��-�V2 'm�pєlJ�����j�#_�:��)���1�c��L�4.�z_��O�O����B���n����<&�#o|Z��l�P;��%^���ͰCsd`�ꚌW� �����;7�z�4>�Z������{9��۲�t���)�y�G��-�S�\*�)��x�%'��	�ӣ�L@ ���0�+��Ns	�X�R�8��Ջ��CJ��D��@���9k������N~w�J��Q"�bו����6S8,6����_u��d��Q8�:�;�]F�A���W���"|�w�i�O;����U�l���9�����e�D������XNӻo_�;TvLq)��=����|���Yĸ+)��YBi��8?�p,5�����Ag��r�@+�)���| �z���>˫'��G�&dȖ7�lg�Ñ0٘�U׼;wׄ��u�4.4��� ��+�'M���K����]�Ӧ����6�"L��/��P7K$�m�v�z���X.綠��H�@E.����L���z|Q���-�y������xF,\����8��D����*q��w�c�Ꝇ��c�aes_�̨�=�g0��h]�z�X4�$ ��|���$H�.�v���Cv!���HBG¦�P��e���{�#s	�dQ�+�i[=����B��)����t��u�@��`�19 ���m����ّ��G��>�U����u9$��M7�<&�Ba����*�rM2�ēz��NP*�AT�{E6����ߐi�����.��a�T����Do��'N�\�?���G��8?��ӹf`	��;��,�&��2�f0��1�X[<=?.��!�j����3N9��P�fB��_@���d���co����%�v�n�Cw�6F%�1�J����p�JFjڟ�Ƶ�v)	�:��1w�q7�D�߹��H���.Tp������Χ�@jX�H3�eCUGKn�	��&A���l�����&*>V��%����
���T�K�����	p�gtk@��˛����k�
B������և@v��H����3Z�j~����(v�:T�V�u$�`'���[p��Y^I�۲[�b�r��*m�M#�L~�ݾZ�څ�!~����vf��Jt�m���i��f���a:s�(r��B�@����S�P�4���i�L�������x$��G����.e�"B��\}P�d ����+M��XŃ�3/�������z�X�gD�'&eظ�q~枆���ox��qJ�|��.��2^��9LP��9���e�q�:Z��u�~[5r�)�������2KҴ�=�P���x����Z�_�K�V;(�����_�m^;���UCK���AH��t��A/��@��<]i�#
ßG�^"
�BfT���E#�(J��k��¢��VZ{}H�`��,u��N	Չ��m߈[O�6 [� �r`��#+��H���ynբ��Eo��2�
;4�p�{�"g�%>�']Ϧ�f�3�w�^��+C����2����� �Eh0إ�u��49��{R])_��S`��t�E��{�;�{�q�����甃�>�&x�&�4]��-Y��7�$.�F��VmD�N�n�s�~�s���n� a]�����d����J�<�@{�������c��ľ-�ф�!�먽�Y���g`|��mqV�����t	CB�2v�"|G��֒;��k�A50?^�]��yk� ۪��3��˱����f!{�����]��@a�K�#s��i��v�(w�<�F�B*��NKo�Ӛ��ں��'x�<�O���.sy�o��:��p��\�qs��2=��5/�B�&�V�kq�����NP-�بz���D�Nw��2v�r��E�{�g�� �%�.6����dВi7�2�Q��.nM��ck��5����,NɮWᆀ�D#jAlн�iQ� ��wWã$�F���#�Wbm~�n���=�0��zV�q{�����|J�����������s�Ub�l��N<�)y� e�Uij�����
�w�`�������kW�d�)���YP?����g�p��4ʲi�.x�o��(@��K����6��;xnO9e��Lh�����W@o�2R8��te���V����Q��}��;2���?����N�a
��u��b=�W^N},]M�b�$�h0�;�,!N�o�5{
�eׄ���P�&��ܧs�	�?
����6�	�ܥ�P!�t��\c�M{��l-��AN�%��!.�}�DҴE2�M$���o3(��Ā,cJ����k������zv�H*����m�4�v�|��R1(��@�_��Nc<�a�~I��9��
�<E�kI���A�"v>~�f�h�@�8��Õ�o|��̧�1f9@`MS��f�@��7s�h5���HWo�k}�UP��۫��:�4%݃p�,f�<���nҟ�1-	@ҳ�Hr��l�i�?��]Wў4�XR	,����b�z}Kcx.!������W��el��c`�T��@�J�Ѧnd�L���xr���l�q^����wZ��s<�=�B�8��a�kɱD	(a&�V�^�7l��`0��7Z!�����[E��1p�6*,l����T����8���1b�ݓ��ɛ�%�gʏ�QPp���|�Z=(2�r4.�@��dY:���o�%����-1֮�z��^@O{$�ǰ�y��Fe1aMGѵZ<����A^�ݢY�uӵD��'|ƙ@�:G�Lx����g9"v���4l<yq��`��s�B�?�	�P���3h\謈��^�m�9�v[/p��]�"j-�m�N�����	��s/	�(� ��g佮� �T?͎�:�')30��_�d�]�5�����>�[d[Eq}�Y�#�-bx�2�p�˪��2��l�V4E�x�JHR�^VcD"�y��<��З��(5}^N˧{� 0��wb��BfCd�5�ȝ��ͻ���B���ɍ7�޲A|࣮���5���,��RU/�[��/ξ)�J��{Q��z�zxv�y���΄��PO�)��YA�W��ߌO�����{�n z�-Xi��r�x���kc�E]�U0C�ryP��P��:6�E�)�������A��i`A.�^x+�y����z�pv�)j���B�h	���nh�IU���:t�i��s���ms.�}e�ч�6�z*Eop��|C�wR�E힀F�m�$_�a�|^;TG����!�͈L��}�X] I�D�j�6X�D�x�'��9i �
���Fzzշ!0&�(4�t~S��T�y�MX�ŕLi�3�B��4�)�Nz4
pq��bs��>5��.�9z6-���@u1C�3�:D4�A����
`:J�)Axj�[�����vю��S(�$#�ռ���߻��|f���r�J  �4��7�!�S���g����3P�w'M�MI�ʫ� ��v���v.0b.�<8?RG:���Z��Z(
�٧��Ϣ������GKf��^�	qT�b�a�XJ%��R1�.N������Θ�������:+�
zA�hx�ճł[l��'j:�@��ʓg%n;�K�H�u�.V�>��u��	� �F�n �\8'K��C�˱�Ր��#��*�����
��'���^*ɍ��]��5>B��pe,{A���\�an��3�ӗt���.I!�Ͼo� �B[�B1`��7��l�!�������>,n�`�����M�4����7Τ�1���<���	��LM�ȸ���˗]��:-+sc6�l"�7`��},m���u��Ĭ��8�3]J��ì�>�.�Tg+�rbE߭o��V��Ѽ��U�D,�t=��+�n]����d`������)�m�5G� d�L�47:��l��x~
�D߹}mAa� �̠���&�R�d�OXտu�	�'���2��"j�t��������)X ��1G/H�Fln����$�o3턻'���J˯�q�.Z�[��I8&�xk)�U�U������v�K��d��,��ϴT	&�g�bC�l���m�*�b���w�����������W:�/�f�6��?֖��?݉�VPg�ֱر�SF^� ��X��e��~�rf�]��[�,����w��kM��*)%k��2�����+�����&������Wk}�88gK�IH�5�@'���8V�.�_=O�Ԉ^�5~�.��zb�:%��X��X�6��Ulٙ�wf	�@*��pLc�F��&<�DM�|	n,q�M�.�XF���+�&�puQ�~��C�)�Lh�%�g��;E)pP7e������{�W���` 9�uF�Ĕp&�4�O�wc<���Y��]�9�A�Hmd�P���.���}R���M�>����Np���~�urEE��MB[�я��ϭM
��,Y���"(����_F�� �-E�P?5�ʷj;�OmBi+�j�͉�H�矈3�f��V_����t���T����))�]>���v�M+VR��I��'\3�Z�/��}H��m��l�z	j��f���>�d�_�z��P�o�~��u_�$��p̫���l[B-{_/��0i/,.���aM u�P"� �!!M��� �F{mf`W�#E��EK��m��31��K��|*m�h���zz��J w�:�,�ݍ8A8��d��\T]��N4���F�w����z�փ��(��a��h��s�j���i��,��,,�٧����f�1J�!��/Dh��u�׈�����kȹ�P��,Ir~����i*�=�긗�r_����@GIǉ��.Ta29ԭ�0���ʘ;� ���SN�e���.��xL�u�8�Yg?�������1�d�� ��"��nSs�2�{{�w�������X����Kb���ۑć�=����M ��<�
�y؟�8�u]���r|cHl��')�M�����iB�f����;hkP�S(��!��)�^ �k&s��gTqP��������ɍJ�lۧ��^���T�vp8�����Kz��8����ǳ�n ��br�y{��1�+��9��r��a�<pقG�v>���K��Wu�!.�4dP�Ѿ����c��5�S�9a�����q��޵7.�W���]���M'��)��.�ж��,u�(h���XW�i�:'��v�'� &��j�Kf�@� å�Q�vn�?�jT؈�\ [�貗<%9�`��5!X�]-���e�xN�XVpV?s��g���ya=Nh0��e<Ȑ"�m�* 2[��|ʵ�wC�A����.���H��}��ٛe�6k��R���ba,Q���P��J* YͷY�
�kLT���%��"|P���OӴps�/�('��?0�btU�7מ��.�(��<x)��ɑ���q�w�|a�߃Ɂ�ZϬ.rK��N%��Ro�{���R��kYhcȃ^+���tX�������kQ�(�y#!D%b���"Q]�`ŧ��e����[E���=�]˕��1��B����կsr��BNb���ѿ/ogB����`��#㑟��Y%�-.�P�x"���
@�������]!�m(�C��7"ؑ_'V�oa�����c[[�M�==��a�����Sm�� q���cŖ�������'�e���Ƕ���ƍG����=�_x2�d0kBbĝhg�<M���2��[���'��j0���y�_�9�<��><�Ȩ��E"�ic�vLI�2�e� >�2�'ٛ6D�aM�( ����<?"�ٹ(R�2Ab��,����݊�G|�F����F�3��\����רe�KC����f�^����t�� 7s���X8e鯂;�匧R��N�6.�!T�䯄'Crh����s�:���DYK��M��SԈl0\���$��׻�Ξ&�����P� ��]�A��b&ެǚ�G&�u���32O������2�
,UY��F��R���W��a��#[�rv����ш(�O�*0��|iG�}��0�=�y	TV*�k�1� ��v�Q�L1��tV���]�=wPB2��j�x-���l��ʎe�s�_b�Dt������KCx3���p�yW���:�JL%����[/t�V���&H��8�Wd��W��+QH�NV�0�]��ZË�����)���B.\�ϓ] _z����;K�	�M��Vi��A\�EQyuw����T����9^��Y"6&�CI�
�1S
���:x 8����tl�*��	X��_<s�k=���v��9���|{����łW�[�W��ӛ��N�z�r��Ť���9Ou�����D�@�����lPrs�ù<�",h�wv�s��τ�&���.W��B<�+TQ�xUFn���S N�YhZs\oL;��*2[��䇧�p؆	�5|��-��۶!���%c��Ǌ���|�J���6��!�T�W�Y����z 	$�A��k�u��x��~9D�Q�Zi��p�E���uT���0�Gr2���/ZVҿ��o���=jtPx?��y.F��I� ��!|9���I2.�L���K�_pVx���x�f>fC6�d6�a�"�c�}�8�t~�qL�2��9���ao�2l��:��k�c�6�r׮S�Ƽj���Y4�ᤃ�<��!Y��>�6��K�z6`���7G��0��a�N��m3q���8��"��@n�6t���_��-�歙���eŸ�=���8�0����6�2����i/�SeI����9�zH�:S�@	��=���܃�i\�#�Ф�|���\pt��niF��üqg�ϲ�.g�_�{�e��YFjZK�w�"����.��i$ '�x昣זm�ZV���!�M����"C��O��.��2)�ן����|k��C1
��Y�_@�_zN��l�SR���Tu�Q>���$ԜH?Ί�⭳�l�ǜUd��Xk�I�m�Z�jt�gD�
�I����א���J��-�mkjm�pg��Ch�����)��Xd6Y���L��D/�{��\���@�$� ���@m;@� )�S둢��uN�:qĢ��"c������� Z���%���۽���	KwDMa�-֏�O�����)_��maY 1#���?�8��q���546�2Wr�f>���ڜ��S��h��e��E�<��8.���?�F���O���`i�Ei���؋J����.Z�c�О���1(��x:V��G�g�	�CG��ם^��M�W�U��U�ϊ���ۛϠ�ߨ|[̓���'1���VO�Q���tqy��5�����N+��ə�i���q�)<k��^T��!�DB�]��Xb�R-jML�3���\V�l֮`�WH�5<���i�(�g#ڄ���3\N�����3"d��VL����n����.�U���AS5\D��,+�:�mt� t�G0������Rls8��rX�:�$H��$\|V�e���P�L�N�~��_��+s��߻K<ƶ�0�P%Z.r��N��x{ ��D�XO�Z�pԿ�8+�ā�@t�	^��9?�Q����������9���V��79�e�Z�-v�o��j�5��	K��˟%���@� }�f���H~ �ʡ�~��ce
�z�_	��XM��z疥�b^b��6D`9��b	0 x
�A�%�L]�:;���E�A��#
s�Y�˯��x[h5펄2QA!8{<�����\΄���L	K.�����	��m�(�L��ġ���I�hN�RC*���6���$T"��]�+�t�.�l�T�9h���� 	�m�!�ռ>���7k�e���nyUK� ����k��B�G�ָG{�A�)��IAԼ��x)-���^������ 1Y��!~߼�̠�t��}S5�bo�m��+y��S����=ô�Um"!�����s@��,N���D��vI�mj0S��q ,Q �	�M��_P���cş�o�Iy(%�B�l�m��Ή�_:�&�2L�ʏE7���ؑ�)T?lo#�8n�g�Y��LW|`�jܑz���L!$�t8����	WK���x����A��y��;-��-�K�%Z������D}�?hg����p�� ~.�2��\L��n"�_��8&��{}�E���E���kuD��
���>��.���;l�����hS�*+ӎ/��`�q�4^z䑚��(�H�'T�(�Y�oٴ�l�����8�]�N��uJ����*��+�Ot I�k�i��%H�V�{l6Zf��j5h��si��}K���� .�k	���]�z�T���d���fw��^���0'�f 3
m��~U�Ó�"��)ҁ��tf��F[�23H���쪌8MA����
�����h�4��?<�7�wJ_��|��6� $�L��kII�I_j�Wy�[1ۖ�to�S(��[��$��?��	��M1��Z�s�v�Q'�����}���T���Z��\��`E�-n��h��ڴ�j��Ki�'c��������4i.���5���z{_�GW{�e�p���y��Q�^���x����k�r.~Z�_�R�T�ǌ��^��k9%e\�]^x��_`(�S;ADW��)�N�0��'�~��]?���ٯ����o����Z��G�G�Q�JG:�A�L�|�k,���w�1���NmO�8�u�<UߴٴD�]��������W�Ɏ���E��f.|�=-x��˱H������V<�k�	2���7��j��,�׳���h���5�(UG��oµ��'-�l>Jj �`�ذ -�~�o_����d+�'A��-GQ��wd��/t̖��&�S��N�T���h����t�["tKf����l�a�Jqn}vmܩW�y��jp$�4�|ǵg:k�d�
�$?����e���XrUi�r&jf�i-tK�xKE7A`�D	4��i���T�0q"yq��z��$9H�d�I:	{|8���QCMP�O�c�:����]N��ϝL(����6A�Wj@�3t%YH���^}��͝_I�t�{h$��A�GsW4�5��Q���P�X�b��ԮMbU%�,��	I��^�m?�ڔ���u��E�X
m� ��B�v��C˅������242&�a�$@�0vL/S wf5Nܗ��{~�wQ�7<Z�m�PE�NUQj�Q�a^�,Vjc�Л�"K �#�pJL,ک��?.x�S4'x����C6�]�+��c{���GyF�Le7n�;RZL����8�� ����8'�ㆯ՞���y$h�ɑ�C����y�fy@k�!ӵ��f,ۙU҉�'0}%���t�i��hQ%B����ga~M�/�t��'T�A�dQNK�ò>��8��r �i*�zx\4��"���qB���S��	k���C<[�� &{C �'_�� ĝհ�y%k�6��w��_w�����k�#�]�p�����{B�y邞��3���l=���I��9j�����x���3���F�qӒ�uc_8X�!�2u�Mz����m�e�.��e��~A���[�[��c?(]Y��)"�I�]Ab����~s�a�ig��p6 �$���}���aJ~@���no���?�}&�0��i���,-]L���5�y�*�<d �̒Ǘ~��/��-�+���ȋ����H�`�"=I+dr��*߳�f-'�;��]���N6�5+�b��O�Wp?p���3�g��dS���� ��"gƐ^��}����z���1扒�/��\{3F�S�B�W�:�ڨ��n�JY2�y�����~����{�6/2����Z	��>�y+��FEU��������f�G�v(�i*h�#'���h��Oݺ!�ڄ���I%�T�v���FN�gְy�S�m���!b�|�����:Տr��O�ѿՇ���"��7�+9�ƎcN��V�Z���kB̓n[-���S׎V�C�}�jSG���@!)}�V���λ��L���п���b��4�9�q,��Y�g�*�'�����"���u�$L$�d�A79^rĿ�{�:S^��V3C��\ˌ�x������ң���D=��֊@t�6`���N�=�nSc ��L���n ��k�xW�G9KTjzNMU��ĉ��ˠP!�DѼpr��ݼI���m�@3Bk��ۈ!g)р]z����9�H/xR\�8U
j��[�^V}�?����ܤ����|��'���7'!�<�ƔG�Bi.�tn�ן*;[�+��v�J��#v�B/%�)FLË�3�� ��!���S,*'G��U��0�Gϧ���؜O\�4`�	�D�1.C�p����<���>�#�\��K�xM��a����J/�ī&bK�лr�e�Ч��~��˩-�U<�G|�K���n%������{��R��N�E��H;��4p��� IC�4���
	�,\�����]���o��n�:��&>٩T:�@�r�P���tՙ��?���x�D�`��u�W*��n^�v��ժ�t �A���W?�=�]�h������wH�H��&a�Ȯ3��	 ���''1��{O9ra��-�V�!E��ۢ�o$�yS�mּ��1�#/Xz�#�������U���������(	����J"	��r@�\�6��A�Kdud�Ym�s��Ś�@�;�A���:�a���?� ej�9�S�g�N;|��Y�W`'���o���>��m֖��fJL���b!?�e�μ�Y���K��u6��	���"��.��PX?�Ape�#�1����$q���H�M�]�c$�91���v\1���=�Y�L��'�����}J��M����#����K��M����C���;ଲ�x��H���Vz�wύ�9�!GN^�3]slq'��4~	���Q\p	Ђ^<�x�����m�����ܸ�ڧ�6{��d�7��k�:��V"@��͜�^9�:HE ��\_>^=b�Jb��M<(����<�$���+��%J�$k����?T� ����J"�H�I(끼r@j�Zr(+5^����!�y�v��(I�3�(�M��}c�G�~�����������ꎥ{%yȃ������9\?���1����F�Zf4�䦞���`\���׵������g����������5F�J�����ޏ�L�p���7@�C��G|X"p;��8���%PW�kH��&�ɕ[��dG����nڀ֠��}ա�}�E��.����~��VuDpk��e���n�V�r`w͞5�>[%sdڭp�sLNN����g���y���n�[�]�E��(��p��x����Qd��x6IƂXlbuKɽ���f$X�YbC��[�<i��\�	���-�=qm�h�� �����x	o�1\W����(�v�;%��!%�x�_���3j����������D9]~7���?�] �b���3<4#*�e�����:��5��i���ކ����*�d5��/	�V�v o���ίL��u[���ri�Q���Z2�����&h�+�<����r:���iykT_9�#[��Q�Vh}BY\��VηWdVv³�W����]O]���Wxi�6����e�T�o��u3×�x�@ة��7ȦY�{�S	w��Ñ��`�K�oI	$�{���Z�-�Y�	�a�:����V�^���#����̘�ޠ����Ϧ�[b�G��	ҭ�e�V��2d�� 
}�#=��W@֌��*rl���^���'��߇���c� ����{�i5VIcKvq�&.h�q��𠼇�T��[%�x�D���cc�?��|�<G��� �X҉�"���ǡ0e����p�{ص��`sp�vx��ߞo��i�Щ�JO��Ԩ0��M+����O�Ij�Ήe��h�|Zd���J�������� �)���0�}�
���>m�z �A۳�]�T�N�"�_�`I6I٢eɈ�!Z������F`@������y��'90�ͽ�y�f��2��"�o����Q�������tLx��&쏩�Ϻ+�m���K�t�ݫ��%�\ �7c�I��*UIر�3�)r������}���{=�5�"��Κ���=�7���݈�<v�� ����pI�����X����糿H��ź���]ʪ�J�����4e.�N��J�inX3�K4���[���>*�k&�D���� ~��dlazi��}�FG��y��=eRu�[�Y޿�2�>Q���.}T-j�q����G����D���	��|DO�ϊv4j�Z�£�E�LN��%�>T01����䚔#8:�qN���W�+0c���w��0�{*\q��\����4�����y�7����m��V%ސ�|��,:���1�tt�7G����n���CA�XK-��>��A~ع��z?�(��{�����N�o|�����`o�j�'O�6Cg|0�͊�����7��2��oMi`7�i�B��qj���v�q4Ŭ�!���:��ΐ�gs�X���\��~��<%���O@�w�H��v���T�I��1��ǥ�D�?.�Wi��a���ㆎ_Š@���0ΑG���59���\����r�6mj��^S�0'����*�ʇ�y�J���w��,�}�d�����`��c��lo�LN0_[^�L���p9��]�)�v�U��bf�kz�M�mT��9���:������j�)8�њȤ �є��v��w5[��{��K��[Gs"���]�����R�x�C�?S���B�w�lGy�w���M:���%����ꍽ�l�������a�n7�%\ ���1v�Ƅ���s �02a��X�YH������.2�:�qwXP$fkQ��z��S�P�����#���^9l�7�,)���Ot�7bw�~�MM��@��Ȥh���\��
����[H?��^������v6%b�2�Oj�$,��R��5���Ƴ��>Kd�����ݫ�7�+XsK�J����,�����fC	��#>=ڃ�׳-b���S/��z��<,/WG�c�Ke!�����S&CN����������m�X���`4ő��CȦt ���1�d1�|,>��8\��ø��7ˏ(���mS���@6Mq�ᬁ�	Njg���LI�!3�9����a?hD��Ӝ0�]�0����[<�E��F�����Ɗژ�:�}��"��b���E������H,�t�8�ɗ����	��s���)�\!�(O���e�t:��B������׺��P� F�f�T�]��o��Eɘ
�As��&���г~iќ�ģSe߭���6�� '�n.<g��1�C�$4_���{ia�
���4Y��y���*o-�~XQ�ʒ35�2 Ԇ^ѱ��2�Η�{��K��cA|9��A���t�����;Vv�ӏ�"9ɵD^'���a�~�����%]�y;��F�s�0<p7�ز��ȑ{ɗ9FQ�:���S�⇟����:Hj&`y�ݾӴ+pzSf�?��ɩ��r���������+�}ݺ�g�D��0��Q�/�kT�Gz� �+�Ԙ"������j��OF	�� ���t���C�����`���ς��3�2">E�.���D��q 9���]N�֯εl��%�j(m�}Q��l���&�p��`y�%��L&�	��q��O!�t:r�������4,:�%�
P.l`�_�+�~ה<pnf	�@E�`�8�௎�Ѣq$qX\�~ų��w"����K�u.`߿��>h��UNSp,vh/�|�zL�׻}�@�/�[��35脏:ț\d�r�İG�F�!�]8x�g�'oj<w�:�������"�!qr���ݹ���9����=U�Zmoo����"z|��{۶�}i�C�Dh���'U��d�e��*�O�(����r���k��t����Tg��'���:�@��R�������u����p!9#}��p�Ɛ�C������mxc�A�- �����������2�0}RX���^�EMZ7���5���E��׸!�e���Yux�i�d��{�$�}��e�����P�,�Zf��
��]Ѿ4+�۔a���<5wC�Ռ�.�Θ�5V���7�w6�+�c��<��NzF�0p&
VN,˗�s"jB����c���s��]����O��!E�O��\XE�/�<[}^��+e�k�HV[�d]�є��i��]y�;{*>���,�b���x��VŇ���=���R�ܝ��?-���KW)��!�zlý�&}��SQ�錓#p�ɢ������Ÿ��M�f������8 J!s����/��%��@3^�|>D�5����c�}��;] 㕖Y��d"$��Knx۰r[1ܼ��� �����6�xT�z�a���V�udOO�M:��~����ʨ��٧Q�b������>�ݯ'�_v��"�"dX��UA|����}r����w7�p�)-�'G2�v������vlSpG�@!.e��J�<~g��a��m6����(���`I:?�!
)�9��Y�����D5��j�3u�Y]T0nr�v�X˜�fewV*��c!����=>7,�,��'�Z!������iC�L��h��\v�璋�
�z�X� 	Ŋ��*&�Kd[
����&���J�.�к�]���.z8dA#~�H\?Q,1�K9U���e���Zҽa�4��i��j��-kEC����z�-��a�~����[������q�M�![�>��^��oZ4/��
'�19}&]���k��꺀RU��M"T	j�<ا�ǃC�7��*%�n�eɹ��W�W��Z��I�?���U�DA�L�N̫#G�X:7�ח:ø�5���"���P�S����X�b|���=��A
$�G����];�0��Oi6���iwP �m�N&E+���>� ���!����������ԑ};�a\�o�	���E��V������)�$8�@�(f����������ݣ���'$�;�7�|����+�@�\gj��c_b�v��2�z��
8mɯ�qZ)_��Dl���>��~_Nؗ�r�58�t�I�e:�+�ٛ��,��2fi���P����O��A�h��a
"�f3���-A��<UȔȱ�$�87�nI�߰L��H�4MP;(MW.ᎫVЦ �98���5���eW�^�l;�]���n�ME��h1bY6}�+��K��8r��	���یיR��hb�Ω�|�p>(�����&R
����6����O]��3��H��i���5[���["���[�ɈN���c.]O�oԣ8A`XH'/�L��&J}���̴J��\�/'V���{��r�O�3�"��(!b�m�I��~O�[aQY$s�)3o�,M��-Q_r�|��u�/�
6F�k��R$ �j& �K0�H��&��ÚdSPa@��D�LNӳ����e��˰�Yk=.trC:y��WՅ%+�8���⁤��P�q�{�^��7�����<3���>��+'� `��_��ì��x@)SX��l����%����x�'�#���ݣ��=	�����G�U�7��_\.��w���x7cg{T2�-�b�퉢�Whk�����2��!.�A�*t�Z%m���J����&�(?SҝZF�.��+Dh�8�O�tP�9g��!Op��n�
���W�O�(���@Sx
���jd08.o���P� �]�ս��x��\#ć�I;��sPi�]��pV��7�$�����x���O�����"L�%�>��Q��N�ll:�DT��C{�}k�k[V��`Y�3�_IF0�B��ñX�S
Ι6M�ɰ�$�Z�5��v�w�������w�g���FZ3��Ggy�HN8��ܥ�c�_l��u_z��~d�V�)}��YL?�\  G��w@�$��Q�%��������Y������ǽ�d'�*9S���'Hz2��!���f7������}+�$�A�t�������\i�9($Դo��K�&E,��R��Z�W�?�]�F��gQH�9��:D�iV�d�|��8�;�#^�^0��
��]��pЯw����VY���v�:$�z�Kis�lg����i����|��Z������ꧡY+mBN�̯�U����Y����˧d.�Y���6>P���R������.���P�5K_��/��z/��3%g"j~�9������n�|Ā�� �Nv��gv ��b5��*2���n�:����p��w_�kr�o�s��Mp!���?�ب����������&��A�\��fpvyJ*J<)(�+9k��x�9l����e�Q$�����JQ���s4L�Z��>+���	�G��*�5h���������HƐB�EH�AK�LT�^9�hii���#��8��kG��IP��i����Z�1S�NQ���Z��D~��P�^A���˾�Wn��	7��x,B����a{��?�r�bN��檣llc��v ҳ
��O�ةq����:3C�t��!��N����7��
�k����@�w�E1%��.Q�J�]�b��3a��lZ���ȭzu��=���"�r�Ǉj$�[E�ђ���=L�7JS��O.�l��ć���}��/ 3�x-�icH����(��^�Q9��
RF�X�������TAz_:��h�c���&��JR:��#�"�/䣭l��@����8��F�|�k�^7*���{�C����#��kom������v����Rs,�r�-	�(.�hޡl���dB�敄���/ѭ����f\���R��dFԹ�Z? T]Fڒ��W\���2�JX���S�
���3�cF�������c�w:�3�����N*�eoZ�}-q톨��%���ri�����~}w3=�6,����=1����6�k�҄Hr���i�,�k��T�_�_�BL��}�-H�o��c�C*��R�a�����C�S�͹cL�~��|q�����V����-�*��ƍ��^)$�2��nv3�L+�p��=��_K�a���Uf+?T����F�k̰�k���	���� �����ZX��'���4<6,FInQ υE�tԪ�n�XA%��l*�qvÖ��4�׶%P�ߓ�j�1�(�.	�d�}�D���"h�����0��G�S��?.=q|;#�ǈ{	���t���>��d���a�����ꔗ����Q�|mަz0���U�IM�M}�U1qi+��H���%�֩�͢�Q E�Io�'��1t׃~5�����Hqk���e'A�Ը!K���鞢�"M�q��w�Y��Gj��������	T2��`����G0��k��ᬾ��N�5F��r|]BN�0����TͶr�*3m!�(?����-�r9�s�)�����,��C� s�s�Bا��=r��zMr��>�'��-�8p�P�|Tw3��{�LE�4�f;~�o����C�E��>�}�A��/�l��;���jG�5�7�6Rv7��.U���� F�S6�=`
���Ery���x[����>	�Q����J���&��-��K#�LzԦ~���f��·y�]�޽�z�;I *-�Z����4�HiEWb��CvaE��y����|�"]�&�xy�WH�Ő��@�1������h����_�@�O��c�ϓ� O���ȩiw�H������H���k����z�� �V[t{�dXW����[�L$Z#,����&�,_����M�U	���Gam!T�&��X��)�k��v��\i��dX
�*�xs�D�k�	#�C}������k%uU�5F�-��;Y�����|A��Ԍ_lǴ�w������J ƉQ$�M�2Z۞�j��01[�]����2(C�H�|1V�W�V.��F�E�ݴs�k������2�U�7���@.f�U�R����$�Gc�z~}П6����3�+'�ޣ��0���TAL�E�f6}W�� ����B��"�J�{b����cF�,���l຀8LY�:����h Z��C��,�B���Y$ގH���V��9O��II������~�]�m*�F�8q>�݋�L������u,�p��)���
~F�,�[�|���)�$%�x�]�@*����
���v��n�o�{�׈�W�\ڀԣ,[v��$������A�4�w�v7l*Q4U2+�X]��f/u�fo[Sx���N+O�ݐCU?U��Z��X�"9�!�U%��3������1�#��%�]2�f�_QF���
6�-"�!.	����y��6!͍��5�!�:��L�
��^�R����i��F��8�dϝ1����!�������ݮ�ZsI�
#������aY��dS�����z�P8f#�%�L��|*�{n�!^����,$`���n�@�pkZ]�IK㵨��J�C.7$��s��{�j�󁹶�N��pD����;xL4��.���KV��� l(r���S-�w9��C����ew�j6�U�ޙ�5C�F-��,�7���In�\l4|��8�Ȅ9X��V�����
 �aj=?����n��P���چ�Nx�3�P��`�u�j���Q�,��^��ɼ��/�	�_��ex�$!N�ڙ�����FL�'M�Ÿ��o��-���OX����'i�n�_�k�ݨ#_Ap�/���3����!hp�rb����T��F�ӃG{�K�ר�3ߧ���,��a,�|��;&yZ]��XG�AfǅW؞��DA����-h�Ю��n�/%c�Ku�<�j���~S.aa<���뫆��EX��&��i�8	O��	�ʅ3wQ+C�; ��?�I~s%<ֆ	{���~s���)W��˃Oi����1JB�`Q�G�X{&"�,dBg9�d^"�Jd�R�v��E":�(~�'��Z0>AD] ���帣GP���z2���s��@��z���}։�N\ҿł��$�$z����fN�f�R�#��zG�CQϘTM�����sz�,�]�UON�u���J�Px�uӚ
=_�)>�I�����ne~���k�H��v|8�9XC(�ʉ�L��f1��ک��$�d��_g�!���]�l���C|�3�O�,,iS`㫮pvhT�7��@�9v�1�~��S⥁9���wK�N��{[��&a:M�NO��9��Y�Y�<�B�LB �>��CAK�/�U��y���vr����Bbz3��ær[��6�F/�^���X�G��BXaS���ta9DIG�<�����`۸7���[_�S :��=wM��D�&�B��p�gލj6����?�%���u���c���?Ĝ&��=��E��M�\���S��6��}	!P;��|�jL>(��G�\Z�G	$f���̕R��}濖�
��p�3�@Qv�9J$��ĘsAD�)�N��A��3_��Z�Em'!�u;�a]�D��P��q;�ک�E����Ӥ���pH\�`�Y����Y����JT(;�2�q��4��y,�-�r�?��DZ�A��YpM��onٶSI�Cw��A�
��sW�+*a�ǵhH���\7�ОV�,��=]��0�F�}Y�4`?��� Ϩ��-0������M�t�%��M�!� ��|0-M���s�yU�#�;0���*�}|�<P�������\���}��m�K'R/6�=+I��K+n�q��d�@Tq�3�� t�&�|]��a�E�jl��jj)?N�Ғ�EJ����B�;���L[5�_�]c5-rH��Eӣ�]�n�E�=8yZ��v v�;�d��7�10�<����E5�͚�.C�xs�r���p�B�?F{4��A���m�.m�md�$�Q�D�w��Pcxc@��׍"7���ۼ�s���c�wAÇ��5�Q���撥��ڦ���������-d�߁kzv87�����Xd�D��z��j�G<�(���$�+\��U[09�,��%V��Ѷ�|P_��E����D��z��MW��6
/����\�H��6pU��l��u�1���'��_��=��^J�~�u����oY�Y��4�Wa��lj�! �	�-��0��ϭ�(�g��.�X�E��6#�jE���v�?��-�IߔsP�!��#�x��1����:à�!"�gT��*�:��^��3�7�+���� u1��P�p)-�v�B�t>J�f]�$���KN�>
�͍�/i4N< �����n��t�$�14emw�n����)�B��s�)���c��-W\���D����VC����;F!^���IZ�R�����4�P	Ö�k��8�xS�Q]�������S�ڳ���Gn.+�}u��n{�n�����[�H���r��֪�vC���8 vn~��*�G�i�diI ��"�IO}>�@���@�(��P�ף'=G<[��(�04[�����b������h���1�[&�eq��G���N�DSp��->|m<� �҅Y�v����U�H*L�^��XS�[. з*ă[�F�Q��t��˶C�c�f��!DJ�Iߛ��C���i�"��Y�O�G>` 6�sdz���K���Mgm�B�4�ȟ&G��5���,u ?>}�e�1�#Fuz�x6�"�ύ��tP�g@7X�^�4S���3�#,�Np��V��������pg�=�dS���L�:�i��5 "m���$oU/~1�'js+ғ�V`���V�q9;K[��{?��V�����_-�68G֫9���~O�(ӛ9Y�����b�����cQ�_�-��%يxP؟���tNH�E�o���V�m��'R(��3���"��d(��ׂU:�Ƚ\Ɩ�b��d^������0��UW�am���iU�������4_fd�qb._&n�P�m�h4�#�ٹ�G�6xM����d��tӒ� �.D䪗J}a̄��E�6�.X5O�������l5� n1�����?b?�F%������sҐ����|��x��9!Vءf�%e�����ׁ�+��Z��$W#y�b
q\�<�	Yȳ�ع��s�x�g6�5kv�=�Ѧ&̏��V��*1��b�T�* �W\�h-�E��g+kb�D�Z���D��k��e��p��_�����<��7*ҝn٦WM�B����X����q϶��"�fp�+t1;�ɐ=����4�j@��RI`���u�T�m��N���#.E��~~����<�h ����خ��0��6�m���dZ�g�f�;	�P��6���=Tv��@a��6���g���[����Y>#b�^�ڧ�Ȩ��B�Ѷ�&^<B�Sc'�aUk-��[af�i��LE�5Zq��j#z�>6R���g�q0���"��4#L4�P��;K{�T�^�j_W���$��Ȅ#�����I��+�9�6���ü��Grh�<�/
���AR�Ź�x�Xr&��㹀�7g�}܌ڃP��b��>*��"}��IU:����F (�Aϓ����4(�*W$#�[�9ֆ'"o>�F��B��:��B����Ю}_BV>����~��-�ZE���X���D  ��V	����[��0^�,�`���)�)O�q�4��c���c�ui~����WX��/c}馵Qpd�x'DrU�0ާ���k@uN��5�Jdv�;��ؔt���0�k�OT�wP�2� �o���[\��|2| 	��P�5 ��!���[��;2tm���'���+)>�j8���@�}u��Um2I����n�"�.|I�����
���O�M�u�B�j���Kw�?������n(���m�h��ݣ�@Gǲ��b�;��F�5��]mC�~��+�$
��2(���a���%�"�`B�x��(�����O� Y�y�#")�먁������0 �+��H�QI�~~0�<-��b��o=��1Q��;a�,�,���)�]lh���.�ǚG�5���Ў��~#-j���nH�=�6�����\��s9*=��9������򟤑�7ad���V��Ay9�w�EJв�d��ܷ�A-0��f��:�._p�v��=�DR�r�T+޶��%{u
dc�7�7���;{��(� ��ml?-e'�sM�^b��i��R���$G�'l�	�#;#qw���,:C��K�Z{CV��e�
��a�hUu��%u��&�	�J�l ^�s�G��K`��i��d;C�*cd���y@����{���{���h_�r�ӳ�j�t�I�37�d�xx�2��=�D�9RwB�,���y�"�b��R~�N�ٖ�Y;�m�b�42�{Zw���9�S�'P/��J�p����?�J����Y���P}ۼ���Wv"i_/��h���/d�^��
��{G��N����{J,�G[�C1�J���n=�r�:6��VY�V�8��C��+����{{�z�י�i@�J��ƪ9/�Q� ,$�u*���%x�m[��Q���_�]`w�YBgJ����e{5��4h���DvnӸ�L���ń��/L�8"��ݪW�������(��iΡ��=
�+�4�u_(���p��y ��1ś��y����C�D�0�����G��tbȧ��T��`�/���0�XĬ�=�ۿ���Ɯ�):���M�nCy�@Z��<�D���^H0��٧�@!ޞ��h���u�w�B�Q�k������15Z���J_e\X��)g�>R��ܵ�F��|"��'+n��prfFW)'G�l��q-�B�����d.�����X�bg �[������xf�'P�g8�� ���S6��|�L�'·�kI"wA����E�l<Z̜�#`��=��[]�M�|�����o"��I>�{�����!�W�S��8�U$KӅ{ǥ3���5*�P�/�~%;S.9%gɕLԾ�z��4�RBgZ���I�R7&V�4�8�F��L6�{n6�'q�p��5Z����z�v-W{�4W�	���;�A�m]E��L*�"� Tㄱv����UOr.,]�L�u`�49�*�Lڂ��J$�&��cj�#"��qF�z8�)�l����
��7��p� k�{ɞLd�J��,�ʦS�E�	T2ɆS?O`X���sdf���vf�c�$Of 4�X�;���>CV�+�6�.1��1�>�vk~��٥Lx�O��f�k�U�*_9��ƐjL�g+Q��nZ��r	g�?�H�y#[��U%:#I�w�2��s��Ǹ�H������,;� ���O��@�|�G��#U|����Z
����84�Q#�]Ӎ��� _��pFM�$O�RR�H�0�9�-�)	u�6��LY M?\�P�{����V��j�V8��d�<���U7M���<b�~��/�؁\���b���u�C��cyq*�B��q��7��Ņ�tQ��̆`��}ԈQ�ui�,!`s;��cДzEu��2
�%s��Z5Ԩg��	pNH�D8$��a��b?/�C��9��a�0��}�п��w�}~M�K �i�f���|.=�N��n�Z]l��i���мd^�z8���z���m���Z9��vl�K���Q������>'�hU�/�]`��D��Ċ��"����j	ARϞ�Ѕ��P2#��k�pJ^gE��4���o�Ii;D�(h�U��n)Ȑ��X��=>���)m.nXk��|D+4�f������*���	�ў!	�H<����c�˘�b�����ƆD^���m<r!�?��%Ic\Ϸ������sɚ>���L
�x{L���d��<4��6�uo���Vs�fɈ�POWӇ��N�U���w��܇�j��g0cɆ6�/�eoF��~�P#ʁ���L_���L$�3�_!D��&�Ut�l�@�u(&�G3�DIN<|K��ă�]@�� �U|P6��|�e�W�Č' �\g�����U����Hcp+aÝz^�lg�����SJc88#�`Pw[��e�V1Rδ����
y����0Ya�3��L���L��I�8=c�Ⱦ}�%SdqR���'�X���ڕ��i�u$�uVP���!	�nK�/;���*��5�$0L��
S��D��v�=��@��1�-y@D��9�bv��~�P
xD�pWQ�l�k��������e9��r ���BR���C��բs!��4S�ý~����m���ǉ3�8��Xp����&q_��X]a,�OG�:��
fW���'��v�� ���úY`����)������]N�nm��p�K�ڊ-����z�~_�-��qn�r_�Ⱦ�)�cB�\`����C�ir�2���x�f�S���h����R�HS}��7C�\Bj�|#*�/���l�lVA�ǅ�
~��4����-?[��[F��]k���T[]��M�@+�����?=��{��:�A$��:Ek��_�	{��(�����r���ޅ���$!Go5��� �wk���������	0�"S��^.$����J��qڳ|�H�+y�����a�����<}�F���v_w����zh�ӯ����̄h,��������K�m�\u���8�q�����`����ȧ��>A��62aYM_C���e�F��b��������HG]0�������n����@{Í�Piy˵`�$���UpC��d��5�pW��'Nx[��|�6Oh��o��K�\J(ϲ�H`�9��_Nе�Y���LyXU�UW&���4�nE4�����K��Z�TB5I(RT1�ći�E��c��u؉m�D�����Sۊ(֪����+�D������Erd��6�ڿ~\��bH@�����1u�w384Vr���;�����v� �?�c�8�d�W�I�������P'�}eGp������+���\.���c�L����<�Y'Kz����3Q��;���Ǚ?rv��N��L{^���=4�)��رc�4���3Lt����r��ϚZ].������s~��ƍ���.B��[���-x*w���AOK�B��ڏq�+����?�G5��ѧ�M17SXE����HX��~,��?�l�u�w�a�C��Y�Zc��CB�z3o~�%�s����L�!�����p<TU:\�!�J�(������^Z�R��gQof�a��Sp��*O�j�	�䀋i����~ �A�SĿU�*K�sR�{�,g���/@� �^�gk����=����&�oSV'�1���� W�%�+� �͙��[�׮��*��$�.#�n��ج�v���Id$\Շɩ��3l�OU����0��+'�v�r�Q�����V���ɭV ;UBǪW�3�!-��n�=9�??4�o'�?�T�:��Tȟ���^����$����&]���=�-��,v�^Վ�p��������<|}��Sc>Kϫ
�f�c"�Tu����5x�����дD!L���@�����7��&Mx��1@��nX�ޠ���7���.�I�!�w���0���I�P��N�	�Y���@�Wͩ��u�l�������	���zRrӚ.q]%�q�_
"�s�nCm't7��ua�qּ{Y�b8�)��{��v�ja����b��ކ��$�As�Ck�C��Y]t���^&�����
`��^��K)��{#��0%>%�"8N�(�r�N�e�ı��h�Ά]BRuB��}�>����w��*��R��;�|�m�=fn�_�+��ѥ�g���$��|�t��쿹3��"��H�pL�_�G�����N�D�H�,:{�'�Pn��{M��>�����w�[b�$޺#�����lR���V ���4�V�e31�t��W�&>N��j|.���2�6A�����Š�p+m7{\��xT�0�q5h�8l.�7V|޺�)���)w��jV�;�is.Q���-��Zzxs�U���)[ *7P)��V?�m����#�9�y^'Q�^��6w��\�n��7gdJ������I�i�S�t�;��s21�7���xf}�?��@"8�C�RpD��7è�,]
]���[@9�F�y��[��רS�\�X�	�זndS�n�X�o�-y�p�h.�=���PH���5�3Qل/ep]݆`���=d�N���FMao��Oxy�7y�ݑxǩ�H�{!k2�}���]���{�O�����d�⯬zBQ[\�`KŎ�U(����[�&���O� �Z�2��
{a�Wfv����p�w�J=K���0 ���d�I�x5:@�F	_U>x�	u��I�'[Ɣ��W��{l�Ju�c �I�u~u�<�kI+8��:tq��	aL7������1фCj�2'3@�w�΃���3~T	)-x�V���N����S?�Ρ�UEPsM�|�2���}��d�RO����G�m���#tZ2��lo�{e��UP�K_;�g������H�hy�ʲ�$q�VV�aC�\�en"����m�S��U���i�U�t��7�O��Z����D\�H�%�[J�d&3��L�4k����*
�/�+hxt��6:k�!��ylP!��ab$�)��5E)a�� �pH�h#(y沍C�X2P���6��@W&��t�F6ҟ�q=�!fRHmecc�X��O���8�r��>eg���:b	�|s��On�����Yg��6�֣�KX���p*b���۪dxW�7�M��޹9��'c#��4�ˀTgu5L��	�aq.|��
���}�����R:"��V��Ӹ*s�f���r��1��5��ӵ�Ҫ)�I*mO��B���X,��?0�B��K��z� Z1`�F{�ۯ�����=W3�����Ic�h&����@��螠��vP���l��c�RG�nõ�H�C�\w>�;����T�NeƄZ���Z�N�kQaH���!�`3�܆:�)`���p*/g����4i�z��&�q�Wk��L�`Sd˨���"{��O�����z����*�9��j�lk�؛.@���XO=|��C˚CT���oA��L����E��zh���v̹N��c��tl�l.\��$�?d�i��mK��FF��?����>����wA|��l�s.����)���Et�0?�A.T����Q<��&�@���M ?v�Ġ��;Y!o�#���@P��bv�~��� O��d�>h�|β�Q���8M��$H�Wifo܇ ���h�*�g2�5��������o���QZ�&����3u�����2�8Y�U|G$9٨p��Lx�����X���%�Ҕ�?:��`k�z����]����C���n�.b�\ya��^{wo�u oK�B����;"Ol����!=pG덊�����GGD%?�?�\�	�sO���P���؝8R���r��j�7rbf �H��"uVDTD������}�C^����"ư_����{q�˕�<G��,��F�#�Ǔ����R�
WY�c�&J`ł����`����8�t���ı�h6�g�k�lk�<?���O��^�8��˿�<��v�9Aа[��F��4Yq~�x�� ����0��Z��f��	������GO
=���\+��孳
�v���-���7*\X�J��� ��`"��s�	�g����d��L6����ʅV�Z���_��Ҥ]�WӪ��{sPL�7�IFc��5�T��S=�3Z1��W��Y�������6��|yS�L�,��K���Ut��if��ˋ0�&��]C�_�5�����㢖� �Jg��>���<9�ȅv��
h�}BB7�ࢿ�����k�w<�`�ծ\�IQd��u����|n861P?�"M�O��Y�(R�/f=1�F�����̊�x\���d�N[ ��p���n���.���,R#���Q78���"~SWk$٤`�/ۘ���/��c#񗛼K��i���88�բ	z]���<�lȥ؆��L����3uX�{����n{�Tm��o76t��n��SR���f����G��}b�	F�1�k�%&d'���$c+�e @���h�['����A�A�gGqm��B��/���,�qnr���:ʯ.���"�o��SY��=�?���ʺ��Zs�I9�ar�N��ⱏ<f{����j��}��n�P~�y�G��8�b:�̨�R3��[Iς�>�(4���D9(�\MAcc���Jާ����x�k�?_I×��C���ҹvϒ+��j�ɗ.CVN��o|��d<��[9�������'���٥����&�CM�(���C�D,��3l��W���y��*q,r�&P�v�q����p�At��wi�a`I�6�m*���s����YU�`��:�u�����d~;9�׶�\�5N��خ&c,^�&U=~L�X��P��6Mś)'�6�Ow�k�;NQLe��ah>cW��e�?}̦@SE'�:��Η�qf�x�o���:�9Go��;��r��V��5� #�q�(G<��.���`�������H��;Dݥw�)_�
\�f�e�j�"��`��4���m4��፷�5�4�<�~������W:��Qʫ`R-��!��1�B��U>�oc8�F�PP�PZ0�����q��H"�h&~�RW9�$l�ӰJ~=~�7�Mgd6r��2	�1�Q�e{�7:;]>���PӠ���i�����gŌd��\$�Y�儑��Q��XNJղ!�1���[~$X
ǐIH���e��i�45j+�j��5Z�wڊ������y�V��+6])�膼���34D�ɅN�7�I��Y��xT�_[S�L�*Tʹ����� �f��ʳ� U�wq����Մ�@y�@%�4����$�{�@���7�D�*��P�ܮ�;�p��3R���n�4����b\�_,ů�Z���(�<�15 �'�;1�����C��N,��u@��}ۗl�[��Q�w�n}�<"�h��6�U�3Y���d���G��a�[|�h�z\;�q&k=ˍlt�K-���G�۾��5:UXy�S=�{Hۧ�{�kƁ�s��9W�fb�6;�G�qk�*Ƴ9��R��D��p���w�s�L�m�����4��n)[Hf��M��^+�+,�Ώ�ϯ���:.�5�U��"�c\��[�z@��G�S�H�#� �'��p偉��"�4<;+Y��<���L��*?���ʬ����������I��=>Ǽ�N���go�����	��՝|6}��&ۙ�nK�,����AE�����CG�?����9m��I0`3���yPlk��	7!�nF���L1eϧ�ֻ��V
TO����-��ũz��h*�|AᆏV��7qSP��	��ET]c��U�Z0�Ŝ�Ñ�T���{\8/�.�}�g>���-�\@�	ΥNx��'e(q�*:E������z�ٌ]X����N�P5��B���hqƷ��[��e�P������N������+{�����&5dv�pB^E�,l�	�tvy��G��^�W�����EH���B�D�7��@5T#���=;�Yh���r��ϔ�7���ò�����R�>	����h2,�����&ޫ������4w����]�ў�������.��T+ɠ���xՙh���G�rFz�	M�����:��leS�{Y#�����.���3y�+�#G�:��of{�l�F���)��3��Ɨ�6��E���dG�ќ0�2��|T����Bɟ�]YJ[������G�y�o�T�6����&k�7�3���~�!r=y}.����	~��%`�9�bި0)Aڦ�����*§�b��γ��~�+@��7om�R��n�o��>��5�%E�ؚ6�Xr��6񇪱)c� H����[�d�#+��}� �_m�4�Ck�MX�Z��GoK©Ў-�p��O��홠[dy_��S��=RD@c�i��L gf�ed�W��6CA����$n_БϒF{F��.q��ᬳ�K���+�	1��&)�-���0�f��a�ԋ����N^F]Ʒ
��9��������(���c�$��]|����7�B2[����{[�r���$�vS0_�7lm�*(��u��x�WH�n��ڧ�M)��GÅ9������CJH��KU��e6)��p���'���_V�f�}$��8��?�*U�X��>>1�U.!7{�˸���)Ho�ȞV[GR�z�,�_��{¼�0J���G)n`�g���� 7GI�Ne�<�j`?������[&<��$�LLƛQa&Y�e�$�hG�L�i�2�&ٷ�V�1�� @~V\����Յ�vmG�Z����DD�v��&u�FY�eD�UA'���:b�M�!o�\�>�t�	8`�R�:8gs��ߩa;��9��J�,�(��eȂ2<d>|*����h�#f�eM�H Z5�I3I"���0�A����#]�tTRt����+Z�
�cX�2��i��y��7��p��d���B�����~m�)�X�*_$Ms�q6����AvT��˙����j�2�>lt����m�}��i�$��D�c��ק�g�Ï���D9�a�hq5ϙΘo���Ѽ���/���c��I@Gu������W~t�?� <v�oʞ��Uwe����S��;d�Q��4$���ڿ��m)�Xxz���ݐ\��s�A�J�9�́���0���T�����g�������)���=�xQW�χ�s��۔�w���nq+΅�ٸ������u�:0��jr�9�I߱�);ՠ���bѾ�<��F=��(�(�����>λ��7��ܗ�A��;���f�$��EX�C�o�������Ѧ��677K���Xw�X���ܦn���E«c]H��K�yf�'�u �A�1ݶz_��p��Fn��3OZ��� 'S�M��y����� ��4ܜ�z��i@��h(S�:���Q�؇ӓ�:�z)���V��0[���/�v`{���K�O!�Ax n��l�d�0���?��s#��Y�3���+���{<�
�:{�������
�z��h˓���6[w��Hi�٫BA��o���o�y�*1d�~<�͔98[�������f݆m���8!�hi��'Z#����:��p��F�Ԯh���v&�`T<�Ʊwb暓���_��f�ܶ�y�.�'���sg�b.�����6m��O�?e�#Wo´KP0��`a���)�#��.l��������#�iWDS��x\�d�{�q��|A#na�3;JY 5I'��s���'N�Y�af�#E������1;�*����
+@��x�hf��,����Z-Hj1�)�	��{���ƶ��=TБ�!P�q}�xm� E�6���gv��3~��z�,���H��pn"�E��$��vN��\q����W�����s	�^���C�R��iЁ2i+vQ]���d�K`RI��P��������pS�v��w=�osf��ޛ��� �|����Z;�">��7�v�ԉY6��� \���Ł�;A�-D��&�W.��F>&jƦjg'����8W��o���$�'�^`%�S�@��Ӹ>ص��Q{+�ƀ��RZ��d\���m����i��M��M��B��h]�D�H�?+��*%{~-J�"RqVq���[h��;��?Zgn)��k�����$9��43���N��������B�y���٦�l��/(�j[�Gp�e�$)E�Vs�`	�#�Y	�l�ȕ�T�O�����[�����|Y����;����ge� <m��k�Z�ڬ��p�M���e�����^XC�u���a�y��b�_?�����NQ�w�$ID*11/oG���z����;+��S�7#I>ʏ�)�-���)ԗ����ZH�q�D����.-����5��'�E��Z0<@ \o���bw%0Լ>$oK��f��\�:�!xs@�M:?��;��M}������KXE���{s7�^�s2�]S)!�"����+p�pځ�@��X*��q����v�%��� FM�J�e��ڑ��{��m�3a㷞_�0XrM�U(fw4i�[��B�Y(?g�]+(l:nҷ~�����o~����D-�o9�S�r�v�K��<Ujbr-�<IL4f8=-��b7o7ucEQ�V�ЁMH{Sț�1�R'Ȥn;�#h;c	U���
d궹��5�� �]�Q��t�H�a}x�q������|����F�?�2����ee4���1}��R;���,��U{0�m�h@�Rӑ]�a��U~�!�B��v	��-��?�4�����V'����V@,��I��w�Єl&gqYZ�O�\��'��`��<4�7��F��Xz����Z'�6�P6����U+�|��#yn�A奭��G�<Kw�*���9�Ɂx���r:���^s#������\z�a�?��*�u�����^֠Lb��*�k�������D�ڟ�ڙ�\i�Lh�i�W(�F�
~G"U��l�zs�n�3x:e*�Y���5��"�~,J���E�����*E%yݽ9E��sU%j#��\��;��	�KbCM�w�A,�X��f`@b�E�?ʷ���M�}�!�ݎ�6���I@Z����A���e��X�_y(5�M�1s;Z�
C�{����jٴ��m�6���4ؽ烎	��	�R��f���ԞF����%�i���R0{�GP]��؆����y(�Ys�@Ɂ�Y"#��X��~	�9���y(��I�M��i��a_�p~ΐ�a{�z/����<�ڨ�H�y��7��N��dWI��sz�����$*�y-��fv�����X#���m�̽��[g��D�H���!m�@27^B D~#����m?jW�%ZTB`�>s&�p���0YG���_zY�L~��潌,��F]Ϸ��kCg�y�v��(!��{�5BRU��!8��7�/w0@ȈcYE�A��2�/V��]]�"�E~����*C����p�v��aC[��&[� l�I[���n���ם��g���q�L��q���e��m��"	�� �2fR�5U���;A�t]�m��&iug���<�&�B�,�#�,����!t�G��>�hA�KF� z�fUn�n��i��d�L�ۼ���:C܄@���PC�Q��j�C�V���K�d���_��6Ut�ǬAs	�)J	D�#Fi~+7]��%z�S*x�ﻸޮr�Q,�
�Ժ�e�mޯI~ ����~Z��t��HE��/FQս����G�<W��PL	�����<��N�����h��EǾ���$��Eyz�a��4�H?|�fh�	b�(�� ��d)=F�z�=	�	�L�Y��P�j�׿�h��s	� ������+�H��湧��,���-�}%*�_!�~�+�%�9@v��y0��O��� M�@JZ�Zͱ܌PG9�x��ঠK�FQ�����"�7BwtUT��R���vSp��Р_׉�>���-"�0���ޠ�H�[b�&{qϑ������z�^4������'�(Ո!$��J����)��,�c��3eJ+��c(N���埮�EA��4�g������A��g;4����OP��ͽ�b`$\� P�էJǳXW�V@/���~��ܤ�ֽ�t����a�0�Y3E�A�.3�yuȷ3@�]��R;�UJ�1��۔�m�;�L�=�L�M.kc��x2�*_ �_����!�t��Y&���)Ƽ��+l4;����:�����J�֣K�����f䫸 s.�k�*��B��� n�tf����J���΅��[��o4aP��C���чJ���k�?����&��1�`t�}�Blн#�O�<�- �@�J���rc=�� ���ڭ �\W��Y���f��(U�������O�Q�3�|�6�����1W@gL@HX�����5()`�s��<�5������>B�x���9L��8��r�؍� Mhg��}4'����K�%-� kZ�kw��G��b~T l��f���~p���[Am�ʼb�P��+�L��;�,gx/�&~&�\Ûف�ov��'���Yj�^���a��A�v&���1;�����ŕ��_f;��=p�2K;+�¼?�M�w0VHm ��?Da�R2��e��R����6�g�����I���G�ӮM�]�7�?~�D�ɕͣ���*Ġ�6]��C��7�$� ��<� �����������<��Y�����
S�h���w0?��){�\�ZTJ���rc��V�ʲ�%���(�}@	��?��Ӟnl+����y�̣�$�|Ss���w�U~/4- v5j����p�� ʠ�y���èVLN�t�9��a;9���5ĶgT��g�+���y��/h���_~�6��@���UO�E~�3�Cg,ȵ&�OT��|"�$�V@$�� q�e4��$q�zp(�gtRnk���q@�7"�W+u�T�,�f�T@�w�mf�g���=�rzRY�@�tg��Z���
l�o
1GE�a{]Ia�]�|�E2�� ���D�C����:��5�a�b�M�:#�N�Aɦ����W��5�DQ�:Jm�BZ�VM�j���)��R- !��3�8��)���d�_�좈a��R(�c�p���9����A����'�ԉ+~[�D��9u:cؒ0�q��Y���Ѕ�o�T�m��r���:,���d��/���ރ���[m�¡"���Jsia����DKoRޡ��y%�R���u�X
��Jk蕘�)��,�S���	�c���5��A�~���4��A�_�_�%N�~Y�wW0O��׈�R	!��)� zO~�:�s�ve������'$�|k���M��@��H���U9X��;��D=��h����R�)��G�L�o>,��8�����A�j�,d�&�����!��L*�]�G�X��-B3��D&��%N5��g�[6��|i�hJvS� Z4�Q�|�7��A�/Yn��W�cS�ЗP����(�e����\�N�I�k)U�Qğ��Sj���c��C�g�!=1�
[�)X�>}�sh+�FlT�x�	��Ħ����A��>������F?�ֈ�?��@3�
$�Q���U��EN8�����KF��~��bkQ�����@eI�(�U<�V�0O�{�d@-F��?d��2p^ �LR���܏�Y-Ή�\$ͳt��Pi�	�L�X~4���01��x�KJ^ ���.Cdbp9�����.���r�LӎAk/Y�_��oF�iCp#�� m�Dp9�T�� ���{u�!��w�Z��� y��'�d>���&�g�wV��Z���W�6����E� q=��f� rm#J(���]/�@`�9d����5�$���UR����N��ZRD�e�g���?�C��-��zp�b�?&���#b��'c��ʁB�N��&	q[���wne�&S8T�Z��Th,L�1���'r�R�=-e���<���rgƤ�5��TN�=W8}e�I���3��|lq�-rb���+�[�;����_�OK&�\��7�W�!��W'�� h]�wA?�����.A�>��Ǘė�3i+��"�b�#|HD%nd�ɕ��ީՀ4�R�?,b#��^�i・���z���<�p��WE�Qp�m� )�As������K�\Uej�Dn9�������=h�"��t���Zއ@U�%����u�]�R"��ba��q��wT�H~3j"t�b��v��������A��|{y��'�(��)��s
J�AK�]�2�!��Jq��J*ן��K��k�<ܝŅX�:���#���xvzt���˲��R���4i�>4��8� ��lf�HQ3��'~g��"����g9om�T,��kRTz�Y�:��؀�خ�w�u�&�����1(Qˎ}	�N�R*y��K�+�m2@�#(.c�M�4l�W�B+�kj�[@������RT�P�ELb�=�k����ٺ�4i��+�e�YEF��[���	��b{�*M�]�r��~�[���O�8]0 ��&z!��4�_&//2�߿������7���5����$���$�4oe�q�Q�<�a�,VM��Red�n)�$���_�o̕����~lj������ն�����vY\�"L4Ɯ�f���w��t�)51��/�	u'��h�GIt@��wO?ܨ<�J|@��։6) X!hw��#T�Iƨ-w0<�q)�̦%,8�p�`��%�ȹ�^�#@���6�֔]�A�6c3;Sh��9����$�x�aw��G~���sC͌w�Yz��~�w"d��*���v[���J0����/�uגj	t�f�-�X����H/ag"I��yW�=��/��O�����i���L���dސ�['sv���\��JM�^����}�� �JN�ðu*;3I��4�v�p#���E�W}����l���б*�K��&?�NXr�����X�Cg&Fg���%h��%�9L\}5�\c�n���̵����I�7x��� �`d����%�$_hP㖹4�i3���'j��zn�G;�_0^(�QZ��m�����p�|N��'0����;\CO�r�Qu��#�(T�NQݩ��A�r���H�� ����F�l�u��^/��WK�`�����R=yVB��,�,����T^ƙ38m���q��1d�ДD8��[��~K��=Z5�.L��V��z�+L�%��utǆ̍�����Z��P���#W����6�n�J7�8V�_b��Hg��E�Ca�:�O�3
��6�b��!ۉ���-m��w0�m�=E/k�j�Wt �$��%�D�'�\7p�%n-��fŎ&2Ckĺ&�Y�K�7C�O��,<$����:g�Dr]m@fK��=��父�4CFG��ǫ��M'����;D���·����i^P�kv)�6�gܱ�'e��|��->�Ϸ�P���Mʅ'����Q�+}���*�R����(�b�o̍ƭ�&�q�'������#���3�NVJ8R:(�_Ki՛���蝷K1�+�!
�6��n@�]��p!��CYq�����W��.�ߟN�,�|�4�r�"O�"-��^�U���?nh%��I�6�|`#���ފ�M��H��4��5��Nnn�,����C���G�ε�W��� �iS���R�Qp�"3�>�]v�n�q�O�Q)���۔��݈�?���Sba� |F~z�s|�R�x�?L�I{ ������g�p͛�6�5���E���=�A�U�aP�B�%�7:����M�<��wڸ��<y9",1���8��h����[��4�X�\@[1��a�4L5�f�oYCI�\Y���nI
��pI�M��on��HQ&pH�ʹׁ���n4Qp���j��Ɇ,Xc=�?�v�z�8	�P4�=���0qiqe�xj4��/X(��kD+8D��X5iEb<8�g��y*�&8}Q����4Qj,����D�HF1`�� ��qV��RzR�����¼,L��5�bw$ť!�}�{���sm����i�]$E�<�D'��p,F��h�G���%�I�����F �0�:�rz P ��zr`��Ӹ#c�~�:�*���h͉��_$u#*PDv3����4�w�U1�] �z�N���,֝O 8>��E>��$��ԁ��g�e7T�W�_c�f� �U(	���zl��Bb��g�%��GrƑ��o^�@��ȯ`�pۈ��[M���Z����o�˃K�I��U`�2���e�޾ۑ���mn��wI(�W��S>ry@�A�d}}N�\�Z��%I$��'|T��%�^�8�1��z�T��ӳ!�۟�V!]/�
 ���2:����:�
���f��>1v�f�������F�>�C	V���Ǭ`�T��-8���m�e�(��I�#��v���R~�C��k�mâ���?9�{3��V�������N��T�U!�Y1�@*	�D���E֨k��\0����K�D��.��h���y�"�Γi���'���ܙ�PK�`�/U�.4L]ڴx2���pӇ���8��]�\��NJ�%Hw�5���)ٿ[��}/�ft2��Mi���R������$�s�ˣ���G[�W;4㩠��9S
�QY�ܾ�� Qs�"`}��!�u�eҩ�9������c%VP�tb�f��GO��ճ��<5M7���A�e��$���K��Ӹե��CE>��A� �!T��ATCx'�:7�?�Zb��C$F�ղ5pz�[�;'��O/m�gY�	3P6aCH-H����$��{I�_5�� (�Vz(cyAET��}��<(y�C�-����٬�����I#�����#�ӌ� X[��M���xখ�b��6V�ˋm��x��Uc�Jq�o��fwrR -|�D�w Ux�J��d��o��bP�����	���Ō"S	�ȗ���1u���wG�L.e6�z���O�
���o]jt��
<w��D�hZ�Ȥ��}~�]l8�L�G�Z��w��Ct'��l�7��0ȨO�܈�P�ԩ���Fs���G�v�s� <����࠺�82��nc��R!����*�6��(��
yb%f��O�C�R6�q��r�g΅r5��wL#D8{�[�@��y��$���2��Y�"K��]^v`*{���Td�4���`���;~ :0��7����|���������`������28�����)S[|+���B}�lvY�"F,6jQ1/OH.���z�v��d��c�2t�õ�Q�Q��_�-s���z��	Z�M�"%�&-��m|O����w���k��ƣ?������;�[���$�滧rqL�Dq/��Q�]��x�͸��0���v�W�Ԏh�JJ�BX_q'����e��}hoy�3W��VRFu����.�PLpkt?�Y�w��Y����O�ax��jn42T����M	��1����dp�B�BRc�>UE�R ��E��i��y�nv7]CY��6M�����a;����q���óC#1hH�e-��,��z�,����\�hAh��q��W#�7ǩ�W��ʹ����K�0�Y�Lk}�:����n'܄z�o��-�*����FR!㏲4���ٸ���G�2x��gv�ڪ�����Bv/�B�]Z?p�x��0�P���"ZKg�xv'{?������F��gl.���g���'˃(�aB?a�������v���䇌���ޑjh���qJǔ4 `jO�峽��8FƵ=\�VlҠi�)�m+�N[ 0����?���6�e}$0~6�V>I|a���A����f&��G�Vb�Qu_��N7�2���Ã6�AP:�"9�ZxǴ����K(ʿV�~v�\й�1E�l�=s��܇��PO�$vܡ��\��Rd��I%��b��O� h��/w���F8h�+����G_"�i��BiX�+{?kOٔ6�SUZ���vLj��^զ�"���fW�H��Þ���zNk��B*��Z����x�<��S�X�� k��K~�v�����!�X���	2��h�l�X 1��m��6�na���[��,UܮM.���.�/�+xs��(��Z͌��C��I����4���k��AhR�l�e��x��B!� �͜f����#]�1pa� ���ޤ��6��!&����%R�ȭr�E���$^���Z9a��N Y'c!t2��l�#-fߣ#��<����
�#B�X>q����6�8A⫞}|���R���¾ �d��&��`a�'�AH	~ɶ��d�&�z��w�Fs�=	"�0��+ku׆�r��6]ŢJ������#�$�3���`��:Y0�Ҩ���d�v9�U�kx����Ր��C�"�ϭ��:�#&�����*�q��v|�Nq�n��?!B���`���Nb��{��lhy1�3<q9�F׸��U�j����J�[�
2�=IQ���g��n�i��k���xDV� �gVy�v���{�>��������H�H�`Y=�U_@@��{5C,t�v�D����'��!��3Hs�ĮT�l����V*k�w&�\��@�uY���\"o7��e!���X��/ d�ۿ۞Nkg0��^�?�@�VrQ��s5 E=��1%�IϢ�Գ	�:4�[#b���GA����f��0ܕ�!�@�h`��?}cg�h�7�b)��Mc4��_��ʼ�%>��LΈ5�nkp����J�_g ��с�Yj�]~Ď,j��� ���(u��h��Hot�躩L�`���5�(����yKF��q���Tǭ�������@�uۉ��=��DDQ;�k	I&=dRѕ���,)�k�Ўr�K9"��H��Vn�����?Ks��o1��le�J�Ro�㵝am��<P�C<�8�(���G�ݲ
i���hAo�71���LN^�R.����q�Rϛ������4����ьԬ���O���Ӵ������K`Ww)�O��Qw�IJ'v	r6�X�<׺�%y�]�d����'�`&�4�~Я1{s�W����Ȉ Xh]y̕�[N�L�Yk@�w`(���FE��[N]���J+�B�5ʧ���j�(�Pp#.ډ�/�X�o�Ci`:+ ֗��?׭yL*	�Q1�|���.9��z(O�ą���: q�{�,���m�s^��	�4��wK�S��1
���8bO5�>��+�d.��7�+"k�Y �jd��&`F%�IMX�C�[J���b���la��A������ي9��$������n�-*	� �خ'7�iů�V
���%��wJz�U�Y�6q>ku�<�UO)�-9rn�*�p\�~�ԠBKm�{o	?<Q�A[a=�k�/#��y�X:ݫ�ێ2^�q}����<��Y�Xg�����|��	BL>qT"�b3n)K�ПSmO�ѫ'K�3n�h o��I��;�G���۬�E�b���`$���+n�/B���-dU6�3>�p!�M{���O9	\�֕���87f$��@������ǽ�Y<X)�P8��lA��'���.zh]#����G�r�x�c�#�q\��BX���˄�WN;�?w
�f�n����?�C����]��\�:Vq}�ӧ�(T-) v�u�����u�%�AyN*K!M���%,haƆF�׾؅$��e�-YC��A�x�!^膞���Aɭ��V]0�5)�ߕX��w2/����3,	~ڇq�x�,�J�U���:q\W�m$�r%R�@�@�������N.$l;�袯ntw7�2U��r��AU�$�Pd���g��� oZ�O ���J���I�V�����P��B�� 4�
��HS�Ҭ�J��_�ˋR(9ُנ@צܯ�J(�Mu��	�޳������+E�c 2�O��/�����%p>J�D@��'ϽC����:b
7����=��y�;����,�RN�*#��	?�٤v�1@��"{a�J��������X��m�P�4��Zc5�&�%��f_&�p�-��J�[ȼ�,�ӷ�"
I���PO�;:0](U1B��:A�
��\2��ٲ�m��	��S�Ax;��T�1�j���X����
�,�\�2��s
>�=�ÉI�*! UG�WE��H!3�Q`}/Pl?V��M�7��f�&�!]Y�O�donD�v_��an;bI:T��8;��pr�ΰ�2�����#���`���jD��K<@6�������t��l)��
���{2˦b(�.��?�J��#+
�f�e�j���7҂�˦q���#�4zE�DW�j�T��p|��+�E�J���kR�!*>����B*�;8�!=�����JU(X�I��,,�Pw��7&�Sľ�ԅ1g�k;¢����Pe��W��럦Gc=��?m��EZ��&D2�@p[�Լ��Rn�\�r��P�;�e9����"�x{㠨�S�o�&���R�;�i`�ڑ��U4�ױ�(�^"��C6mmM�-q~��߅��O�d�9���G��֚tZ#�O1]Lr沗�V�tN������l@;��b��St��*���<����h7�);y�����B�G�T������;h��;-|�L�c��184{L
<\�z˩�/�/�G�4��(�����8�'�ڏ����F�%�	��Րḧ́#]j�4	�XQ�~L\��#�?,��dڧ�����62���P6�l�j��k�/b�s���`/Е��Ǻc�Џ^YC��b������)���v�����Y���9w�)�-�$�4+���}���i����r���1E6���5wN`C��pyX��c�♉ʖ�/L�,���T�rzf�fL}�U�v�Ej͌g�/��d<i�C�&M��PzR��*�nM�w3�8�ϒo^6٬?Xf	,=�U���Ӕ�#��,!�� ��,F���lU��\K�%`����Q:�B���ѵ��|֭��a��Z�x,�J4�-)Gv��P��I,v���>7�(�#?5�G'���6��^�h����`��<@0�-/s���g?�����y�U�����x��l1�z@����W���t�"�=�.��؀=D�����/�d%���)�%�Z�HC�� ��H�!E�b�q��t��K���H��L��Ս�E��!E7\E���S6d	6.\7N�	���xi����E���?�Y;��'k�j5�NaHwPe�vKC����y*#k>լI����pn���P�U��H`~�-�p��C���;��>PfSQ�F�?}��/�{� �N��'�)�[Ĥx��zh���a�RT6p	��<N_�wbk��n��ބ	�r&��Ҳ����nq�*�t�9l��h�L���Ӗ�^�W��_e����k��mj��2�ͻ�",O�����L�(�T���N�u�bCrn�B�s�Î��qY��jmz8c�S�5�� ��+������L��r���:B���^;C�ߤ���(�`��!��D.��b���ol[XJ��@��6K]����CGс7���OO~���Բ�4�6��C��m�ܼG�$>~��#Q�#��I]���Y�����0��s��RQ��4d���":H�$�b�Qi#��S�k/? ȳxgk$���Ste�gX���~��UޠO��RO���#_�N�B{��Y���ܗwR�R�'�	��`t���?'߳�xvX�ɠ������l>�UQ�C����RY��bB��Ø�E���
P��uE��lh� �SɆ��a��ѳMZQ#�����&z���go1=�M�hc@R�K��X3^��A#��m~w��F��sE�˳����RC+hw�*<�쑝.��y{��Hmc�?�oh��(�������L��Q��,W�����>|�0v�w���}-�l�k!}�%q8�G���p���I�~�M�Y}�/ӍErܦG�����QL��{���.�л�x�����x �����((��g�7��韻HYI���L����Ax��A��<P�}D�0�R8٨�{n/F]��$����-J��j���8��c�ʵǋ/=A���J���+10�/x��p��hWoBV�����P	vie��)����nMn#��bE�zQ����n�PA�1���fV����=�]頋�/{;D�����))�e��YR���{+z�ؼ�X^ݜ5�^IZA~W��c�GscV�y;-��X�d�P�2�o@�$�F@+�;@RAX;��8�|���9�6݉u���g��b ;�ڦ~��`X�׶i�'a9��r��C2Wź=�A���2��������vv0�����*\C��x�>� ��β����N��ync�G�Gf���+i��Sv�a�3�>�J	�F��M$êb�J*��ƍÈT%�rL��r&D��G�h��W`
��56V����+��"5U�����P��I�6��̼2גo��p����ٗ; �� ����y �Ʈ֙ �2g�KٍaK���6��z@� or����nw��Cf����_U[���I�z��%f�MӠh"�����^��1�j­S��,/�Xe���&�C
)e����_�Q�����87�?��]ϣ�j���Nb����QFQ�y���_5�/^@a�
�>P�1BC4�D|GW���]��A��?�;�S]�of�}�*��8^�!L�=w�Gj�9��Fc�*�:{K\�6m*�l�eu|���&ڗ�D�Z��@�a���&~=2U��q%C����/��]�`��唺�~zG�=��)V�a7��C]k�8�'�MJZX=���}��9��Ҋ�5T���q#��(�ly���'u�#�M�?,�VH�\}�fu�h!,�_#���[1Iԉ*)��ʖ��TZ1�8�R��M����B˝/%���G������A�
���f����i����oY�~I��?�k�U�@���QzWt��d�N2<b��J-mI�����N�x
�(��wQg��*3={θ�y�x7����\���(F":�߸��B٭���s��;|@6�'R����R��vi�,.38����u��أ\:.G��x ��r��,��s�U�x!U������ ��=D�~�f0%O�"�]�W\0{R�\-9]��R:�c�Ʒ)���rb'qX�?�T1�O���nf���"	�M�7]ē��_&��b�3��v��Ο��u�'���H���M�$ �|���� CZ�x��8|ܽ;y��(+(���8!]��|�9n4�Sf�fS��l�-d���G�Q��t'�g /(
1��Ę�J!R�Farf����:��"��Gމ��d�O�e�a���I�h��_�K��%A>Z~u샘�i��D1�n�Y��M1��m&�g�����0#�<�n:�\�_�t�[�/��W��Z�{�qp�����M�� &��H%I�B��+���G\��"1.���ZߏN-���ԲC�_���uO|U��c�XF۲�K�6xɢP�
�c������mE�6Y�;U��žt�8QB�썔�^*��[~����s�w[)�VI�я���u�r�q�t��z2���n$��O,��r3�4|(� �{���K��~�����翺��A���p���i��6��Rx�I/�j#����u
�v�0���Y�/[�Ǧ&k��vﴥ�:� kR�V����WV�
�\1!}�+v3��FJ@�#����q��h����ɪӈ�X�w�*y�yw�=m�H��m`�x[����x���#E[����� �R�P�Rg���� �N�Dq�������%ۺ�a8�:�
���=h�0�����I��eS�hM��y�]�܌�$��%�p�d���i�}*P�d���V�R���HC���Cyqr�Z1�Cy��y�z8<�pJ2=;�9�1Jp�����a(�c��Q�\H��f��E�_�o4֮X�.��,��Һ>T�iU~�۰�| �7����lh�����Wi��䢷6�@ȈDԱH�����泉���&A����m�tA��zC�bt}}{�2/O����F�)�vs��lX�vw�x�-�d��ɶ6P����G(����dd���G�і:�[��@H�L����n}Hp�C.��R�o0����@N��K: ���(�����D�f{�@z��Q6�e��~aa ~�5Q�l"�,WH�F̒��4>�����<*a�T;䏢;Y�T���E	�z���7u�gê1\�:�R�<� �gN��P@CP}�敺�&���3�H��B��V���c��_1E���
^d��q���T�by�⏰-�W+7}�*�A�Y�ڂ`�i[���xoT/�H�����?Sd�A�X�Ђ
�euR��XL ��B׮��s璫��n�[~�W3�!qe ���1xqqBuhlj~���&�T[�
�w5W���cj��c���
����r�c���UA�Hx5�q���C���yz�!n/��-�t�( ��@Ώ�g;���x�:����%~�������I�`�k@%L��叝[7͆v�|�ט�F*��KO�%�|��!'W$�غ��1=���J�ѐ���C�f�"�^@��=lt�̭_���9y�:�o�G�v+Ie"R�RpBK1G������W5����
��,Y/V]l�/3�A,�s=^�v.Q>�)��ZK���6�eK2%T��y�F�u3Q"�ˋ[�B*~N/�x�{�`k���v~��k��~�IE/<�}JJ�]���mg.��P��$�x��)�t?@K]Y&?�6H����ٲ&�������^�[5��~MW�����ݺg�۵Y���n�3�4/9�m0[�mU���=����J� ��r	K��G���<��Ub�G^��`���X��A�:rem�'9|�>��a�4^�Z9`�Xh�G6�D�K�|�ڜU ]]��Z���V��!V��ɲ���s:G��	�Z�af	��d|��	�w۩��`w����;�g���5�����.�M a��ڇ9�s7|���XHI�����E��]��$�A^'H
�ɸx��y���۳�`���DM<��\�wn?`U�D_���#=`^�,t	�T<�^GJ;�w���ʢ�8�*����j"�E��YP?����g�6E�Rl���&�W?��=����(x�Sg��n����-AM���I֜g��7�����H ~0��Ue�sp���'�E >Y�j�P�~ׂ<=Y�i�Dkŭ����8t�+Y�A˽	�[q�����U&��A�"k.lׯ�#���hV���'}�!���(�|�=����n.���V���?w�im3^~�"�?�ٯ1��L+A��b
���rĻE�{r'�O�M������s�F����B���@�󱸊�I�r=��Z�8�5F�Ҋ밪�`�Q��Y߼��dL1���_��5���EI`�����S~�g��:�lM��T�w�ẢY n�+�q��[n����(^�y;�g
�O�����[ް�)�ڔ0�|��
��n�α�~��/�lZ��ξ?��	OƉ,�J��-х����e�9�]K;�Ab������AS�f0�]����e�qC��� N���,%K{�����A��T_�i�|eԘ	���ʠև�؃sM/5
n�
s���"�*-��U;}N�y+t�(��ܧA��D^R��-�?:�kP�J�^ \{anA�g�=O���>|Z	���y#���jes�VZxf�v1�����c���e��U(^w<I�[�N�T;@BS��YT�� ��TЌ���Lh�2UAˀY���F!�'�򈁐*�������V.��gT�������A��{��W�ɬ��i�Vf����B�&�Ο����-f"JOfД/��V�
n2Da�)��2������)�?#�lۢ��9���Ol�L:�Z��P6b����A⣼��DL�!��R�O�W�P��3:�uo}�@\��0�âZ�d�7 i�K6��5�,<(1�L({���{]��&套��?�z�U�ވjnٗ#r�2��+7kG9#`������?TX���ji�&�7uW���e�_��2m�:��y��T���mS3�1���݃O�ݖA�r,����ۦ�����X�n��ӸʩKź�/D��1%)n�K#+�̅���R P���C��g����~E�MmeeZ����y�e[�Xa��_����Tl��Wy��A��j��������>�*�Ǭ�C��֫ Eo�9L3ژ��iszR��-!u%wN*����:����K�F
��c�  ܌&�!��� ��1dPRm`���	hK<�J��6�P����l�\S�M=��e��BFPk!ѵ���Ϸ�S�.=A�v�� ��x"$Qó���to���� �	xsd�*b5���zbL|j{��vǡ]�*`0�� �GYP�<�D��ĉ�g@I�׹*���Ɖ�/ǅ��бx�?ImA�0��^C��U�����M�w�7�27-�I�r8�yd��*<e{~�>_�8.D:�)�/�}W?�:������Kj�f����7�(��x�p��`8����d�͜]Y:��Gd��=���n�%7�-}Q�4��v����o�QH'[T���x���1�Tv��iAr�b��5�p,ݯ�条�c[b�P��V\.�?a K���� zu*|ѽ���h	%�M��F�z�>�������+�[R�辫^�:��n!���1��3�=P�}���	����6Iv1���NU�6Mk��>|F��b���J�S��Ӊo�.	��6�.�Y�vy�DQi�F�{ �?�js'���%�~���	3V>����&�7ӭ=�)C��	�3�sz}���`$���{�`���[u��D��%�M���"�ۭ�O[6�@��E���&\�/	w[� &"�6����sm,1D(�ȇЯL�y�T�l|�u���wh�l�<ۋq���V��.�n��>�6����6G�Qa��&�?Y�S�M�n������������)@S/Xg��4�
!���)Q�*ci3�^4e�z?>�#���R ~�(^7��ɒ�
��Ъ�Ĵa.�}
	I��	�p?G�ɬ�a�����&�^�9��/�_�#�"��Aho�����C�v֙��,"�L!_y
�"
g���v����_
4���y�aǧB&��u������m��7��u{���I�)�2e�m�
Z0���vT�'`���>��Ц�����S�
�E���
�����ͦ�嫣Qd���c�k��w=Ƿ������z�$��̲kc����.��JUgjE�*@Q�~��Kf�%p������!6�B�]a$[d��#���;$��X����δSDӸF�˽7�_��(C��z�c$m��22+����e�3	n%c��.�
�љX�~�M���TD������6&��`���% ��86i�a#i?��,�g����Ώj�,��Y@m�$U!.��k9������m�̼;:"w���i���w�4x�u��)���	�
Cb�,bQ�T�֘�l]D٘j���9�H9���<a��;5%�K���@�� ր%���j�,=m�1`x���䂫ʯrNR�����g1͔���H8�Nn��3g�ױ���y4���&���uN������q}�7˭�H-��r��O�G�2�����+|�����WU��1���`1���a�C��-8�(V�f��)&C�C�T�!� Ӭ�t )��y������=M6s�P[�vȳZz�
&����+	f�ҏJ���J�����d֞��^���ʃj�����$��G;/�w�JYb·�S�?���a�Z[J�2�el�+*!��g�,��f�ve\D��t%�DI���|2��*��h�k�n�P��z�ƪ�p�8��dN��\ՙ2��|��Ȭ�=UWeh]��4ۀi��Ħ�9��j�>Lm2-Ngg|����I�s��o����h@D�	nsWJf���D�� �d�;j�$E���<i��9�s_Ki�u �s�&ʚǛ�]V0l `��eC�5�gD
Dh��O�p߆ս�avI��Z�j��p�"�(�j���Aß�.0�u�"�� Z�.j�k����l۳�"Ns���ŀ�i?���x!#����Y A���m��/�����?�;�}�Mw��g[䞡�d�E��ʑ�7���H�g�C���C�`�V@AO�[H�m���s~L-N��b'OfG�K,Ń�K2��Jŕdj��f���E�v��6�<�F��)��S�k�ԩ���������pS��*~���?B{Sh����e�s���� �	�l˄I
#��\�Tw� �A��bt���W{)�e?��4"R���l#lܪ�a��M��#���ԍ�{u% ��é5pz��'���nx�:Np��7������;��v�~d� �ae������U�W�O�5��)'ݗ�<�nW�۳L&^Ք�~�J�Qr��t)g��j@��m�Z0��gf.��u{�l�9���D���-�u�x(�s�����^�j��?%�K������	�	�������t�|�̢�Q@���8C� �����ɨ�_mAO�-�Bk�%���M�X��=�J������m+H1:��/��S�o�l�5n��V&<l��ˉ��CW��N�ڵ���آ��`��2A�_C�6��m�}p�`iO��QoUjlj�+��Z����,�Z��%ބ,�1Jء�� ���kl%lF�uHm{�D6���S�6�|��&�¥�=�0q1���	�x�u(����{�x�gV$��Y�K��O�4AC���2�+���vneS�� ���˻�O�_�ڶ:&>�P����$��6�mפ�ʏ
��æ݉�)�>�i��	;��$�]��Bl��Cd5�2!�������ˉB���\K�@̵���`�o�������AÓ�\	/f@��s/#���jE�"h��|�򁓿�ޛ�̈���`F#iA����[�RmH��nC����B�H
�M=D)�f/S��<�����:JL���YS��:���9<��?�\�/ɫA���<�`!�����;KLO�О �uz%j�8�H'1�6�|�M�w$�	"�o�M��	=�/�`��ݳ:����N�E�&ɴ��cV�L߂�ӑ�]�8I�����K���0���[���vǬ�P�`s��C��� �˸B˕,"پ�}wm0T2���)�EK�2C�ֿYL�[(�!�*�_�r��	���.��A;�rF��9���f�F��?J,�}��Z��ƪ�u�
����^U�ܟ����q��`�fEM�.��gcZ��!�[��d���O���a�L�O.
&C��"zXL��k���Mf@5^�b�u��4
�n��h�9�	M������_�(�u�u�}!�Jl�Xl.,t�"��1�섣�œE��C#�<�l��!uS���yUX�Ǳ�^�&h�ʞU/L���g�q"/�]�J/@Z6�(N`�Mu�V�^�QI�YnI?0�
�2��S�B�	`��y^q��U���#�6�|���0�`ȉ('E�ήp����ܾ@�}� �ƿ�o���]�+�`�C.:��v׊ ����8�Lı{p�2y�p�ܣ57M��J��T�$Z�T;��ߣ��u��;�mPS`͂� �^�z	�u�:���W0Gx��s۪�`�%37^UZu(a�`�'��?ql��:����kVӟ�:�6"��Z�[J'�D�ƂR߯�[�	:��L��v��<�^����kJ��hg����%���(*ب�mZ���e�2^;q J�B��HT
�C4���_�X�f�B.�,� wn��:�D��-��/)�ƴ��|�9n"��*�kh��_��֗L+��<��~7eq������}`�K�t;���'�ī��_9ٺT�AfJ
pp��"�8g�Ş��tBsSnT��,�_���g�����tA���aRYaX�E��I[��O����L;01i��-<0�'�p�jd�b+;6��p���~�eY���7"uO��S�0�R�oGD���)j�d0�_pON�D���|�e��¼�A�)�WE>0��V��/{�zh�$��I��:䒸�Yټ��\n�iMxAH��㮵��ꔺ����\��PD6a{�ۊu����>�>�=��1�\�`�q,م����̀V��Y��qY��� ;I����G3@���9,�x��=�jw,��V�:�s�� $���{�ͶR���
��U㩄ׄ؄��5��!j[cF��e�U��D�K��N^zE��wSѧڒ�s�si�9P�Rj�k
f�O	5V@��E��}��"y�܎�f\H��NCSz
������3�e�Pt�	�U�mߜ#0$T����@'w,]��d�/���%r�?A��9+��!L� 	szQ�TgWYaY(X-��e�H����j&�f��-I��>��Z���V������j���cSD<�P���f]�P�ҙn۬U��
a��D��)7�|���)7��Ն�$X4K�걡�\�Ҿ��7�)�ڡ�	܎�Ѵ.m֣�Jt妈�w����WʄOs�|���$�J��v"�q�<��a�ǳ�:�u{`���t#&N��R�VYRh��Vz�w�E�5�L_�
;�+�<P� r%����w?ke52�s��U$��H�@�S��O/P)X�;]�{�Jé��͖�P[5� ����J�����{m�~��٤�PwsY�� Y�]Ԍ�r�7ߡxhR��@���:����*E����`�m��
���a���O F4�!1��#%n��dX$��)������㎻���Ee�t�T?/��O�
q�tOR�BT�eT]�k�sw",v;�d��b�`!�훚�D�����L�U��v}c%�<x<�^��#[���(&s4�]�I��r��;�J���!�����)�2�
�}��+�E��+w�r�ȝ��31F��9��0i������_\*�����Z#4cMV\�Q4H�����Q�vA�{��N�3�9�@���Y�_�T��������u�t�.z��m�,q�ئ�d�P@�O��p���1�NI�X�N,��RIv����sϾ}�xoV�/�L�qI�W�)�i����-����F��Y��W�E�{��5.���M��o$�0�+��u:3�wM�O��E�H����ɔ�-�+Pէ��ʕ��ʹ�M9h�٩��D�T�d8ylI�]�tR�%M�&Z̮���?�d5H�A����%HIK�u��O��޸8hʦ�����q;-j MB{fC�d��q��/����K�/���uk[���
�`��u�ݦ�j���>�=�(����<�ة�@D=�`Iا+Z�b�ѱ��a�����.Ld��z^l���5\4
�����n#��/���U5vU�T�Y��N��Is2�8�k�=0`m)v��;`t�#/�@�*��4i?C��OI����?�b�K2E<�ts_0V�E-��I�'L<#����-p�		�C<�r�ln�T{�ڽ��?TO��:i��	�CjD�@���:#�ZR!�Q�&��БO��Ԑ�TY7�^p���.�`~�k��֖ݟS�F1r
�G�o���[Q�����?1*�G�=�=+���Ĥ�n�lAB~N,_ �������aFm�iG)E
=5��݁q��w>gq?T�a�R-5,�t�����~�+���\�t%����U�����a���:tZA�QK�y�-�-�D�-+/�gG��2���;xB8�.��e)���a��뮖�
�Hp��$���ٵ�z_dBt�57��H���Z`ȡ-�1S�=�j���C^��>����F+䚆�|�z��y��[�Lt8�*�W-���i�'�
�/�5ZP�c��t��E�� Ep��.�"'z=A�|&Ƽ�R��^%�mu\h�b����'���؍���nE�B�پ_Z8&�}!2����	 Z�� ��ڇ���������y5�qgHA��O����!�Et��%ϸ��]k�+|��Ȥd����������Q,]���m��i�����||~
�ה]a��c��Bd�%Iu�3ryH������W�h�4���)���iK�
�{<�@i��@�[a�����`����f��4��`�v����qz����;3Y_].�o-nJ����uWpv�`��T[v�ञۻ-� ds)A�G#�\=������xu
y==�T-wp�e|������E�j�����?�ٰuC�4U8�&�jv6��`��V���/(�q@��FrXStlc����E�_������o>������g��)f���u�*�@��Zm�Ua Z�	u(IsD�g�=�P�]�L�h��׷
�-l�(���@<��r]���4�XC�r���pƈe1%ƿ�˷�_s���X'���p��)��+�?�99"KO����@'n�H	1��_M�	��.��t�}��~�UY�^|���(�B�]9O�*7�ym���pJ4Q�����4q
�v� ��:�zt(
�M�M�8ϴ��d�9�����:�.����f�S ���G�8��ko��!�=M���CU�>��a�ė�d^��"f�ʵ ���i�8��B�+�v�W$±���-�Şep'�lm�K�6�I$v&�������)���3T�2q���L� ������e*�ʣ�_��mKe�0�bB����8�:�Y�֫�״�M�с��.|���Yt=�b��ǽ��3y)K�3L��%	�x�����2<\$;�`%��ʟ
}� �����x[�*��ЯR��0༲��_|9o|�Z�+�\�YDa�O�x{Q"�8R� 湘+D��b�b�
���%m��9�cX5�S��7�`��ӊ
�EI��؇��_��	�Ksv�5KW(-�fk�]iJ�v�o�ChD�Y+"s�aL]4L���&fe�6��\'�4#��r��
�̯mJ^J��H�Kl�BR��ܷ:�o�W�̒�����2x/n�률*�60�g/���g�s���.���|�p){�}��0V3��ԯ}�Wnl���c�&�:j��X�_�ꁞ��%�u�iڲٔ����iS[e�Q�t���E�}��\��x�����2�~�S��)l��{hZ�s�qG_��> �|�c�!i>Ǡ�¹����J���&�IX�ZiQ�<hRUb\��e(��aΐ��1��Mb�4T��'�Pϝ�v|���ֳ�?�+w��k��V4�Ӱ	�d��r�gLU~!aΥ*
��X@OBwG��]��n����q<]�Ao�����Ɂ[I�P��*�^~������t��
����;�':v
��+����21�6드P ���q���~t|�)(����^}�G��qk�B3d
�w�Y��(��`�N�F���3���n��$�4uz�'��#�;������5E�dG��n�;)�e��͢���w+��H,&r�A�i�Qq�\<ݸ4烒/�T�z�"�e��������(o��e|<�\����i����s�6�C��4�w�  E�&�5:��l
A�w�h�0�Ft��+;"�W+�G��W��S��q�JذkN�JRI��Χ%c�G==
��\Ld���蕤��o|w^	�1������>͇����Yd���јk��Y`^l��L52m��tsC������+�ʻT�������R�Ϛ�i(��ӆ�n@ԡw@��A)~Ɍ?\���j��h�+���-_��7�آN+�Cu#�5���oP�X,K7[1>��L��0%͏�U�*{�o�H\�=��b!ۑ���3���>�؈��xhl�7��:e����NYt�J�5�w����p{l��e=�q�P]�XK���]O���������tV����e�N�N�F�z}�QnE`ؕF�*�5q�Y���f��W�JT�~I�-��5nq)����i�h���J���qҖ��<ُUI�7ՍM#���3��4��8��D���,2j�*{�5���g�8(������) xŕ��K��r�I@�9���@W���26o�2(��n�gP1��ol��>L��x!�資��[�F�<��>�8�y� ~�C~,���p�+�k�C_�Ko�Y^ߪ���TZt���bVS�s�w�W�����(0�[��{{�����8���:u�(�׺�Z?1�Ӌ<��()�������8ޓ��ᨆ���݆�sz��������!�I����� �ߢ���v��sBjg, �?z}���״8JT	xj~�הm�E��-Ze9`_H�8�% "&0��F��&��Z�����(��P��u�t��ul�	���k���P�â���L�A����؝-@�<���Щ�z~��u�� �3H�H��}���gK��B����Y>[������0����l"U�2n�������~97��4Z3��l����|��&��Ϲ/6r �qx���/�`*���Z"ɴ� |�|g�HC6��{���vP���o"��1���V���D����\�9����&[U3dQ1NZx�"��	A��y���w��
�;�t�d0;��A-T6'c��SH�e���PP�D4�Q����}�]��$*�d�V��Kå���Z_}�L�*-�ʵpeK������Z��m(�bȏ�"y���$�,ʁ�ڻ�}5WLEL����=+5�IE)р�ڊ21�
Y�_DZ,�P�x��.�h�*x�e��e'��4#�����������v�/��
J)�Rn�&���A�FGs��$�;6�}g�ӫ�}���YljsX���ig���EN�
�$��i�(�G�5֍^iTh��N��ȷ�k��@���Qؤ�r�J���>�����R�x<��$!�B�>��bOH��Pp���7p B� i��.����.-�@�|�$c�s`�X?�轩h�1�,��oV�����N�����u����,���G��	*NVUǶD�Nw���Ռ_.�Sܒßc8^x��5����C�$�-�Bu0�����^������<(EohT�[�v���`�h"�ݳ%Ş�C`*!mӒ�(�9�;E��]�ǣ�`�'�q�����A|�mY��n��-Y�_x�Yx�s19x>��"Tr��Zv��t	��#F}�?)l��i�~��U�OK~|]n��,�_w<Ј�]e^	8+�����M���'OV�H�_��Ƞj�r��zMz7�ز�� [�#�XE����o9�i:���Y������`#>�<	��˟Ԓ�+ӧ?kQ���zc�vc����2����;�"�Qv�J�':�0j;wQ=EKt��������B�Ɉ����C��� ���j�[B�T��s��:z��*��,�`�E�4d �=�D��0�0����頿�Jv4cT#f�;�k�(��N�¯�<dY���h��@�
�*j�f�8jO��NfAh7a�gt���j�+�S�߾h�� ;�Fdԑޒ�u�j~S&��]��Z˸����kl��e�D�`$Iˑ�l�o�x��(6��g�� Ғ�##D���c<OX��_�&�;�gjp�7��=M;l���������H�
�3U�lt��Y�s3-)3�4��64�l.�����N���5+H	*B	�]J0����EX�ʡ�=�*o�p,�N��-�G��X=�1���i"�k8�$��M���#:H)�]�E��C��rQLC,��wS_�5}��N�Z�. �n������ƛ�O�4���C�7h��k�B-F	�܅|�{��<�G�ܛo�r�n�A���)��([X�-a��T7Uu�Ƥ��渋�r7���L��m��TPr����5u��3���^�:�7����)��ޠF�ڬZ�]G\����zu���o����h�R���)G3���"��!���^�D������Ӗu�.+E�4�x`�k��4�s�ؠ�Q�Bw��Qvhu�Ǔ�!�%��\l��M�V(��@���!����y@�E8U���1��q$����οL�]��qi�������� �u�0�x�5۟V�&{X�R�=��'?�ڢ���{Q��K��#%�<�ϯY}N�3��Ģ��e���ɜ`��ĐIY�Y�Qq���Y����/d��7@._$Ŝ���`��k��% ��t�X�(��d�|}��Z��l\��W�z�6{Ճ��!��Nęܕ��h�n�9.��Z��*�?u;�vI���@%[N�l���/7�) �'X9�F�H�R�,ʵ7� z��#�S�g�G���S��w~�^�Q��E�ׯ�ͅ{��&&���m�Riˠq�Ң`K���ǔ��I����GPV+G翀��.��8Ѹ�|�+���)fP���%T��?ӱ�66u^���Fxc�_���t���q[��/?�:e��{R���;�]�4Qw5��j��Wg��rB���%ᑇc�s������z5�x� �B+�1|%��p���8�'lip�l6O 7�P^�|�`0V@JA�R��Q>4��W�.��`�ja�xf��T=�X	�_\�C'��;넵NO�1�|�t�b߮z�z��xE�J�����$"�l<��/ۥ�cY��HߖQ�ň���7��Ygm�����]���X}Y*u���@�Ͱ����Po'i�2�~M�(Qr�:��t�	z�J^�����q��½�9��Z��'�gSk�u r�Ex�ve�%5���K�Ե�b7���1fړ���B���F����Fg�x$�s�7�Ǣ���\�D�WSþ���\m�
�Q}�g���t�C�#���'SOIk����IZ��l>�#,aS�.���i�cL=ڗe�X�6kpT802�Y���v�{ZE�r��>}�Z.��}��tn�F�u���u��a� ���!"��!d�HD<�����I�k|2M�߉zjJϚ�H8�]daM~uD�����ֈ�q�;Q��w��!]?~�M�/��'$y��	���3�F���ҭIr���aa�0��tW��{)KCC�X/]���H��سU�`���(��?�_Vl�<Gi�G��x{�&�H���m�����Z %Ƹ��l�g�&�X��/�c�_��o_%�����T��;����N��2�a�0�H�c7��23>��"��_���/���)�q��Q���!�4���+��5�3Wu6Z��{#�}:���B�U�ý:%{�K�����Xm�����vlb�����j�r[���{�;�Lc�C<�>B��]����/���og�@̔�뎌�?��^�a4���-�*h��#U|-+�ޢ��V��O�>m��P
�^��X����������7�Ws��o�9��M�]��h�{N����b坩E��N�����q�I>z��[�0�t���Nc!����2���ʙd6wPz�sr��BH�g��f������	F$����#�^w�b/NZ�Znc�"ƀ��~�H�UH<b�*�i{~A[�&P�ɼL��7��5��]��>cΎ[�8!�ؼ|9��e^طT�l�M3T�<V�OH0�\��/�E����T�������Y�Ve�!�z8�������Ays8ߊ��6kQL��X����N���aW��f�9���,��D��,�c*z���1���	�Ӑqz�w��S�P��Ϻ�z��R����3V&�������{�(�s��p,7�bQ����s��'��N�����?߶��3�O��l���|��FD�lS/N+,[�Е[�fJ�]�H�ߵ�~T�6�l�2gO�ɠ8����	�}�G�S��@` h�-8
hX�Z���;:��8F���hY�<&u��S���)�
t3��	X����Rj\�AYe��6�X��Q�$7�!���:�ͨ7Y	p�y�b%�e�������'.�}�rQvGOTĽ������ܹɛ�?xm�Fv�"���mr��(���'�8���j�͗�;9�p����n��(r�;�^���ٱ�K'T�J?�
B��oe(��9I��J��gƵ�'����Om��ڐ�.�O�'Nu�έ9�{y��Pq`�Nk˵Y���)����x��`o3ո	j=�GJ���<�3��ݔ}"����m�C��:�2K�(�����Vd��i"S����ㅧ0~u}!z�ɏ������p���"iT��2�P�1ד��J͗w���Ҫ#񍢷�A���I�\3[���J�]��Vm2������#�����ޗ�o�G�Ax���Ѓ�Z���TӉ����J݊)��Q�:����3���D����d4/�j�65����[H��oğ�JځtR`���>a|��3��㧽�s�Q5׷�x�̶�Ίܼ)�, m����v�vV�H*��[,��I���:���M�^�$�]ql�;y��+`�k��	S@�r�,+D�e�$�߱`u���Eu5�!i���Z*RI)h&�b�� ����I��I �WV���$(x*��BڦE�tp{aF�"������߉3�k��x�wg�N"-/y�OxL�����%�VC2J}�r�K����Obє�������O7 ��(54��� e­}\�B�pQ}˵�v�ˉ������#���3F"�$:��`8��
���Z\E7���8���ƊΜ�{��]�+�y1H<�޹	78��m�E�}T~�=����Ö%E����4�^���K��1���䦫�*��,�<�BA!u@��:i@D$k%[�J��wC�Q����$:a�b���w�M���� p��~��D 6g�@)+���%G��E#��tc������U&#L�ʵ8m��S"ޏI�����n�����~������0K���H24 @���}�s�p)�̱�`1s,1�7���c�'F>�!h�5��#)���b������
+��y��}��Y��}@Qz���	t��C �;6S�j�ǣ3ճE
�8��q~�k$h�T�%��K����0�E��hJ8�iKr��]��r1AM��:
����K,���|9ZpXX��=�w���o�gI�bjq��̐*�G_a���P��{���ݪR��fA`dy����'5���x�U:߯Z>�#ΐ�l�ф$f}�5Ju�N
-�=姉"�rb�>��<� ���u2�3�m�����0ª�؜�t��}X7d�xb��hZ�h�+���¡}%n�O�!�H�*i\�ۺ� x�����kwU��?O��R��>7�`��Ny�%u�߽���Eh-
�p�'�����k}���`f9��_�@���&��/�d^hp�J��ַQY}E�a�ޟ�(��R4QW�	C�ml��[!�m�A���k�p\W1狢=�i��
�cypS^@�IG�W#1�R��1Z�Rޛt!�������vV�G���C~Ⱦ������H��S���Zjʐ��a�/�-�q+�Y�|��I�Kߴ�k�DXh> ���8Z'�����y��xZ����(K��7�a�����T�&�RM?є����$�P���)�߀���6хە����H<N'�&%0�CL��0�	���)��Qk��u����;\B1��@岎�ⲣb��?���a����5������P�3��e���ʔ��<}���(�[lӞ5ƪ�C|����w�~�3� f2qK뜃.9��D���5��8ٝ[$~�yP�%�U��r�P'*��Ff#E�ߌ�a53�~j�
+���	Z�.<1��`�������U� ��ı��Gri�H������:���>�e��]ګ�����h�^�0��JtX�	vQ�j�n{�I>�����<��%z��$ﲍ_2/bD�(�~;62]֫hTQqg�!� ꇘ�j!둻K�@@����(��Ss�돷gr��
�+v_$�"���lW]�m�܈-�#c"#��7I�I���ek%a��{-7h�R�(l<��_B-�c���{�W�5��'�z6�[�E&$b֢�v�aȸX�Fd�.��@�.�"�,.��z#��u%�{v�^�s
Qݑ�t]ڗ��=�� /R��"ק1YS�o/�s�{x���M���K��K��B֡��q�VJ��$��L��i�u�:�grE�i����L��r��3�q�3�z�eo.U[X��5�+� ���r����Y�\j�j�L1˛;��j�:�vyގS�Dd������(�	�:l��Bيk]�������K25���ÍG>̟za)mf�J��j]��jذ�����#9h�>~����_��6�]x}�,��/�.�H9~~J��w-��î�v�R zy�5[����I�	 <�@,o�i!F�X�{���r��C����#S�>��"�����dñ�O�l��z�HI� ���t�"�𩣼��
 n�� ~�EV�C.[٫����=%\Ad�å��	���}:����y��5>��7:ǁZi���<3 �����r�g��r�̰3���<YNWSNW"�/(�Ϡ	{S5�[�`,lwY_
��;�n(|ز����X#�C�Ðp&�3!1e�J���i�V���ىq���i#&{�9���2���)cs~R�C��z�}�Dz��(�&*�N룇�����8�Ԗ��q�5���Z�s�wބ���|~W��iI��lK��(@8O���rg��Ǻ���1[��S�T�(���wM���1#v)'3g����kMգ�����F&�Z�	�r'�5���a�RJ�R7��V�\]�����R�-e�H��̵��2�Io�q?r��Vgˑlӏ�
��po�'��[��Kjbq�"��yF����dQ�c�b������	�h'�<n㱕�F�g�� 	��0�`�MH�瘬]m=���	�n! �o[��%2��j+;��E��3�Y�N��K�JЃ���p?D9�ps�gŵ����l��%
�e�'��v��q؃�q�o?�.m�B���$b��eW�sɹ��3���{�xQJ9�j�ٯ��s�|�����m�#�}Ywm�����g�:�w�x����<Q=A�b��k�\h���x"֝U ~���w7#�A5thCE�{Z>��_����)t����'OH��D����s����ƵWJ�+D�ZфE�F�c�����Ly�j&�+��P(�z�bu�{�6\���v�`�j�4�c�`���>L|��@Mª)i
��|ݪ��W�k�お�����M��_&��؎�gC^����X�w��0yr;�m��U�@�����ipV�dq�g�x�K�Vc�O�a�n�*��%/n(�E����.����l��� �a�ؔXXS����&6^��|AAMx�򕰅LwB,��l����^��x�Y$H5o�-�$ك����S�۔v����cHi�g�-)符�K�;�p�9�g�CS�_2�]�<���r�;wp^���zt�7\�]�&&�7c�?��D���Z�7>���{6D�4�V�<Z�:bӾ�ʶ4J�L�}7�
��4�ҡ�{������y�V�[�X��J�>E�a����u}i�V#C��T7�^�69�7�Y ��/�7����+P���0(�_���CK�3����X�lrD�`�!��w��ʫ��.R�U�K�������{ܓ�ǒ$Ǯ)D݇A1�ØF�x*F�yE& ��xJ,=��/=�'��PG�(��4�
Z5j���s��0��D�Q�G7���?pT?���)�s%�R��X��O4I|��i^�_
�F��X�g'@�Ј'�cw��O��!A��r���@���D�Ԧr}u��=�$�A���{�ՅD�������r�S?�����{�7�Rﵽh�|'��(�C����D���\��!�T����Q�0Ϯ��zE�b��:U����6R���~����(��i�?��-�_��*"�v�vl�y"����e Hm�%������R�h�UO��:��!�6C*F�q�N@6[���U|��ØBt&�!��s$G�49ڴ���{���M)�];Hk��1�U����nm��s��F�����XKR�3��b3���LN�m_[�\/>� ��A�:=����(�A|y����*+�~�*�w������HH�����6R֣)]�[B�otk�&Q����5��b �V&w߇�^'7*dˌk�o6�	�ZC
#�>#f�)�Ģ%����j�6[|^�95r�E�O+��?H�7��8v��P��(�p�A�����|��ϱ��)��s$��Yv��^����.@N�>uP 3}*�ȯ@�A��L����3�h��H���j�Z�2gR��H�����0� ��Zw�3aP$D���;���0�<��@+�q�H�g��(�<�ŅTc�'.�i�^>Qb���s{h ��XqKv�̚S���O��.��1H�����7nw%�<�y{���'ͧv���*�Yce'N�?��?*���/,kctw�d����[H0�1n6k�(;���A�H�RFQȼ>��!��\�P�)i𓱪g��7q<=Vڲ�V�-Z��]$���@}�~�%V
��{�����{�K�?6<5�ԗJ�UT��;V�	&j�[�|���]ŀ2\�ۙJ�������P!}P���Xρq��Ӡ1�ڴ��*�5���������=,KJ����z)��Y?'�����Fz-���b��bp��.�L$�2���e�,!�1�4�4�����&x��)�AcHj�Y^�Y*�p�U-��WO�8�k��#c[LXs�72�zg���o��@�S�uko�o5z������1wx�èa��Pw��U��u��F���v����CZ%�E�����b肠��co��@�Ģx��{Y�c[�:����?Hݡ��n�kc�����F[3_`XtN]�1Ӯ6fٔVR@���@����*;`�,{�
G�&
o�8��m���ly�F��C�z]��Jh�w[���d�߯fʗM�h�ڼ��\�aVr�-kӤ���VM�|��&{̖gkMm��(��j���,@W�-H�3�����3��S� ��!)���W��r5����=#U8�z�T��|i�7j�B��:�k��J/��Z�tF�*`��<�=)4} �t�X�6}!��B\M�����N��h�.[�y�H��!�iَX��;]`cN#cd,z��;����BE����`2TmIg��TG�����Q�1��-�3���Ϯ��3~,��H��S�Kw�1D}���C6p<J�����u�[ݱ3##�:�̗��x�@�T���2��6P� �G��Ų�ި��D>T��!��z�������XUs�A��{��	#��aL$%�H^G�>$nUI*�Ro��v����#���@)Yp<�0g����yV�3��Pk�'=f�	��Q��<��,0MrT1^oOB�j�����ѫ��EMkW��Q�c!� K�)��Po�-�����c�P�L=�%�H>����5~�AhB�_�p���M5�;�"�$��O֗l�r�c��d��á'֙QK��̿��&K����ߑ��o
��!Jpn[�j~vY��e�4FW�C
�����"jε��`��SR�gSUzs�8��� Ff-��1��Y��y�ҩhmu��0_O�XF9Ǿ�@�9԰����ś��H�YqE+a�%@S������gt�OS1&��qBC�q�A��{s� w����Q�D��x��[�w7����CLdZ�W��E�L1�����_��Z�$�� w�m�9ې�g��M� �t�t�"�u�Nߟ�V����/�1�y_D8��Œ����o�),c˲R�^
cQ����R#{�݄����}	�H����t>�8˧�sG0�z�whR��\`�&f�>Y/Q!���e��dIl~�W!�2���}�O��ῃD���O���?�y�A����?&�آ2Ch��6+�d�*�K�HJ���]�Y?xUQhE�hۦn�J	ԇl��CI�����w\��Oz�$���\L��-�1�ޒu/ǧF(���1�݀=���-w��,/���h8rD8��Ѹ/�%���E��ٹ��M��CxhM�!o�ty�H=�x��p%�!�	{岥��e�dٵ��\ �`��w������UM��!����-|'�n	��	�' 6m�_��kc�چ�5`�"��C���]��M��;���Dٲ�F���b�UN��t~�� ��!�!�Ng����ûY�T,	���]B����ކ�y�+Eg�3��j]����>�H��1�u�J��$��Je���|����0tE��}ҡ����:M��ɨ�D�?-���z�ˉ��k�*�O&t�>�5�?��o�&��3襉+�9�@���*V�vx__�M�v�G����5��W�L�@y�0�(�9v�1)H�p ��5�i�O+KET�
���VV��Z��?'����� |�U"L���_uk-4���@��XG�#��,�w�yϚ�S4GY��wb8�V�`e�4��6<�� |�H�8���|-q� dK� X\.�Jʬ�?��	G��I�?�Fza^���ӡ���LH V#��/(>>g�)*3>���n�+�(?��� �c�)���`������B�>���Le����i������`�?F���=" ������-��m������F�����[�K�t�(ċ�y/��BKfkV֚~��dB���҈�BY7c�p-B�5��T��6ѕ�OE�W�T�U��C>�tq�q���o����I�0T�����"�,�GmS�0h;$�ԉxQ4X��0�=#	sȕM�"l`�fLqŋO(a4m����c��A��ۤ��k������B93����]�$���w�~l��Ϝ�O!�]�f>���Z�1<M�m����܏|��h�K��+:��>L�@�* ���T����
�T�NIb��<���&�.ﯗ1�@7�a�P�����u�q-�)�u�D� ��t��5�+�ו��T���!:{�X�������D���C���[}é�gF�<�7�vW�|'Y]R;�Z�z8�p#�m�Qj��.ݭ��+H̯���g�*Az>��<�%9�g����Z�#�i�S��B2K~!�A���;1Od��P��gz��2���"	��(�;����DX��X_oS�TZpf&�wJ��&��hHּ%��8
1�[�V�ʸ�;":~���.T��H����k���f4Y�OJ��R:���</4�<��$�܉��ӧ BL�a�������6
��tZws����E�
4��,0��.���	���(��tp�7���e����Hr�e�}b)p����̍D�Scܾ�,eH�zڈK��s���\���)���7p:�$�;�J^���>�X˟��
��k�DU1�%���5�hP�,*��g{��	��[���Iܘy۳���:>1�Q!�I����6$i�����D.��b$�h��q*��#��%`�_+���ƒB1L������o��/����q��>��S�=���L��J���W��v�J�!\���Fqа^%���&�.�Ɪ��M�8�Sv�K� +���|�3m��T4O�$$}.����Y适�Zt����gq{G&�^k@�k��k�9���Ǜ��lp��d�z E{����
+/���ʃW6P{8V:-�[�R�R�-3ɶ��������0��M^���4�s�n���#������UkJ�8%*PC��� R�U�2��G���Ϊhv�h�w�c:ˬ4�8�IL�|���Ax�&����3(�E�S4'3�d�n��l	�r���XsY�ч�D�Cx�_wZ]ǧNo���Ň'�|0@}xdS�q����5�;�/��ԾW@��C¾l�Z��h�ԗ���O�I�2;��<*��YQ��z`?�]��7i7���v�ke��Mr�/���q<����^g�ׁ�cή@\�5��T����6���a��ߛ�(rOm�Y��loM�2�n�����\� ���m^��2��)�6��^tx�2��w:2)����~ `N,_����x��]����
l���VĿAkjˇ�2�(_	�q���"9_U*�$U���=�$rv��/1�ӊZ�6H|ܽ��O�y�:�z��f�F� `W��V�ZfU�iS5��ZEo���`��]��0DG���/�|�_0���Ư�Z%=�T�5y���7����>�b6�C+��������O�ky �@_t9i �WX��߲���	<P��ې�ʒ��d��&��a:Bp\�OsF����]�7 }��bk���d��Es>1�Ň�DA5"������#P��q��b��n<ebcs��0w��8�_	�۴%���OwZ9�0����MK6 �bޢ��Ab}`Қ�t�����S��S��k`��X>�
����֐+��?;t�Oe�ժ�U��cXr�넂���`���}����^�E?����b0�;[jjӳ��<��)Pz:��(����rOpY�v]��\���UT<�rIn��	���u�E�/��iO�R�Uv�0n��`K̒�p<��/�5����HP�9.c���ߔ*]�5X�����ͫ|�݉]%:���M;"9ۛ�'~?����:ٮK�W�c���d/�~��$��U_�b��,�<"��Tw��̕Ș�,�ṵ��|�5U�)� ��5����;j�d�G�T�e�p�:5$X�m�HóE��7��9Pn`����\��T!zQ{Xf�ܬ��FID�Of�Psd�VO�0L�Aη�>��\��ķ�==�|��bQA������������Q�0�ʙh[a�;�	U���;���)�Q��g�g#��9�Y2����^Û��b��Q�x�$��Ϡ��+�B
��P3Ĩ�\��U��
�6% t��+����[��WI�M���AV:tն���2n���'V'&qT-K3�/'�ԑ�6w��k��b�u>KB=���YhIQ��氧�%a�n�j����,F���:��ܦ�\;WPt��뽌q0�y�[��Lb�>�j.�bᦘof��>X�R��>ƧO�U�uu<���3�b�i�kk%�s�<,�D~��G$���Cj=�Lg���IH;/9L��e.y=�w����mk�[0�#J+*ź�1f*^�w��8�6�d�`�EI�@)M�j��Zo��G$hcΗy�a�W&%���pv5���Y�<H��EҎ�jC�Y9���`/X���ANݟx��=�S\a�4>�#^��:j£��������+_�^~��L��=��Md\���pkf4�Ѝ.��Y~RΌ+p�vsK��y�D,f,L*!|n&v_mN�'�p\	�T�r)
Qf��<ىwK�a�K�����Z(]��*p��N6�xE=��l)�r@�}���k\�([a>��$�-܊<U��!��"7��r��6U�6$�ٟz�"Aw~�|�\e�?{Xk�_)
)h�|`Wm������U�P?Z��A"m�LjQ�"(<=j#B<��s��Rm73,�%k�)���ǝ��f��Qx�#���g~�My� ����L���
\!��Lcd�Xb��-�E�"�H�t�C���ؠ���q�����2���Y����T�{۩����{G�9Ɍ��!m�ߠ�V\�? X-�X���ם��9Bj~�ym-����^M+XK��ݹ�H@�ц�O�:_U������*Ь��t�<���Yۅ�����r{&K�*h��0�����265�N��8g>�2!��T5�7RT�>t��n�η:���0�E��5��
יo}٧�vC��e���*=���#z(�ʐ� ��a?T�53��7����S̜��Z����O�z�9������>'ϼ����s5��|}d=�䉌�$G�xS~®=R|�?��7�( �Op=W ���*�0�=���@�T*p��ޒ�ݶ��(7,�V�0����Qs�=Gy�"�͏�혟��� �H���ya3�ňSw6)�[�. u��u�堒�WQN�R<�2^X� 4�;�����ot"�
�~�!Vy�M1_Q[l����M'�{���3ꆸd�l	�ۋ@E�fGJ�4 �o���>l�\ϓF;�{"ǲ�u�ζ �B�?�4s&�~~U	�jY\�xt���� Z����L@��J�QE�ծb��(���q.�EU<�	�aD�z;K5,�*96�g�;g���z���v���xQ"dp�,D�9��gg�H����m��{���1u�Cǟf��}��1�x;��e�d4�PN�祄J�Z_�.<+�ծ[�ڜ���1�en/��S���/M�edרŗ,?�@��8	2�|�~4�G�y�T��yw�6$t6�g�H-�9SHN���n }z�ϷNsꒆh�N� ?/2��|�*YU�Is6u>�h�*ʒ>�������?d�Ƭy�b˭�)�A��)f�H�!w�A���T'P�\F8�З��d���
Ց:�=�<|U�c�4uCGAl�2�o�W35�zb�L�AB��%�EiL������M� ��h,��侶"��>'qꡯES�FIf�`��V'�P��o��������'�,�����U��
�f�;�U	v&��j�0ۑ�Zq��]D��������)�]0�sU������F���f���-ݷ�������I�q�(��ô�u�9������$8ݏߢ\��-��*�?�J[�M�ݧ�TC?����+�ߴ�d+R8/�"�RM3�mA0��-���D=qC��}7O�F�G�����m�u�R+�_�I���y�
W	���5(hy�3ϸxFlO�Ӎ�x�"�dI7�G����d���W���o�nʯ���?^�#�wK^"0DO8���;��x�\|(t�Gm[9����GrpK�%�}K�G�2B?�lW�	X�pr.�W�tT��4<v�b����uB�zYY��}9��!�~���C.�O�I�+1���O/?�g�1��a�i�R���1>c-U�_����j��Ϝ�eMJ�
���f5?��u�aM�9�òS���������C�;�o�>��u��z���҉ev�y���_ʊT��=V�Y�xTAA�J��?�@Aׅ܇/@���ԫu���g��v�����r�T~Ƹ~��� V~=Θd�qA��9���]�
P�IPҏd��A<�}��c܁���ؽQs��(|h�_h�M#��1�ϛ�<�F��uze��?�2QzZ)���Qmo�Si����'+e1s��ꗦ��1񫜃"7��O��:j�z"��R?�9����k�{�(ыW ��%hY`� �/�r�J;b��b}��˰r2FR�a
���@jzw�,i��C�p���uNt|�$� ø���d��+EP)�`t��_ج��P�Q]J��amܢ��Y3��-@���� �,>¢9���y�|�Y�����od�&�e�� S�yp����R�.Eca'��aA�l
cXKJph�X��oU���?<o4;o�-b�RH���B	��Q��f��HJov�!��Q�E����pX���L(����Lʦ�Zj����}P�Zs?�<�?N�c�gG�� �c�\�o��Em�	���9`�t�%�ѴyF]_]��X�+��4M=V�t���D�Y/p���p���@��B	�i���Z�f�f�H��Ї�r�l�`D�.��l/�<���M��u�y���M�5{�;�bNw�
%�FMՉ���ρ��h�v� �=���d�[Ӽ!���xt<��������נ���1�w*��n�P&}�)�a临����e�y��9d-P� Ϙ)J}!<w�>���c� N���������T�Q,;����d=_Ԗl*�t�:Xӭ�9Ā�2�i���_�3@/T0;f�/��������KHǋ��(a�}����U|1��%�x�#���g'�M�.h{y5ױFd�߽�ll��8@�ɾ�O�U��t/O��fFR��x����;��Ʌ��+{�� ����L)�!��Od(�o�ɤP�H��O��RV4Yf��Ukȑlq�c�_��ŀ|�c���\)I�����2Ƚ͒V�}W��F34�NP4��@���Q��ڳ�3�}�ХQ�~�`;,Jm���c>�yc���~�t���Ƅ�3�ͱ�7��&a5��tc��3�~���7ۦ]�8�~Bٝ,7[Sb���R!�t����DR�41�Bf��ޛ�OV�1m��,ȭ푒�Y*՞4��(U�	ִ����s�� k���Sj/�g�h�F�M�&f�������.�C"E�k��T̀z��\k����eз�	^��.,�*�]L�-9�^k��0�g���qP8i�E�6Ƴ�)4~�/���h4��ƋV�7���-u?�sp�*�ou���������h>F�~��D��`�~pKWQ��p�O�H��V	�Y m>(�`��ښ쟬]_9<.~��:��)@�/��4��3��;�p��Ó�\|s���E 4/��+���D���r��0�%yU���I�M�B9�U��҂�8����l���+%_��"`��/�f���1�#䃊�A���p}<���nv�J�e(���)��J��>��*w��������S��{��-F�u-�;A8f����m�d&55\i�R��L$�I'"BC�^]�Lf�%��ݓ�1Dg+�Ӿ�l6C,t��I�6-(����J��}����-��՜���̢�E�{a�,Ni����i��~��c�yoNF�e�1�s6�}*�xwì� g8g����en�m*�Kg��T��% �|IC���;s��^�fR�6�s��N��Nʛ2���쌤��K^�+���gjnc#�Z;�~P-oȊ�=Hl���l� ��\��(K����%D���w���@�3���8�5l5f�_ॽ�;�T��ÂYU�������,Ňʅpu��1Ĳb�@����f��!cQ�
�� g�R:_gNQo��o+�>)&B(�J���O%�}�ʶ�lT��̠^ɥ�X2�³���#f�T8��� ��u&��hJ�jvǡ2N�����a3%�;���Sn#��2��R�b>�U�gH������>���v�J]J`%�z�g����w��PEų����o����eo����]�Ct�j���
h�O~�&���4��#�CaT���BW�$��!��{��8�E���o�R[k����#�-�b������Y~o_�^��h�餿 �6)6��<i�^�j34ʼ#�=(a[�2'P���""	������ "�g(���af����Z��ɴGo���n鸣ء��z����e���1�r�z��  v����w�����|�z��i��S��ݵՠAU�Ua˩c=4�1-�`�צ������	E��HW��W���X�7|��r9b�yt*�wV')�P��e�����&��OM�!�s"�dvV'z��3��Jx���,���"�co���l�`Qg�b �G!VJ��%ר ������DǺz���K7>�-��k��*�x�E=G'���͞��wJ?����G����J�:�皂��H�����Q?M�~�N2���s!�D�Bs6`}�fj��~/�dH��/�[����]+�y��@�E�<��L��6c'�@g��ڂj�Ʊ8���e�2ldW����6ł��,��V��7 T[�8�d"��	�>��Z~4�m��h�֥j띔C�B<��S���/��N�����5W�^v$W���p� ha� �|'���>��J��)�*��>H����Q��Q��*#"�頎�u(:��)����~j��N�;�|�x#$�
�] �P&F|�P� �GD}�!VsU���hI��Vz� ���������K�<%�j�)���]�\Ň��.�R"��i}��Ѧ4��r��,*�̭k!{�Y�bVb�s>+�T%ę�'�6�@�i���"òr'��fQ�w�r!�-��Ad������;am�n���n�g�˄*����y�3a1	8%!�&�[��!�v5��.�7*���(�˟�=��*��w<�� }��_��E�2�,�*���[7�
�T��i�8(ܬ��Wd\�q��E	�f����U�J)6��F�f�0�Ѳ�����Ӂf�4'	�.Ro�
�쉦H�2�-q͉�YrH�G�|��N�/�(��+��,{�߻�(�D8�\�9��V�݆$���}n!kq�{`��e{ܪa����Xj!�*-%�3|X_mG��H��\5�§/��g�0P�	u]�5�j~d�T�Oi�#S�
%�%aؘΉ��\�p����݊��w��t+~
c��s���\	uTU�,���rd++G�o�`�X�d�@]�º��2oK#$-��YE�I��`dj�:o�M&��a��:�b�����o��"wꠛ	L7%N�H+��-�z������=m��e�V'�{����;mh��=i@�eo�����C?����E�5-3��F\��- �.�����l�Z�L@C��(T辕��T�K`q5F�Ĝ��۳~&��)��%��ʈt<�-H/�%\a�5�hJBWC��)Ks�K�ف����[d����_&K�]RƎ+gEϯ��8?mAP~�gs�wR���]7��y��{?�|�o3����1 �`�-(P�'�(�y��ݍ�l;������)��,je��~Q@t��!*��d ٦2�׆h��
�)��u"��v��\��B{�u��U��:w"�P�m���&j��X�T	��NazoQ�٤i���4)צ�*Dc�p��tk�x$��߰�������R���]�]�N��F�N���w�F&*���O��)�c�9���߼�w w��#�W� ���^+��|Ǉq��R.�?��E���VD�ɮW���lL ����?��)#��׶PkPz`l�ԘAX'���В������A��/]E���͊�aF�B�Ni17kBN�hq$jST�i4����#���r驽61��ld�Υ�J�7Z]�lo"�״����#q��#H׏\�^��zmE}�{T=!\�ot���"й�G\]x~s�n��=����9d��X��j�HmT��qw��f-�>V���W�d��¥�NV�����ߕ�o��V��j�v��G�A3J&ߒk ��]р�S�&��3qW�k͝)I��{oV�=Vp|Q}�Q���1î4�h?���e"��|s�5�A�~���/��_:5傉*�74Dix��|7j���+i�^l���_ߎ^�������%&�I�;��ķ}~�62϶�����`���4x�Bݞ~�_�N���a����l��H��8�a��LMV�(1O
�+��7v�溘J)�+�?u�2C�bP(�u's�B� 'A��5*�Nut��1A|=�'$)%=��� ����ZH�@�W��ig�o����I9��?��*G��kS�r�]��ݬ�(�����O��[���fg�)˺�h��|*��e��X��J�qy�*��(:G?F˃D�k��r%�'Ѓ�L)�L9�;[BL;WU9�*a�b��.�O�Yw��`��o9
�p��wH��ZXS�J��r'i��w�5�����F�W����(Vᛑ�f��������+���.;�pg�T�����5�g(֏Q:�����!ag�.���7�p���_6��~o��&�н�Qp� �"�<uB��3�b�jƕK���Z��F����Ƿ�r/�Gw�<���T/�JeKy��G���@g����-|1�K71T{��ռ�ccJ+��g�m�t��P��D@�>a���I�v�l�c �CN$��ȴy=j_��dPNZ�@_�߼�Tw���.�e�voW6���"Y�g�ҽEg'	ې=�z�')U�)ݎ]#�8L-;œzs����g|$B�� qk�BK�f�?�V�2�P:��1���K�w�->�&Ĝ�k�leR��p�,g��ݍ��\�K����{˲��bI?�j�N�H®���"_����R�*���V �D�W�B��1n�L���޶ɭ�eO6ME�x�`��g#� �d��SƞؕO6(D�"�����.�� ���*� ����2�j��.>D��� 6N8>O���)�"�j7�ç�8���̾�#�kJl�r.���+l6`��%�rxm�癯uÛ���\X��`X$�R�wk֞�Es%Ǔc�w����ʸGi~��'�������$!hOS���ٺV5Se����Y��� B��E!���D�ai	���v��~oͲ6�7��ye��+�Ϥ:�s�ߝ{ܔF;�|�7=��Ђ��<X݂˒6�^`����|4?��?|���C�M C:��̳0�#�l�Ew�ǈ"��6B�w}3@WaUE x%;��NZXT��G��B�}�5��i�p��J�H؟pvZQ�S�5;�;����W:I�Q;_�����_2����gv+%�M����1u�n����'�֣�ACuX:�kP%��/ʛ'����(�BA]����!?�c�GңtV����&�m������se�`2� �M�A�2��r�/5`]:�LQ,T��Q��?�K�Jb"0-IM�Z��r�麱Y���G8@J��c�d�顝��\�uT?�i�M��<�C��)���#�d�b��[���	��eg?�e��l�q�*)��5����E�\�7��^��]E4���!�U-'�C�6�[���1�kx<5P��V��{
ƎS��ri?$����\���S��r��ޔ��x���{��ƿ@���s�`���%�-v�Um�M(�e������2����
�3{B�$��e�R�Q���%�J^X0���vn�:l�#��y�	u�ܳ�n)��q6{������ w1�,~
u��h�'r�X�[�w��/�x!�C ��;�;�[R9$�����u��-��?ŵ�"�WS�%dK�������ӤAΟB��k����#��c�{a�ʦ�5���d>^�G����z	^�J.�k0O:��@�R�Z��垇�i�2#�q�d�ẇ�ɰ�� H�Zk�Ҿ��W[l�"�ObtfMX���"��(���%(X�N�X��|α�]���`�����b/��;8z{�6�I�����d�5^�oU ���C�P|X��𸰫��,�$/�h�]x��S
�%^�yB�8�Y�{�נ��b?X���4�G�x���e�g���t>���H�#Xe����A����@�K5k�	�e#�#w����ި����c�SvK��S��iI�j+u慚���GC�'��i`���rDu�lCku�ڶ\������;������ ���#��Ȯ�C�x;�����c�V5��Ac	�c���>&U�aM���B��/l�2����Q����ё��3[��+�ƿGYJ����Kȗ�^�����[p��͏U4����wNW�C�d�:��"=�A,���� ���w�z@I�:4����4LP�	0�O^��* �D ��O0���w����m���?�&BAb��Z|�y�]�SK�C~%Rg���aHOm+��jI+b�h+��k1j����{q���,��ke4̵���<ZE/����wa�c��r���Ϣd���w��[3fJn�'>l��|��^
�g�^���Y��\J)�]�b>�U1��S�~�K`��p���{���`�X߭�СJV���k����krU�P�0��&on*v�V5�l]��E>Z
�]�����YK��'���먭�!�^�7vB��9�
�32=+	̻�U\Wx�l�_�ڎx,�F�#q�Ww�'�����G���M��g�϶�y���Qe�TG��ĝt�ؚgϊWפ)�L�P��@�\�Z2�OVO@���j�೦�"(������q+�m�&��Z(�Oz���#xr:�>�Bz*7� �����Խ��U�`�N�ӥ�8ضz!���c�D�?ʶ��X QF��-\��梀d�.f�<�id�^z��P~5<��m�膮4�w��>'(*�n;]Y"Ь{������\�o5���ًg�Q��p+��)\�H��@��)$%hva����;C��$8(2����#�`���o&�P`��󦠭��X����(ʽt��xH�����3%F�K]�;����9)�a��
�����34g�a���H�8:���3:��>���$�N'�?�
qm�e 0����
".�W�ͤ%��wG���˷�$�?����8�Qa��dH$�0>-�I�gWb�K�b�ui=_�Z�P��mY�=)=�U���{Cz��,��?��eTCP�7EŤD���Ӈ���y�;�y�8�vK����KmZ���ouü��ĥQ�����ֳ\� ��+ 7_q�K"��Y4�[� .�֨M�Y:�m�l�$ŧ���v ��B?zo	�s������$,$Vh��ΔU�*d؈�@?��&�τ�B��&b�4���>�d�iɳ$ў�����V��O�c�k4R&�߆T7e&�Xl�]�Tq��Q�?qVh�m@�-��F֏�9b�p�*1��C�}l��l�XÚ\���խ�?|>��j/���Efa
�Ŧ\�J}���NS8��jS>��J�C��X"���ւ�$2��Yǂ��Qb��\g	3ӟ��,�f�B@ˑ��q�ntưٵ�e�:2�dc|��c j�T�տ�6�m�ԝ��N������Eo0~�����(��r:q��9ʜ�	7�&I=.Ka�O鏁�*^~'��2o� �����=�T������d+[+m��G�C:3Oפ�c�7�J�(큄;�^�wkB��k'���:=�Ȗ��n��R��:���"�(�"������.�jt�CK��oEc�G׵�Kw�B�m��ef���ӽ���x��T�o�2�3�����qu�����~eÂ��YI�v�
�v��p��ܔ�"P	�q�'��ا�=lV��y�l�}�D�7/�����$�$�����5D�_�q9�,.�t*�4I.e��'��eM9���X(�+E���M��L؏MR�[��4:v�即HE���L��#"�̀'�0���h�R�R�8β�kI�U�8�C���`������C롽Ͱ�	ƅ���d�ة2	��J��MC�o.����-�7x��x��&t�<7� �H\���dr���q���o#N�X�D��Q����.��d�L�XI�!�k�����r�R� �8$ڹ���6:�����օ�B�
e>�臫���[��:NC���tH~
Bm'�_�vn���o�~��%`�>"��I�;�����`����T�:���I\z�6����)���k�쒦U܎q��v���Ì�@�T�
{EB�o��l�cځo�wr�oe����ua���x�o";�B\֌�<�~��2�A��r���K�gY{�	K{�=��&��Y8jZ��>�	`�����Tګ�p�T�W|Z���&юv�L��L(�(\�.I�4�=#���@p�M���=�y+얆�|?K���9R�I3׶�N�Ϻ։ǒ�I���Rx�A$��hlq1@�{��l�קȴ0s;��iⒸ����u0�壕�r�FGwȚ8W�^_��F�
2ʋZ^�Ǧ(�uO=�mc<�����eZ��}��s� �D���˅d��5��9W�*��Eux%]q�r*4�Eo7�aw�wIȴѪ $?F��� 
����a���w��h/��%�c����h��Q8��Mش�]����t.�)�%6�i$7��Ç��j*��9%�q3�&�̹�L�Hx�塚�ݰ6��Z<� �����,i����l:R�1�O����g���p�*c�]&¶�/��5^�7��ηɘ�㼮�o����?�O/�+�C2W�$Z�3v�alJ+�V@"T�����c<�*(;�t��lZ����U[�^(x�����2vG��iG�ۈ�vz�?KG<�'F�P����6�-�
b7�2����pX蛫3u^�0�4�]o?虏����aT���k�գ�A���$�e7��@�j�	��lyt�/�����t�	�amU��G3�8�ݗ �Al��*-Ӻ#��H4���$���|�{�!�[D:1��c���R��`���NX�o�^�4��X=w�˜;[�"��_��&�B<��f��Zfp�����n�-��z�g����scJ�X�B�:��N�=�:����U�p�7{ev�P_���8ŀ�(Y�6�?�����;��W�l�(���Q�4����B���f3� Y�K����KV�k����� hpܕޘa���Z�!�&�:��c���vx�xJj��Ը㨍!��vI#�̸����,�]f�� d�ԓ�9���T�_u}s�O�٬ѥB�M_��:��\�� ���s��8�]�c���dT��&�Q�G���o��?�oXfeC�\E%���V����ݾ��z�Y_��Us�8��qx��<��rD�_����s��C�?��a���S�����Q��#�=�.9�V|-^��2/F��hD�FþS��ڴv�d������9�rG�������C&�d�?�內�����X�y��Q��g^����������e�9n]1�T��&Ǭ�Bk'�#<J!�^�}a�Mi-��
p�!B��Q�j��?Xq���:![���e!$#"�g����
��]x�d���J�ݪ�����.q���!2���X~!ic�v�d&���O`���^���a<��H3��#�((0^e�������� �a�.R��w���ꓸ�%��ڡO4x��Y�^�{&ځ�����u ���0ߝ<�4�mtqe퐧���az�B��6Se�9�;�vc�`���ȶJM6��՗+R㭆QDXg��A�-�P|��k�*��w(?l?U��M�$���X����M'wi��I�k��PwEE]����*@�ma�"���[���+>���,V�>��p���RI|�s���S6&[rX}%����+h�j#K#���V�rf��+��=��-5�@�ۇ^���)y��&�Q��[Y�"�l�7�I�k���X�+��?�Qͯ��{ӂ�J�lmW���� MH����[�7�œ���^�uH!2��#!R� ]+T�L��7&��Z�/�~f͉���O�h���o�k���%��.T�c��5�S�9�N���_Y���3p��8MnO�|t�VeCH^=\3V��b����J|�i�c6!A�$7��U����$9�W�5��)� 3hhF\�x��j==]/�6_W��ܙN��� �%��Z�W+���AR�U��#����y�h*�p�Vz���q0��hTkR�@�\%�L��oW�Ri�G���),}�Z24���#[�ј�kp��"��솠P(��� �!������(���M��ޕ�a��4�c�r��I!MqgN��=�]�� 8�;=a[ov�4Lk?)(A��'76���n���ԧ�k'�2�]��-[u�G�4ǏhF
�<,��AIE�ܠ����K��t�:�#���1����	��bR<�P��^�?iA� ��,�e��>�L���{:GpҔ��%%�0�f�u�J���o�uZ�hLb���_5&ծ�j�s%�!�E�>�ٞa�B�|9 �R�����ȩo�A��c�y�'MY�8�ɽY@V��y$N{,[Q0��`�o8�"�2o��t�$5풯6j���,���p�"�k�1�u�e:Ĺ����U�\<�x$P֜gw+�^���O���f_Y�"������Eܲb{FJ�T��6�e~YW_�EN!���z���D�}�3�,�Ө�=JD6��`%6���^冕���n0�@f�� �$c��n��z�h��}8d�j��1}(��/`Q����P
�F��dW&֝|������,X=���U}��MhRL��؛��)3��E��#
c�l2%t�4��:إW��}�h"�t:�1���\����Lr�����&	Nn1m�fw}L�'W�mE)�;Ŏ�P:(�0g��p7���U!M;�z>�m�A<�=GO�|#�C��*�݀��~Ntxm��>���=��|a�a5~3UQ�9���C�f��tth��q��>�2���k�����io���Wh]�<H�O��v"�x��m���F�9�:��s"In��%�|9�W�,����c�ͼ���/�����t�kn�J�@pJqb��>���~ԉ�lÖ;8��FG�ׁ�y�p��wo-�����?���Ԓ�k�T�k@�b����[�hz�&��9�Q�\P李z0��j����>ش��֜0��/�UQ��At�<�N?4��K�/ӭmjO����b�F�r���C�_�^3��>O�����_�]��nD�K{�}7� W�P�; ���+�/�U�(����p!�s���uS9�A����4�d��ۀ�l��i�#�I��ݢS�k�GV����?��ע�y�Mj�Z��c���J��9�?7RZջ"\&��Qy�j�Vf �i��%F�a�?c�K&��\�i���$�����Þ�(9��B�)b�<��3��,�ְ��gr�-`��G��{���'�.3�qT����P&���.��
�Y-��;�!K�A���Z���/]�h��9��K��2��	�3:��ڿ����O��X
}��Oqq�����惯	�Tb�)a�j$Q�Ս��WFR�C�]qҋiڑ��&_���`�D�?�\��5p|�S�p
~�#�dƚ�
�S�~�B=�"ܟ\�臽�{6=���燫�v�L2.��"���1V	�:�(D�՟N�*�ٞAܲ�%�o�F9��
���f"�����1Y%,���+���v:��[��tT�j���UΉO���ך�]��~-�:M���U�^hFy҇iI����v��5���(����Zj��^T2�& �)��f������-Y�ܗ�<r��#+9�lA>!J.��O�l�b���lL����x��D͡���IY&�_T� Ɠ ���~��V"+������9�V�P,-,��L���܉��SE;(�4����؟�_�&�x�Ėc�x�����%!'�> ��&����в5�1z��O�?�V\p���XA"���n��q�P+Q6Q�ʠun�{�hJW��0�}�PKK�~�d�8�Q�w},����E��Sܞ�|��_�ĥ ��ɻͧ��Y	 c����gԐ�1lwG���yY�ĕ7�ϳ�v��w'��Jz�3�s2�מ"��G���5��w�Z��S~�IY��UiV�]��G_�g�Eڼ>e7�4s�.S��9�A[�D=�.:��9�{�S�QA�jO]'�P0�U��:�kP���NF�$��bkX�g�Ă�b?��I�kj#Ƽ�_��A}�@_� ����+Qm��Y�!U]��a�LFG�F-�eS\�TK�t��{:L��H��!��k��z���Y���]��wx�fm��T�l#�As�m<�|�BE �b�Ȳ�F��5hMRŧou�ϻ�y��J�ӤmRu�vip
�Zi���7'e+�5���e�bp�^��TqSB_����i{���?1�a��hǦ+�P��j
9Ɍ�*D�;�exҵ�h7H���Aw-a�e#HrR(B�.p�"2�dl:�N{�,���d{�ٍ�Q�v$����~GГ�^b���脻z$�<�|�[�&o��P-�=u� 6�YL��^�j[@���J(C�����`Q���[5��y�!l2)\�N{�ˤ�LIw"��R�xZE8>�P���$�4qJ!�N�RB7oTg�	C��[��싑���o�tX���#��\u��A�{?�G�'LA`Q�����1��}�=W�T����FU�_��t�n!�Z�ϕu:��r"�L�B�L��
�nv����kZ�h�!��|���#�`��;S�j䈊+�!�D�Ih�
�/[�9�'h�I��o�X��:��d8|��V�[�6����T��~���l���{v�Ǟ؊^?P�������`�T��r����]�kd[V�c�D
+]j��r�k������a<�@�������@3����}_d�#��zE�x��s��)V��Yjkg|F�����<OϨ���u�@�y-�@EC6�s���#�����I� SE���XN�ޢ����L���mr�l�H^|�x�v�/�z<�Wc����e��Z��Uo��u j,��)m���t@�S��y�F��
�i��c��^���y��F�H��b����M]�� 
B�$v�C��70��u4`�Y_}���NH��d	�1	
�#��%E���=�2�|�D���,G�듔<O��{4�xK&u���A���*'��Ny�����7*P�S� v��E���ZQ��^Lg�u�\��,'U��p��備��蜫�Wk�B�].���7U�Di$�qQ(D�h{����t8r��ZV�S�X��y'�2�E����f��X|��.�B�>9>��p��H|�#-���x&O'�)
�߈�ҟ�1��2����h��#��y�"�9�9`2C�<_2,¡fGʟ�r��xb9CB�cI�嫎��°u�2���"�D&ʹ\x���aL+�%S,��,u�7����iƩ�*�"��ɸ��@����<�&��0�Q<~T�h�Y���x�w5��P��v��@����ٳ�:�����e��z���I�������(��^a��
s�!�o�a�,T��HAJ9�|���b�v���t��W��u�dR�BZ��g�j%Jf�2�!V<�-�������%���ʫ?�`bMV/,��-�/|&l�9����3M�~��כH�ՠ%���#��?�H&�_z2&zИ���ĝ���aK�٫�+[}�Z%oa���HRF[j�O���Zf��Fq��i��8+b`�Xy�SV����*���z�����E�|w���s�b;�����RnV���q�������sC�|0�6C�j��B�븋k s�~��2�2;�O��e�8���BU���Xa N����W,��j�V�3B����?��[M�6�h_�����|�O��թ{e�HQ,�Q��.�_�M��~���@��-��e^�ڵu���R�1�Љ>�sF��M�v��V�U�Q֯f�ځ�v�#�-[y~��~�*���b��=dC*�)� �Єlw q	s�/|�p@؞4�T`f��,��be�X/��J�3�I�ȡ�t^�_[\hv[�F"(�Xv`w�g��/Cg���luD0U�qTq���>�!2ǚ���XM��.������/	�nh���0��#1�_��{͕��&��s�5��w����=Yk�av��+���F�S>|����q:h�~z�tKLǉ�����R��S�=Z����:|�L����U@��*Rk�v�n��@k�
<�7��<R����6�t�B%�q��tc��r\G���Ae_p�e���{m�_�@n#6x����#�YG�\�Ǻ��@�����*|b��{6W",l8Wluc9aF�p5��v�?�&��`�:Ͳ�4گ�h,�j��3�rb�d��؜[2�<>V,�t������镕�w���?|J�L]��bվz��]n[
�}�:<�(c��*���w���Vdh4�ͩ9m��S���`#O˜�;2����у���m�\�.hNZ����ٺ���Ǘd=;�$��lߏ&�t�>�̑4j#xn��'�<Sx�nJ7V+Gb1Y�$�*#$n�`U��3�c�+��U�C���`��"��7v��t-���_ȩ$j��OC�z��kv�b�ԽO��vjy�ư<�8P�����L1}5��гiw�c�\E[9[�T�E�� �X�z��	gz�(�!
��4-��K�7��\�iyO�sZ�DKã5����.��)�z�^� Af��%ϧ �H#�x��.�������M7^0�E��;q��&Lמ�ցO�13~��D=<��4s�z7�l�_u�������n',B�dAX�I����J�����b���)����;�۷���$��x
��y`�]�
H$O��*�`+$5�gSϜٟF[��$5�cg�g���{f�$�L��SZa����uq"��\':�:{�w�t�ku�ЎT���嶆���l�P���7t����<-�ӂQ?];�`M��$�L`���5%$]NO��м>P���[)}��페�Q� W��O��ϵ���f�H^,}�A\��s���5�!�o�ɤ��O��%��Gc�zY�N�(�X4~�q8Vk�_��4��-ߖ��?J����ӡE�c���4���J�o��h/�p��q_�9?n>�&X5F32�4��$�!�v'oDM�і8�/�_ �r6TUw]5
`��I�"�ߔ�p)`���3���!I6�d�q*3��a7i�\���a�\6�Gv����m}޾J�[��N߫��������e.}�p�e?���$#hB"�Di�l���pz��r$#�����,ջ�e%{�19�������l�-��A Fw�V7�b���`�5�7c@-��5�2��� T���`�&�(LZ|s�ǽ=ފ���?���?lu��'��$w.�E��;����h+�&���U�Q~gҕ����:)��R�7�5��;�:f7!�y36I;->��=��N=��2�4��jT�+;�c�cvf�F�o^
�[���3Y�nz�ɤ��daO@U��! ǽ�^�����|-{��U�z[�4#�,�%�7�(h�,ǫ1�?<Ԁ�C���e�m3��v�{��1��>��g)t��,$"���j�o(}[u�Јܘ]&b����LAO��#�s/gu<�5[}�(�R(�w���C ƌa�����G�Tt�+,����h�qq]bx��T��?��K@�m�K�����@�S
��LE8�7���T�?W�Mr���
A��?�t:��w�e0�'�