��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�!��
��%Y l�׾���b�����CK��P��Q�$���}
�&<�Ī�7=��}�7I��q��p���f�8�Q�L��.?�-N�#�F���OX�2�p$W�����. g�w?y �I�k��X����''��J6F�2�`
����Xa6�R�`onЃIϽ�G{9���9pQ�9G���7��xL&M��C|u��2~�����xg���A�.�,���g��T�H��	!ǘj�X�f�
��1M	�u�`�c�n��X$�����A����_��L�0$����i�>O��B�tK�7�Kfѓ����i�}ې��は6QL��g�+��]��Oh��i�ub���k`V����hP��M7mHx�Mu�I�6�����|E�\t�u��$�be"��=8��8X� p�Уր٥����"Mg@��<�B�8Cf���@�����q�n8��N!k�V�C�y��y^d'8Sp��ʃ�N��F��A[���7�_v\oL�����^m��d��щ����1�ڀ�BK�EC��nkA����],2��6��/������cV=2:05&�V8ܩ	[��|�,m��NcP�c}��Hʓ����V[{}uf�`����d^m:�Ѱ6.�:�udB=/�~`q� G�l1�M#��Qד
1@	��22��n��Sg�&s^L,�S&B'�����h�nxwT�q���K,n[��c>�/�F�p4}��������_C\�]0[�X�X���ΡQ9��Xƞ����� +�������6���b�2()�sl*"���IH��^� �o�|(�j\Z��~Ȟ�t�5��b�h� {�§�́��\q�YwMO���� M�?��2D{!՜.�(\oh�a�}a�4�K~�YR��/�Nl�"�%"����"NT]a�}�����5c�I��5�u��ȯ�3ÿf��q�ed��(F�����n��d ��*6��!B�����|��W3���D���Z
�U��D{�]�nJ��2��LǔlP&�s��UI��3rͽ�+���x���>� &ÉRw�>�2���������&�;�/�{�-�r���/l�ӿ�p��U�/\�W[�%Q�$�/�<Z}����Q"e���bfs��z�G������gG�ꊭ��Pa~� J�
�����c��p�Fɠ���I��ك��#��s�#&q�Wu����d|M�F)ލB�jŒa�w/��d�T=�f���ս���e�D'�z�eo�7���@/<a�W�e�O��nN�|��C�S?�N�6�$��p���a�����.��qj��X��?_�d}D�b���L�C���E`������1a����}m��5�Q@�M4��KΓ����AR���Q�DP��J�`�����@1� ��˂�׷8J��F旅k[8W <��8��M�	�	��\��4�_�_]:AA�{�à ��f�C�Őb9��@d���t�`��{�Ʀ�V��
�픇��=�G��L�g�m�r���`�\!���f=*9�\�c�_�������nIN䅂���aV�p�*d�}��A���_�^��<I�bZ��:�d̛2�p"�[>AE �6܏3�H�
-�¶����Y�ڬ��J�{b֪���v<�S؆�	r/���a��{C�K`�
¼�ĸ�W�r�Qc��I�**$��򣢡J����-�0�n;[d<�IC��vw�B"$�>����E5�%蛴H�'U֯��Z�z���U�������_�.p. �M����cg���v�Ů��K։��,D�8����2R�M��u�l�+7�o�߬N� kD�U�����������$X��(�l��Aţ%��s��¬]�K��J�NC��Ⴎ��կ�!�F���FW3��{�ʯ	7�7u��.
b'[�C�� �3Xo��Վ|-�K?uq(_�� �i��_v��� �//]�OO	�~Vx�[U�E��Q7ط����.n1ǼC�6�R�L�����~ԅ=����=����*��rw>(�d�Y��
�m�}/KO�+�x����F�}�����ʾ������P�j:�9"���I��kֲ��#9����5*#����8�~@r����)=���5��d�H��Qҋ����昔���f$J�5��T�ȵ\��t֘�H�ՠ
SRT�u��m�y�,�u1u�Zb���	��*��;+����;�#��0�*�r��!��,+��g��dR=(���NT�c���-B����+��(��9�f�«=���Mߖ���d`!�q�޳60��D�!��L�z��Ź���>��Pю���_ĆFu�,u?v�&�fɝ��5�:�cŕ^JO�V��CE��4
�8���}ڶ:c!�tԆܮ7�4Ȝ���p��eA�d��E�k)_o +a��#����VC�{������d3�H�H���*���!�!��=&�`�R��y�7j��ub��f�D~�G�2ܕ��+�y��5��g�Z9�|"GЫaߑ��A����&�q.��=(������V۷-hcv�4{x���`hE���}��(Lu�@�\�W��u�]?�k�G��q���Af&7�l��X�ip��I�{�=s��e��j�Bs�[�Ej�S�8$���w�`NE���v�{�E$d�z���T�v!��!h��k�h���q��3�����T��k���DMaEm�\��A��ǭM�Z�齗������[��C��ŧ�|�:,M
���{Eߛ*�3n�>�Dby�7"<`	���s�ko=����F���_7vbwѿ�٭��]ΚS��;��S��B�t��h�f�d�KU�%7�2��K�C����"��0�c;%dSK�c9TX����!�,2|��RJRwN7��Su����x�*���4).x~�5�� Wxh��:����KqK��m_�'�m|��-R��5	rG��$�mn�z7R)�$|-L���:�iO�v��o�0,�:bFq)��e��~����Q��0g'��b�u*k��=�F�{[axY!R��=V��+ �ۛ��'�����h=�bT7.����=D��B�w����x���]��%�Wr���/���Yڟ�lDCʙп�v2�L�Ԭ�^ �n?:�.P��*o!��^�����_t���4�a�.��؜���jY��)�>G8��WGA
��:�l��＝�|m��#�}�@��V���W�n�<wz:�cx���f�@׃[Q�+���Xm놞Bl���e�ADJdQ��9W�l��8��>Ğ��'0���Jj�3��S)M�Zr�0���Eko;�/h'�M8$we��U�\%v7Z35r�pd�GK���x�HJ���	2#K
.0#�F���[4����]<Y�.�L�!��6I}���2a.޲��>��8ߒ���r3y�����ax��(����xՈ�4�%F���Sȟ���;��O$f�Nm���V�\�wQ��y���!ȁ�E6��x+�!;�-_ �FC���@pq,Kyt��2��x6��R^��>�"Qe�Pԁ���?J2��@D}���\iC0��e-˂��:p�����}q�X���-��E���5�����q�����tD��֫�Q��dHk�*��fČ�#(��C�/�G�1&�	7v��Ɔ��u�%��\e��Ro�9z�6��O*���S�0�I��*b��ȋI~�10�BECu�u�֭j�[҂�PY9��	2�!RHm��ߌ����b7�� i�uK\��]̈́����y��vg;gfդ}~Vc&{�����]&Ü���9l���w-;��9��¡oMF��'�(������ǽ�j�L�\R'����Mm
��-Gn�/8��P&���PB��N�X/`�H&���Le}�֌XlkX�@�K���s ��T� @O�$��1�~�$)&b�)ˏW���A:�@��f�T���,��vI#A��P� ]vwԈ�O{�:���PÕ(��x�Tn�'L����1��_#�'�4�E�@�/�6%Q�d4�+1&�������<�����G�C�Nia�E���C�X=���^t}6���w�\�0Z�+3>����\��f�^}^@c�"��(�z�+p�3�o6^c�;�WG�`T]�>�v��V��L������q��;�YQ1��]�
�dF��pH����z�I��ٟ���o�U���93�6d��ʥB �#����ajB*?���9m39bm�k>86sE��Ϯ`k���mC������R�OLS��Iؽ�s/eĂi�6���O��:-��lؐ�<�s�񇺲RO���y��(2��ѷ؁h�	}(P�Y�Ngj!H����3�_��:
�P����$�m�s�'0!��d�H��c��嫠�J�ĺ�s�^��H13sJ����@Z��bdx�W���?}�.��VJ��&͑|^ӂ�;���G�ю��+���	TVՖ�C�3i��"��~X�E���c����z$h�Ӕ��S��d+��^M�ew�j�VX�N}]r�Y�T>�?s$�,�dy�X��z���8R���K���<H��hi�4�h\����ߖ��W�GƐo��H6p����@K}��2��
�TvK٪V�`}p��!z��<Q"wK�R+/)��L$D�@�)��<C�wޓ��  ���5��q��H(`��l�z�@lD�C��)IB�`��&�$�ʋ��Ir���(�-�_��2��y���M��S}Ц���ah���8�O�	*�#BfR@A�M7�z��?�Hw�i���2X�4��i��}��Yzy���j��0%5�p5��IfD~��q��x4�>5G���q�0���M�t���>�t8�a��* P�#G2۷9cv@�_��l�K���?z����\N���o/��Џ2�|$�]�5��Uh}��������9���s�.�Ds�}�r�r�S���ϐ���	#�2UG�0:0^�*�_Ys���}�m��"<�:Wni�`��v�CH]H�9�inC�� �[$��JpjD� B���(�.{�������B�5�<O�L�fž�)����>�}��4)3fcT&���Rb>��? ,P���������s�UR�L��|�K�3�D�btE����
����{jY�����7츅�s�.%�o٨��nX�/5 y_O�TY2�=����ui!y	Ǆ7��"S4����.��kn0����$rt�|���&5�vCcx�ܽ�-o3t��C��*���â����w�EФ�����1�X�<���+�D�Jl�Fk��tm�M7�!ߥ��t�}&|��"�O�?4�-�Q�~1���̱��̓u5_*+�Vέ�#=5����T�t�[I~�T�������Bv�U��/N�#�."�]�� IZ��Bwz��Y�q��ܗ"���lFr�����?j�I�C�����1r����<���[�XGPS��w�y�������/7�pUy�QQ��0��.qǃ�n���qQq���	���Z3����'���F�%��R�m_��H����2���6ҾN뙸�>Fx�;0~n�⟶)��۱����i:=(54��&�̂sm
��_���LPm��I�w���Z���)>7=��x����o$�
�#�¿)<�,e֞ł��&x#�y�B����֬/t�1"sJ�ٹu�����Tb����K��g~S�	���ey�����E�(bNӡ�1�'��h8t�ԍ@+%�"Xx#b���W  `�.��
�q6��P��������L��� ����v�Β����ρB�Ox�o[���1e'���w1�S+��iUT�=U�<ޱ��+���	`3��s�����_8	jjw�94��Cy�G�o=pd���"An�L��]~��c�K�T��N�YqY�v�X1�����~��p�/�u���o���D���F��S
�Q>ɺ}���oeU��/���U���Z�z��p�UTmzY�f�3H��{�E�I��;�Bœ��e�5��>��W�@\VR/��43�҃�×�=�5��� ���ׁ���K2���p�v��n����L]D��Q��E��S5�����v���a�%�s�oo���*á��f�uX#4��6Fl��u�a���,��	I�������O/z�-����t���,��	������4��G������/�K-{.�o����X�pU��x������_���p*B�e��;�[�R�����H����<�f��<PN�x1M5CǶ��������eKr�' u��x�fo��e�Dw�6GLw�l'ϒ<l�7$�X���+M�P��-���d���/��t{���6+X��J��t��Ů�w�R�nC(�B��P�рo`��U����{+-P9���b4��+��ϧ�iP��vg= ��TA��H���y���)� 3�#O�j�S��������Z�����fv'$,��:
�{$-��l����t��0Nl�Vk�iP�0�"ߙ|�n������!���5E���#���
ܾ*�A�1��/h�[��\!��_��ň���c�����Up(���*��O�c�)勧�At�]�ï�����=�����|�����f[R6o�e5 �t��V�u�p@+aW�`g9�J`�m�hU. ΋z���.����(u?��qw�еi�)��Y�4_揍Љ�ÊG�(8퀾Q/���4�}*�`�	 �HSn�����h{1$�F�r�~��y��WD1�	��ʉ��m&��|B< �ϭ��O��Ka�n�q�8�f�%������+4�fX��vs[G�(�Z߲ۡoR+�M��W�������u�*�9JX�WɌ���t�'?�=R�EMa���fܗk���Ͽ	�@�Ɏ�v,�s�ƞ�`=��#�i�N_O���?d���;�$�����.��M��۶�(��l�7C�Sm_��� �t�-�������q ��
�H������:��^��c3iX����^k�.��yЊe$��8K��:8��=TTmO�ʟ|(�JDC��ʄ�C�aL���:*���;p<��ռ�Uq��o�E~Ɇ��T r���b�%���^u�BgB��Bm�Ӝ�(��̜�j��xc'=f<������<9
��VO>�G�a�io[���R!�XB+���~?�=���οG@�
�@����|J��u� ��6M+z002 B�\��=.)��y2���j���7�a^(/^�J��>�A:�_���B���]�.M�2c�G���"�W�|Ч�C�I6IX�K�2s�p5�66�l�s���x"ت�9�O�����$�S�_�Aޖ,a�.v���n����- ��;_��$lC]C��",�5�� �T
g;��%�ty�,��JP`�L_��{ D`E.*���ܛ��`W�n��X��>l�FM��=�ň�	^ڕ��4Ұ�~ �K���h���D{\s�?,��k�__�Z0cz�E�.	mX�v��ġ��1T�eڷ�v���8&/�����"�rw��E���e�R��4�sz;�"V�r��a�l�Z�RQh%]��Z��5�ؼ�e���Of�6-�1:��Ϣ"�r2�ALG����7K�;'A�;�C����r��9/���4� =��3�N�h������w�g�X�l�[���v��~cy�g(�ł�kŇ;������>����Ko0Y����A�T�tq�AQ���DH�f�^��৉������$K�6Jɶ�'꫱u:Qvr̎,�ATE���M��J���Ƥ��.;�	!`����?�o`��#��@��z�e�B�U���ϖa���1g��\��4��-ʉQ�	@tV*�y�,Sx42T��.֠����$��~�~�������U���5�M6�d���Ҩr�c ��;-�����)�2<�%�?"�J���Z��]n��+�:<j�Tg�9��������_�%$��� �V��$n~��J�𷓲�,�Fd��~��b�M7��J��#BoƉ�,I�1��|d�a�A��`�%�}�m�B�_��#������-�<�t�YIw��e�Z��Ʌ�Hy���qS�ccٲT�B�b�����}��Bc�Bj��D�����?��|`�y#b�CJP'0z�[���9Qx3�Mb���e/4��-[��I�M��g���k���}x���D�$5ׄ�O_���V���a8�H�S`@S*���.��l��!y���Y��#>�4aO��ѪL�trZ�"I�;:Ց���o����V������0V$j�0/H���R#֑|TQ{�`�TiTU}`�w��C�����U�!��P�b֮�ئ��' T���W�%���^��t(��41�| +?��a" =��������M��[}�Z:y��h����a���IKFc������>*;�S���nC=����.�� Z��x�.i<�s�2��S#�9YĻ�k'��׽�o/��F��j;Ә����٦��M���(j+��e�&�Lc��`A9��j��3"XgϚE:�O��
+2<%�[ ��	Z�*-�5&TP�m򡜕�
�:��ǒ7����'��{�9_��˒M��h��?�� �
'�ao_=m��eT��&n������l�Ϳ��������ㆾ�>fYJfH�̥�����"하2���w��ԅF#l�:�5������XyR�=Q��Cy�)���4�Xt9�+o�R̍�{I�Ե����1��g/��n=IF`���dB�~���xס�fI�z�kU�L���*�f�#ړJ��pӹP�t�Ɉ���d�!��EϦ��F�������$l��80/w��X-q/�PL�>��>���%�v!	gk�/iγJ'�b-T:��ZfE��x�/G��	��B;ءz4�A��Y�5��V���&�S|� S�?u��b]��7J�ݼ|��C�Є*�$�(�[��S�ռ O�g6%�N�.UF����R昧�!�w$��}DĞrWhH��^}�AS8y\����G�ٞ�c#m�vU��"���Ѭ�r�[y{��F�c�CO5�諭%��J$����8����(=�P1���!O�
�$/�_|[���V���}%~�Y���3���NP��% �UK^p0�6�Eu�"�cQG��<x������v�%��"�iL���@���K��j�����O ��[���$i|:_�)x��x��x��{��I|#9%Q/���{����n3:���r}��RWֲ�g#��W����E��܃��O�)�����H���\NE���������,_��u�*��^����H�B�]$V7j�5�?KXwݘpf�ہIXj�6R;I���^V�> �l]���B��}�R�ald�Ԏ�j�w�
#�`�P�tR��{,z/vǎ�ˌ��t�h"]X�7�n#����kC�e�yG�q��kTQᪿ.�qJ1UR]�Ί�z+�G9������W�}��
�b��k�1��l���s^�*�Tu����WI�����Cj$V]�@�� ����a�Er�Ԕ���k�޲�K�8��W�hv�ƿzR��tZ\�k����gfI �6�*ۻ5�:��~F�^݇�=<-�����Q����A��;S��&���0�:|*�W��ξ/�S��'8lP�6��.SU�u�w���!�V�|�s�-�GR
��4j�n��	d�Ä��=�D��o��+l�����Vh�-�i
�'���!7����|l��ǩX�h���A�����ʍHow��C���t��ʒ*��N��h��Ez+���=W-ˠ*�><_�2O��VG�V� ����|w�$��:źsW8S
d ��t�f.0�o���� ���	�S}<ޫ�w��[N��
QT�9k�^�RLqnDru8�0(C5r��Ɯp�/�y�O��g<�3�c����}�iɛ
Άz�?�T&X���G��T�p�O8,2�P����R�y��Ʀ��
gZA��Ԩ��r��.|��$�.�^��/^8\_"%2�JˌRn`ps��yA%�}�;ջ_��y�[�%\0�eV�Ef������7� �$��ٜV�M��[8�I���/7�l,����,�r�����~%@[hDs����Mǫ�a�W=���o��U�Y��-��K����q�@d����r��2?��w�����P�N�%��3F���Q?��.(���ª��+�?gIo������<gF{�5��\g���GA�n��;���A�U_rYO`I��17�q�z*r�?���_%6!� ���p,|�_'�T�C��gfg��p����_�Dܕ��5�����T3���!(�eT�� ����v�>q���"k2Ж�g�2��}��|I��}|h�oo㏜�\1�J(Ŧ�6���!���!BX ���7@=l��#j�>�hW�z�%0�Џ��[���3k1�R�Fs�$e���1_�S7���'��(8�iK�K�S�.�GZ����4��r��y�����G��K�cm߀V��)�ﾞ�������O�1_]l�:�ձ��N�_W���ھg[�h��;�fQ��fP>=KȨ��:ɫ1#��52"�B�a(�����y���|k�_�KbQ�j�>��m6��� �PU�E�ՠk���ə�Q*�߰;�V1�qğ�:�N����賵�����@��HQF��i&�rZ�`W���~5^��D�Af��7	���iSv�1Y����'7E�����c�����0��(�����l{���]��,R�x
��j%m}�
h[�*v����e�	]=7zD� ��&H����H���p`�y�_.��L%
hb��N휄 	b
:��{�����<��F�ۤ����5���Y�6�[�\'j�7�<��.�Wǈ�;Y{���dVN(<?�����޵�����F]�פ2�-���?A�äۯB?GgdD{�x#�
K��C��>��d;�Wqv��g?A}S�\�%��l\姲R���	��\���I4���O��2.�xfk7WP�3(1��3P�d�y!��u�(��jDi5<K��G��k�@[U�t$����_�͇;8����鱆_\�!�Iku���
o���I�-p�7��8��LX�`n >u������T1J-�o��+��ʳ	�
M��q'P�84H�K�W�G�z:�J��-ҡҤ)}���V*`��ʶ����\�NP�y�S�����!a,I�����Q���n��\�����<��8�,���KH�-	l��]vU�͚{Y|�{������a��QUt���i�,�6ym(_���O�(�����+�V�R����F�76eq�m���3�ba�	1��Xِ����I�5,��%�:����eUifU�BNP�WR���V�کPU~���m7ͥt�8E�S�a�p�Z�K�3����{m��p����.�h���6���b���zn�y��|�(+�S$k�*e�-���mL
��X�y���~�����{�-��	�zu���
�>��������ʠ�������Gs�R�y��C�[�QʟwT�ֳ����~�7+�>�ΛCQ�r$#��)χ���?Yԙ�p�R$�$S��%kZs��X��KV�@=Q2yߦ�nuBŏ�zN�0�hdĴ�����ύ��X����Z�Ia�ܴ,2�������.�NtzL,3��$�krտhx�s�.��x�)��u;l�%�~XǾ(� ��7� ���=�t`��ǹ�`��.c��Ӵ�Yv���u�0�r���+_�zt$���ض��栨����C��vx�f~b�������ι�ڲa��􂧲:��t�C��m���Z4���͍FGI�WD�"p�\�v�1%$�W�2�'��uN�:��a6�J꺃L��P~���_�SfȼV*�,%v�dc�dvW��Mx�,�8�,��n�Y-V��N����_3(*�jg��t����4�|��~>Tt�'�09�@��a���ʶ��5#k�%�Y��1r鋌Ul͛k����i 黆��f�~

�1� ���O|lAH�]͌� tS;S���x>�8���XN 3���:�<�w ��*��z�4�o?H���W"����x�Q(4��
G�!�w���Y�����}��;��e����E9$��c�:PD��b�Z@�g<�����Big����Z�m�P�:�����"�Gn���?*� ��5��L�#2��[���L���Я�BLa����T(%)�-���HvkZa��£�̹Ĉ���-�s�Ɓ���"����vIDkϘ����n/����P|��H<�ߚ��a�a��m���nd�4��]/S�BH �Xp����x���&��x��J�e���"G�!�;6~{�~��W������¶����,*�J��/�,��,(�)���X�_ճ],��u�T�13��U�/�@e�'m�g�� hٜ>s�r�YF�O˘muQ��p`�˴�L-���D�#�@�=x�I��D9��M�XQU/]H�s�i��C1Li$��)��6F+��L���|�8���kooF�޵o�rI�����G��y,��2���&�1=ӫd���z�P�5�{��l�J)���N/�^�(jJ��F�X��\�t�;sium��D�w�F,6FU	�B9��4�r��� ��E�=�������?��.{�Թ��x��;���%�*���uX\�L��mfx4��C���aGyɭ�h������i��Yj��B���f��n�<i��s̭�]�g��˵���-q���Oh��Զ٥���N�	6Vh�V.#~�{�4gp�{�kg�̖��{�J�~�5��%D�a�4H��H���6/u���nލj!w�`�� O/q�
x�ċ��Ӹ���h3U�&�-�v�--8f�z1�ܡE�DaG��#�ޚ4y"X������C�񦮙Y�D$������'[��3�D�c:�l��R�R`����A^�e�r�=	��޼)[�ޠY�$�{� �H�{�]:g)��]ef��q!�!��q�,����<'���8�	�N�Ρ����ƘV��[��es#!��(�Z1m�4٨����I��$�<�^�2Q@�<�+�H�y凔�Evs���=}������GJ��P�B���vk�i�j�����0z�a/���{8��+z�Z�(������Q؟�:ޏ�O���}|�Z��!�S�D�~ �߬��9�>rf��Ů/��[[)ͤw>[5�Ț��twc԰hx�E'S=T�Τ�ۏ���gN��f/�Z8�����q��H�����
���8����U���',��=r)*=0>HI�$��Ftun73?��,�������8�9��L���:�%t�CcN�]p`[p���Ĵ�'w仭ڌz��-��vZ�� �Lz�o�Q�j�;��4N�`م/�J���{w
T�n���W�nȫ�h�)�;�~�Xhu5��˚�ڂЪ��й�!��ro�t|aA�R�a�<߰	fS�L|V�y%R�Cލ�o('o���;�]�@�q���S�ߖ��/S3s�^@l:��cv���:2���2�����7�Y�1/$�#����"��zF��2��,�)#>�\���L�����ٟNҨP��?v���XƏX[����T��� � q`Njn2gz��q[
n��g3�v��x�t㫾,�N��2����K�P8gjXU�\P'y ���8���?����-��-uA�d�D�Z��'�$V�,b��h`A�0�[\@K�*r���8H��M�[��B. �"�cՙ	1�J���T �����5�������nW�(�2(U��u�����⮬� s�^s�3=0!����b���ˆ��c�R��J�h��I6v��jLٮ�G�h[��Q�$��.�u�0̤L��U�6��K�yMo�0�z�Շ��_�n3��)��� s���FVdjk�����r�(�^|?�d幚��d��T��n�j�%�Cڒ�4Ɍ�{lBX��>/���\n
�|��9��/�H&�p4 f6�l��S�i�U'��^�mk3���c*���>KϻXg��؆��{H�M������R�S~�xPHG��<ʔ���2�BC�D��'5ߊI�B��:#1���Pv]Z�$:
|P6��Mib���b�ن�Y pG��2۸M���ۼ�A�M�60�Z��j�*-��~\�GxlH��E��DH�;^�_Y<�Ƀ��'o�@�����N�]��җ);7�'-iC���۱�}�??Nk�@T�(�JZH��
?���_�hQ���m�D�v��Ʒ���T�2f�>���x-�#���,�A���	
ӥ!�5�"D��o��[r�B5K2�2�8Mb�3@� Ҿ`#��= e�7[�e�K!�:Q��3����ރQ
]!Um�w��L�^��Q5�iА�b8�=)�� ��ou��PD�;d,^_$�8@9�_����+���A������H{ۗ����ؓy�][r����5	�=�)�J��?|���t�c*F���l<�p��Y  ZJ!v��e9n�K�Y�K�c���O�]��T���*Q.�˫����x�p��.� �/����|�?�c�Aqhl���*��6�#r~�O���I�Ң�xw�R��	)_���w ��=o�ϿB%âw@Ŕ�������I~���=!#1�^�1�\t�T:�ZJ@��Y0���P�8�r��(>"�O�=�M�B7ʴ�F����D.�8i w~��1������xa%��O���-`�r�F%�RNK&U ��w˱��"�Ejo�����:�z����a�d�|��;�;�Ċ��"�JӺ�m�zx^��8�uPV�Ԝ�p<)5!Z��Zb�	U�@"����%+�Q(O%t�f�ƏN�j'���*oJ?J�uxE��o#�@�i$�9'_��JȎ���Z9"]<
�n`u'��}��:h� ���W��Z���v�*�VC!�_#��Y�ju�)���jrrނ�����J_Fk�P�\b�kz���r�U0_��u$֓�8��2�w9�mMd�!�����8�n�pQ��m�8��ǮRs��N����oO��`��!c���F��^�ԦlH���`96*ɟ���N��q�G�
���t����{ ��4s�/��"�^D>͉�{>�b	
5���C�PO��|�TWS,�*�W����,ѫ'�/«Z���Ke�AQ�W�:�Me�^�(���d�!g4�"�uƗ�^%�`Aj�b_�tj�_U|�۔Σ*I�wT�GǴ{Y ���B~�`:��@��̤���ڞ�)�T4,5,@I���=%�e"��1nH�t��(�+w�KS4�P�lt+2	��h�[��!���ň�����N��O�C�/����Q.sC'f��3����2]��.�����K�G`����j�xm�F�z%f��6����$��U��	cS��:苸�h�|Zr��L�S]<2[oN�~ѥ�9;�Fw���@1�`����YKG�EX� J}���ʧ���=½:ǵe��7=��`��H��e2�7��c��+�ܬ��&�Ըo���U��ifsbO�x~��4�^JnT���Q�=)TR>���l{G^���/�V-M�Q>C�R������uN� �~��ɥ�K�8\|�֠/u�@+��P�µ!t�Y8c��pe8��I���l�y���@b��M]��w`k��U6N݄�IM�]�L�4g�pq��L�\��b�v�L,��nd���Y��v�{��>Vu�t�����s%+���r\�[ v� W�m$��]��7�5Kn���#�S"	�� �)�2����(P�n��Ԗ���h���}�:+�`Z���i�S(�֮�/	��r��7#�L���25�0�탵ݑV5�EG�}t9��VR��L]���%b�ߐ���_�̤b��2,Sѡy��y�b����#o1�P�_I�y����:
Z�O��M#�Ũۗ����(ǜ��XM��Љ\y�&��h�0��\߆�S�^Cc�F�,֙Z�":-�se!ג��$}�B��
�ez'ϸ�	H&�8?����5O�M��_�3�2�v�v�n�	<3� ��s �?0�ZN�ΐ���z�Q��c;ע�I�(���$���e�p�I���}��
#�GNF��t;x���z�`_���>��,�n"K��(	���P_E逭��Z2�!��%R;�;��D�#��5?�������>�#�̓\����<�6��la���}ۍyD2�ªI�����%���5���X�V�7����"4.�4|5�����)(ux@*�}r0��ӻ����q��l�Ţ7B�J�6;y��$�zr���=n.ٲ1G�I�͒���pG�#�m:$i� �)	�P��2�@y&"�u��w����<�Q�L�J;�Ε0��8p��	K�
��t��P���>}�Q.h��ذ�N��՜ϳ)�n��mi1�z�M�z�T���������#������ls���l�(Θlݟ��,4�:��ի�&�d�8$�|q��h@e
b4��H�k;�.�̴˜�aV�<�ׯl_���Kc�V?��7�bFrw=k(p�F����w3-,M���c��2p1+yn8{Lj��STJ���a2e_�Q�ͺ���0�oQ���R�#��eTe�M�QKy%�S&&�_S��s�J��6Br��,ܣ �g�s�Р�>_�s(����b���X�nb{���RdF�c�Gb��)%��A��b�ѭ����~���<.�u{y6�d}�U$�1���V�|�Fs�R>��	^
f��л��Y;�^;���� �H����[�reu�v]cꥳE�Ev���3N߬�5&��=�<�O�˃���S�B�A�r��n"����x�ݺX�I���>��S&�]?�d��0�C�d-=c�Q��ߛə����qev^ݤ�f>e;�9R"�l�:-���ȡD�� ����v�c�������rU��e>�0�W�J::�����(�K��r[M������v��!¢%�rX�M�.�,��J C/�'X�Oև*Frjѷ.#)s����i����VW&j���qo�_H���Z KU�o*]����<���4�1�ev#W/��ӏ�_�5|eۡ�6_
�GI���2��Bu��MF�8��W�����@�Ր?�ߔ�_�H$�GH0�~�K���=@ԗ����� S�`�:k��� ���|I	+훧�8Lb��"N+Y�&{O�Q��>{��r�񝄣u�����VTy�3=Mm��$�ccL-�K��OП��x�9 �#|:t�C��mV9Tec$��8GnO�����	թ�l�ZM����-mјM�+U����,U�x�ߘxr��؁[�88��}Ǟ�&_"+j( ���}���Y��~oGoA��1��ߝ9��A`}P��Bx�NF����z�.}�-ٔ#�u�A�l|�]=�[��ڕJ�g�J�^(��z�
���t:���0h:P�T7�גDKhoY�gM���3䗙cZ�PS׿6�ﳬJ��}�E<�a���� ��L�
��
(D$y��M�+�G�=��\�U��9��̞���x�pd��Ϭ0�uv��\z�<�e�e��u��"�/�5�p}��D��}	�Q��v�G������?�g��TQ�PӘ����[?��H�����{�����K^�e5#x/�h?P@,+�G,du�	/�P�3��P���葲�l� C���|)Db��*|�/S��>qi"VL�M�i
y���y9sL���	H�-O�Z����;)I��6]��J�Ш���_y��)�>x�����X��nϸ�@� ��p0o<.%2���VV��vTjh����2C6���>B���<�s�Z,�v�z�t*�ni�� S�]�9D6_�ޡ~6Y삇T�p4�W� ��� ��j.�N�p O�L�B�,�2P����4�� �?+��7-�Y��[~��>{7�G�,���&~�ʏ_/�V,2nR��F4��+��t��V��?(��G�x�lA��6R���ɼ�x��ʣ���m�Z�D��7L�gKy(>�9G�\��;s՟���3��I����Z���@m��!t�'V9JiK�\�e�~�I�)b��(R�xs�PS��Jه��2�NM�k!�u�y;��sh�C�NǸ�e�$ۅ�4U'ԣ�3c[��q��8��=���)E!Yj����1���g�4�lH��ʝݛxʄH�iXdx�d�-E�g��@q�%a�jԠ��+�V/�tJ���z7@��wt^
��3�����~:�cA���"D�C����o���R�Sj�|�|���Cx�Ё�����:��5w�t����L�[�����{��]_"'�O�v2�JM
���x��q��U�V}zb0�
�F���ݓǇKa�*4�3�3b9�(���f}���@��Xܝç�̕��J�����P��i�Ag]�1Z@�}sI��ӕ#6���f���~W�-0o���<���`�~Q��ͮ���ޓ�!6����`��{���B�T�	�ov�]Q{�D�����:\�>P<����)�(�Q� ��6�#u�a�L���:��"�R.�縧Ⱥyh�B;�g��G�R���k�E�֭/aB)��6v-�����g!�i�ѓ_T07b,2����龀�]V�17�}`���A�d@����;�܎:��+���4���fM(�cq�[`������Q��ڍ�P�$5{P)������ ;ś�*Zd�ȡ�b���5| ���<ζ��1yɩ�Fn�#�͛|���G�����e\صؕ�]�0�Q]Li�D�gwl�*�Η�a���U��ѱ���t�0Gs#���uDvN� {���g�g�ɰz�U���=Ls�5�0��}��`�1Fۗ�bf@�BE�����r1ܕ-���U�ĺ/?e����ge�b�d�@b������tWv��f=�EQ4��,����V$�|���v8�c/�`�؁�_��<�ݪ4G���
4����B4��H5���%yʃ;�&)u�,�:���F�q����a=��EM�Dt�ǩ�t�Ga�6mX�G�A�{�@,0g\�%Q�l| c;��f�`�W����#�W8��c6�S_�p�v��
��lHA�Lv����s�f�ۇ(\�z�[�^bc7��A��h�������P��Job�7_�Ke(����s��z,?����̏�L]H@� +��D�lY�*Op�0��հ0ܳ�V�i��]��.���I{�#�G�kq,�C�/�*Zެ�Ҋ�m�.�f=����2�ѩyV�?Uv��ªƪ�V0�Q@�j� H_'�w�4~/I�(��g�g6+�-��ZI"q�IפW~���������j��/��c�t\���&�\�7Џ������� �q^�A3�:�٘d��~���:J+ӣݿ�@5j�Ыݓ�moi��6Q�&z)���&CX�)M7 \����\�!�ǟu�Y��P��u�A�פ�[���n?���޻ے5�1���z�Y���8 #3r#7�J?�B�����
�M�'^�2[�a�@���ʞ0��3�W��r�W�f�?
3��+ܢ:7�����a�g�ܦ���ɫ��ylv����4�*!t;�w_Ǐ�8���9]���]�H�B���ATv�	����!�eYIgt)s(���iG�Ӯ="����W�a�Ȃo���%Q�!��4��*�P��2�?�/�`?{�پ߳�:y���պ��tM�n^}5��[re�3��ȢT�.��s�L9��K�'�t6����#h�������_��ڬٍC�R��"��P"�|�V�"�W6����Q���B[�4��;I���
��fw��#�\Cs����X���������>��f���A?�um�w���ϓ����9r'���N�i�ɶ�e!#���R6�U�a��2ƨP&^,J?P�8IK#y;m
�����{|XP1�h�'
)Hpp�R���I�Ct�l���hVm�\�Sd�j�+X�-�����C�����\���!#�t�����!�z=��.o&�poe���������Q?�F��{֑�A��)�=[#[��G�k���P˨x�
sD5�Rv��?Y�Ʈ�>��bO�=؁D%���Gu	�Wx�XK��Ϲ\��࿀U����Fvm�50%��K~@��<4���5!������oP�j+�3��P0(�6.Ҁ�JS�k]�Rq���w�;Jg���jQ��f�C5�ZZM��?������Te3|��Ώ
�;��|`�R�-��B�������hN�1u \W˕�7��op��sݾѿ�谏_���50�"��MD,����&3˝FqGȦx+��w�7P�A�ݼ4��c���m�%̲����ߚֹARk�'��[S�x�Y���t��H$ྸY��v��i��#[k�v�1�8�-����{��ʅ8mW�P�j�m�x�NY��q�I?�O��]�ƴq
�W���9��J�)�ǉ���*�t��
x+q���ۜxr$٭�gWˣŊ��a,8���A�����f�.y&4~+5��[�  `�~*Aݟ�p��f��]�)
�(����U�BV�L�]ƭ���/G��%�ҏ����'�b�[�����L���Q��M�\�<悄��|�m�)�Yp��q�
�;��{�p���i�)\!Rr`3�B�s,捑�n&g��!c=�̔�#�����:�P��3�Y�G�;t=��%"���Ϝ���gS{���w�|BS^=��U���r���Te=�
t�ة�J+����W��������2 1��!D2w��k4�Q�v%O2!l����5�	����70f����&.u�H����G ��>�����o>����*�Y�J%��QуIu���C��.�J{,)�~��]1k���f`r�_*�3�u�+
(KwiQ�b�/&Z���%��~�/�V �H����m7���FrKz��1\.��$��Ν@f��+��s(��C�[m'�d�.�ư�HkW�s.}����$s�e�;Z�R6�XG��1���>�����uu�p�����F(a�_0u�|h	�������� Eū&`�lm���#a�S�T5� [�x]W,Cֶev��Z���8vx�/��%	`�#I�w�#s/�EE�ᬘ��PvPf������� ��������Q6��C���B5�o�z��V?�p�\�C9�}�?�>�/��k���G��Jѭ��ƭB�E
s%	����P]��W�Ğ�|�Z}� 
��j��4����`�xG0�CP*��}/�5��
��%���j��Ӭ���7��4�<�5�������1����͉4ĸ�Va�	�M5�*�0e�*�:�g����p�#�����5�+��&`U�@�R_A�����:O�����9E;?3�y�{J�ULo ������ݬ
Kyׅk�+*�K*p ��J'V1�ɱ0-��.G�Z�7�w�b��F_q<�-:K��,��>^Ք����L�-�� �s
�I����*ס-6�d��g�&��c&���ׂ��r{�ܰ8����5b�T#<�V}�8	D�h=���_� #����*͋��Pj�t�@��EP(���z%g�F�/ҝ�5s�g*�%|���GV_Cث2��q��9Z߁�(�3�P���-����l�v:���u�Q��������sR7i�d��z�������� ���ݟf���V*)0���KcI��}s��rn� ����!����V�����U]��(>|��(���n��؅��"�;���0��y̌ѳ�ъ.�J�^�0E�K���d� g���,r!cD=���L�,�F�����ˬִZ�Ģ��G�Ҿ�͔v����Fy�v	"�m?Y+^�Ȍǽ������i����A��lE,.��-:�X��H�ˆ)�/+@��Zܗ0x[6e��<�7��(��E.��ȶkT�{y�,[0�(4�^�͖x�
>�[Zc[o�n9*�9�r@�Է�&dV&��/��V�n�����t\�0����>�Ox����܌.��/�_ڢB��9�յ��țUb��-2�8�Fj)im<��V~�P�n�$d�� �~��j.���0�:f�^9Ӫ�x�>��JFc>�
�|��"~L��t\]}�9=�! ���<p��,L��*�-��w;gW�%��Ń!9���fY��:����$��c¬��c|��&C?��I���&�|.[Ԕ���.��ш �踆�T~ϙؽ፿ Q2�'R 7<��KX*H*(�	X{��(�*�%�a�ɝ����ح����1���n `��-d�Ӵ��t&x�h</�F��A��������V�+�N`ߗ��׋�D���ߒox�F�]ŀ�s�4L.�
.��kXyɋ�#os;o	m����R*m�ء���&�&::���S''��9��x�dנ��{p^�k�l�\��DJ�E��@8�(*����m��y��Z����-����y��B/���@̉Ż�i0&%"�tl�4��"��(%Īh���Kuu¬��i��h�5�d�i>�:k�6fz�L�TR�R��Mr��3�q�?p������n�Uy�{��͝Y_�s��Z�sV��dpQbλش�\Au���f>���u�;D�H׿�L��5�(���2�#�5��[~��	+;B^��k��:�*�]���3\ǵ�a�$�qǂ�,��Q�	c��(�ځ��	�x���a�g��n��Ŗ��MH ia�Ut�0�m��8[�U��������s^������5��]z�� ����谭쌌��R܌��d6�W{%��٦%X]���Z,����S5.dO����0]teD����;��؈.�<e�P�R�YU|}�T�(z��(������2M}��rn�_57�@���q$Yb#�opg���Y�$1�4V�Yh��L���������������dQ�۝.ϐu�ݶ��I��$�[5��dJ��E.{��|2;9��-��S>��jd{9�N�O�ޫ�E����e���ܞ���K����+���T'����lM]������]���J�N�y"eX��rg��؅�F�P:����F�s*ѫtu5z�I�.�a�8�1)�M1�P$������{�>Lrlqi�z���^��o��?y����H�����RuX����>>.r�Ӊ� }��+�U"�I�C������J	x��M����>�R���a��K^�����/����m{��P������?�9h�[<���U��x>��c�~�v�?�8������0��ǔA�-�됲�TT���xhG!_IF�`M,�. %��
c��$'�1T�K���"8v@L�Yu�ЍSt���$�11��v8L��+;Yq`xö>�/�7�?�76�7�g�84�1����9�Y:�4g�,��A���J�F/Xw�YO�q����_�@��A��1�u}L�1����#�B�-�?��˭~�u\�+�gR޷/ք�|�U������`��7��ȝ��@�窅 F_�|���Y(vΝ�g�*��:2�@�%:�=
�S_�T\�e1�T�����B�$E8EO`���	xu�H���G;�	bn@TEc��r���yW͂�
n��J�����2&�����K�i���p�.b�V�eR,����/H���?��?�[Uo>��]S�O��z��(���B��`n��m��-r	}p��/8��yd	��ԕ,&�#&\��&[�g0ON]�H/��l��.dm�3q������z�4N$�'�ɪ���;��锗';_F���>�[�ʨ��1������Xb/�bhؘ��d��:���m�^��|z��������vt!���A���*l��0m��Rҭb=w^y�X�ϥ���A�D�f�?ʅ
vJ����+2Cy�=S9Ä&D�����f�����8�q=�� K�������>j��sq�Tm���?6�)Q7����t.y���a�a��KPh��=�z���JD_��#����:�1oQT=���]���4qX��5&G�k � ���w@WO�Z��9�N��h�f�Fm��B�n��}�{H�[�f��!�:�d]�A���x��S��Ђ6�U�4[�Cy���VO�>����/cV~M���@�7�Uy�I�uzUʝt'n`�� ���&`$]�v�XS'��*�'��mϥ�>>��.�r�^�PP�P�`̒�*=��KD�j�mf�h�U`F�TH��sP	�R�^�t���N"6h�z�毶�s��TB�� �&���|���.}v���D�7���i&)Ϙ�SI�2�&;��!Y��6�W�ӽ}��6Ӹ��a�x��n�e3
X�Ί��+�3/:��yÞ��9̸�����7��+�_�[�f׹G��U�KA�]|�(�T�.�#9l�B6g�IK��o6j��h�l�}�,_�RFp��b��t����h�٦7F���6���!Y>$f�,�?����� �}Ѵ�l��D//w?�;���3j��R�8�OG�l����)?����,�'�2�(Ɓ{�6�N^j��C5�f�]y���$��Qy�!���|�*H)�,u�i���D�E�N#a܅�c�o��Ҽ���X�4n���
 <�H��?�F{؊��i8)푅�*��h��lxqyp̮��?lZKuC/��[��V���'g؎�kA�G����';�4V��TE~��*��$;���1�0���}:-n��3�[$�\���6���k�Յд�a���ؕ�q����{>���;�A�閉bRC��3c`RI��ݎ�����C��n���/v�B���w^��@)���EK��:�ǖ��.OOKLL��t�e�K�2�H�����Ɖ�Y��G.�,}�P�5�|`3h�*pNϘ��K���#�W��.��î�i�cR(����y�}(i&C�s}�V-:��
=Sla� `�$(�-��T��3��~i����`pl�@�D����EJ�����3�Vç�q��R���;�*"�8��r�(��b�{��-�I�B)�]o�T�`��w9��<�9�|xi�&+g�T�\J���:q�r��|�޹��Tz
�qQ�i�C���$|�t
�:�9�����`��(��v6X$�i`w�p�������ݺ�[&�"d/�T}r�G�A;N?팞o_�
�IY|>�ϥ�7�m&'���'�7����@�������?�V>��E�%A:�f�F-���kY{bh�z�Pq����Mȯ�dl�˨C��c��ic��7lxl�.�Z!ݎ +�����"�$m�'��w��f���8��h��Yӣ�_u~����=2�
!�h�����dq��a���3�{Z�i>_G�5�h!�i���@ (��?^c<�W��d� �lL��U�?�/�/;����6�Ӊ����vP=�������X�����Lv�8bG	'�&K?�Q�g|�x$���� �Ck�dT2�ϜG�G��P�(2�
k�(�\�jLI�y5v*��1v�� �s#j(���5m������Ӵ�M���Ҳ9�%ș��b�t\��Oӛ�rn���i$IXcV���A\j����S�j�ߩm��Ӏa����bl�4�\���
��C�tu�d%H�i��v��v��-��/����Y�qj/������ ��?0P^ L|U7ܯ4t���7�=���#w�+ƶQF�,��/+(Q���/}+)°�)�?�(��ᴖ�(�M��;C>�	�
̟�*N�Z��# ,�Ϟ�6Δ
��u���� �~���ͨ�l���k7��Z�ywo�H&vj���n��cU�{�o�{�j�*�d|L�N��'��Zڠ1L�#U�4��j�sGұ�U�vRYS�0~D����H�s����s]����1�Ƽ3�����=I)��y�@�I%��}�E�:lH�_���-
X������+�<��tW7�0�����*cE{�GM,�A�\Α�y�2 ����H���]�]���/ƶ����%g�@T����&�#\��NX=A7ʾ�uC�{�v���G�<O�W<@Z��i�N�4�9K�dl�Wb���ߛKw�oi��{M��o24_%]W?@�+Ltw�e��A�&a�":r�)�!�v,�n�]��m��h8%e�C� �����{L����|�D6v��|�X�'�rt�Z�&��CõT�p�Mmg���K�K3.▗��z�L0�L��O9m:ۀ:�Cw3���<�W�H"A?d'���L���?�C`;���IK�u�c�z����*G���D�qޢ>�|��x~����jYe���!�UÏO�_-	���k<!,�܂�F!P�kY�$�1'��b���bQ3/��0\6�
�H� S�?�\�r� �[�G
�Es�Z$]��;���KO�>[�Is�F��zM��O�E���d:������kS\^�j��1��: ,-�V����I���OZ�dS%��8�(�֫eYY��������Tir���[�z����/� ��y�N�ǒ�����X�e)��XN�c��� .��0�������`��)����2��8?Q���	tk�e�$+��F34�p� ��KPW�:��M�*f�����.�'�G��I�',<#:�C����2�{�#R+��W�~���kl+�k8�[�QH_8Z+^��?�5b���/,(ϒۦ���iC��۩?+��HE� �1o.�I��IXP����o�Z���r9��t� (H��9r訋��ߩ��k�%iG勁�@rp�	m�:����,�{��=�"?]�\\�yTu2ʔ��Kf�P4�<k�xB��Wԝp���m���وZzG
wV��x��^'.r}�-A@���N�a�ݐP虏K`/�>�������>)p/��{�����c�UD���v�0�{��
ͻ��T���9����h���
3b�Mȏ�.���U��:��}�+���&@��y�V�kh��u�[<ɜ�Zfz
(+�M0�=%�\�;�1x����ڏ �׭�K� ���(F����kМ����C>��1�H�V˵�JMR1�֢s���l�:^�O7���C����a����+3Z� �gEF���7�ZX'4Љ���U�_kҤVǭ`ޓ���8���L���??tvY���"8&ϖW�9�l�
����+b���쐏F���<�����-����@�I�t��)�g��eNS	������B��Cg#����@�I�S�rB�] B&����`�V��(�2��(�.�tį����`�����=X������-��]��* �`�����I����si��Թ��~�6��Ǫ�p9u��#�6�,\W�f�����Ŕ�ZaC�X#�Mh��l��n���W��p��1Gt|E�ڕ*�B��S����6�0N�(�#� ��Ӛ�Q�+�M$τ!�}�<�PI�!�0��Q��5 Q�c6��\zz�[���,�m�1Fd�U�`w�pȞ�}�곾�1�L;[T�D�dv�N7m�jp̝�>S�gF�̳5�e��	8�ŀ��3����a8֎�Q+Z��Q�b�:�`֒܁�O�{���Q��%	6�`�M�����N-.�,�>�j��Q D8�fsPZ
��~-�fY���_4H)�E08�(n��d��p{wd�z0�Wbd*�#�Y�)�aH�Lğ���/zV���\���1I�G�Tq؁{e�`�}������\��������^M��[���,����`]���o-���������qRuZi!Z���=��F����ϡ(�^�y�`��v�����1��L9�z������Br����|82�� ����1���pH�Y�'է�j�.���mwyxn�����0f��_#����L Ԧ�ֳ�u�@7���~"X믬��-h��t�P��ɵťU>vN�%��>��\��j+�-=|��|�q�A:�
�~�U��6Ԋ�_Ba�>�D?���d,p��l���k�f��B����Ar\0�*�1�!Sr�������gU��ey���E�v	�:�<�vр��ޜNz�O���7�oŹ�t�������T��I��o|�R�^S6�|][�ml�[/\<�V�Ve@��?��v�*�T�%(��0v�Hy'��yfǚ�d�]j�Ìdt�l�-˝v�*
�(�#^������#��s Z=�v���"���/�׶�#)��I�NJ8��J�C�8�d�&L4*�܎��.���C˙������**���Z�(<�J9i�2�={ ={ށ��C�!�<&�"��;s"��׾��8}>�J���y���񙓫�*�cY�
�����ixN�%aI��U8ߊ��S�X�a��.��Te����hE΍��n���ȩ4$�K1�w����W�(6��UcL~i���ث\S������ �V-��,e\�Ŝî�a{���)�=IN��h7�I�ei�I�K�}.0`	? ������%(w�2nTm���p���n2�A��
W������D��/�e�:
L��0R��as�h��ӄ/R�g#&�b�/���g�r�)��+��
zG���JbKL#�4zu�����4D�n%ÌRc(�����)q�B��"���K����-�GR�B+���R�֗r�(w�/��[��LB�GAf�ܾ�_j�j�L>ZKݬT�\�%��J���R�y@�[A�Ƽ{o
(X�t��4B�5�7!����6�� 8�
x�r� ؅cf}?�p:�춚����֣�NW�ט��̂
��X#@D2�dL�����t���v���c���97��I1��&��<o�{�lKˢ0q6@^��u��`WT*���kU;��=�������v�|��4�hI�
�xF�Rj���nJ�{��"<��&mDL^����N7��ެ�'z�0Ir��R/tL���0e*Hp�"q�\O+������֑�*&�9�W׃� 	�so�;F�	�ɰ�Ft~,M��� 5D��o�m$W^��k�͹>e�䒆j;A�t�C<�&F�S@G4I���u$�;z�QM��#`
�x[��;�1˥�YQ4��'�y�����eg��RS�dNPzap �����5�N<q"�KNEx�dM��qK�M-��bq�[y��z�5D΄-D����C�Xrz��4��
#��9}�컬���o�`�����]�]:�v3�'x^$���A����$﬍C�%3�?S���w3��uD*���]���I�!x����M�����$�'�qAs��|��ƇH�0�[����/�Zm�����C�g����^6Eb/��؆>֗v`o�=;���u(u�V�_��1٤�]16Q�m ��]9~���e���~.�mX�e\Y���LR�۹�v"c��d���h(�	`��UG��K�v0w��SFpITm��~'̩���TCH���`��`c�]XC��J���۪���?�\�3��:}VܯfJ�?�4?�Z�*c�'�ΏII#��p�r$����N�p��@(v���@@hV��q�+{ �Q�����T�na����~�(���uΊ��X�
� �2d��O��ݗ�O ��Ϥ���ucUJ��+��cс�M���hbU���%�0W��0X^�M6�8�$-b|���;d�TB;�2*Lk`����F� d@ʜ�~��ԈP��v�0��$זMH�πoY�+�k?Π#�0m�c������jJ�m��AQܷC�%t�2�ܺ$���@&!{������QTlt|fyU�kB���t�N�֐��\�i\C� �ed�z)����N�kO�!�[ݱ����u"���)1��sB=����<	eFт��q�@~,/�&��BOƶ��V�i@L5�]���?3,:~��[Ś!SQ�h��A&����ꎊ�'k\m�BT�N�c�0��+m'���:�Z�a�#��䝊<����ԃ�/�!�9;���(�i�sd2�Nȓ�[��V9���'N"T�Ch.k�1�V��Fo�����*���M�����+k�ĳq��/^�����(����n!<F�B��%�a6WQ|�i�v�E�l��*I��jA�H��u𪐕���-�C�g5nEI�KD��-W�!v�Ʉ��@�O�Ń�-�_H�hs! �-?N�\�ohu4��[�m�=��D	�7���Va���D2��[-�$�z���� ���L�
��ֲ�w�	-O�Vr�޶��A�3�`��?SOoȿH1���n���rN�������������J�3�J变F��`P�#S�5�� ��s��ÕѶ\�/u����i���`�W���%��=l�{
<GpYA̓\Z�R'�A	�}晲r�v�3��ҷK�"���j�J�YtAܟ� {�G�I�Z����
�W�C�Ǽ�'�}y/����%[��	=�����ǽ�:-��x|	��x����� r�U�CQFrf!�;�9Z�U��1�!
,���uw.P�=���W��'+�ޢ�q����)���f ��c��[\섈N낯�h�z�~��sZm�ǥ�%(�$r���~�ĵ^��v��厚���ieh�I�K�w+k.�l�̐3�HI��%t!r�>t�5�훎�y�#�7Q�0�������?D2�VꪴG�R��kہc)>��r�<�Ҩ��M��J�3iֲm�{�s�-ڈ�T@��7��p����6\�+M�� 2�Fsvt^�����޻)�4I&@U�\og��M�*�&�W�FR,v�-��
��^�9��GZ��!��0&$��.vz�8Z�9�7�T��������&<I�T��Q�h��n��7��!+��]�T���G��v�}�D�ި����)ɚw��R:�sm9�.�
-.�"������KaKuM'�?��Tgut��B�p���Z���4���U�P�ԃ���$�h{�ŀ��1���,�?v�sC��4��eN qBƟI~����@%Jƞ�:�0�B��,�@0��͌!�+�h��Q��� y�O/!�q6C+oy���j���:x�V����u{v��$���.u'
4�����$�B�V�M>{��\��n)})�,���,o~2���.`�]<L�<r�6�zVN�f�.�I�*Ԓ�&�M���42:�"IO]:�H�!�_Zń�82�=��HrBk$�f`�Ԡ�eh�#���Dm(`�^jnU����<ތ�о`0Yo��?��N��SꖁX�;Y�Z31[�'�z��H���%�]8���� �$�?�tσ t���d��Ћ�6�H�'�A�j0����:̋��dt�P�h���h���"���|�s�;�����x�<<>/�䵿F�3��?���{&���[K!~d�c޺c��so�*�!��)Yk�L"#��a��o	d�/�Q8���פSu�����p?rR���A#����.<��+�ȷ<ヒK��g���F}�oVc"�^r�W �YΓ�V��"�8�6[,!q�d�K�j
����T7�6%�̡T�7n��Q�.Uw	2H����o�m<oF����Vjm&�� ޚ�n|Xq8��tITvY��s@��,�����cp0en���hi��Jh��F6�,5vn�}�Dv���A��4ځ�v+�qt�$����m�U���dK2�=Sc	Nx�'_��:/�-���s_l��G�&i����ɹ��4�6n>j�	�{97XF���9�6��M(1����x��;9W&�������I�{b��
��m4���ݯ��]A��%�qA(�>¾��L���@Ď�߾ŧ���'n�	����H'Ys���?}���|���.��=g*W���X�P�5���d����j_C͆�,�+�B��}Ȩ1��.7��m����t�s�C�&�ϸo2��X(�j�VH��>���0�\�9wP�4��ꢙ���ْb_wJy�7x�����iFJ����қT ���τݒ��HeXv_��� M��3���͆���+,�JK@T �t��$�O$�̹�yd)��&tu޿Zȗ�0�e�ĸ{x�������6
\�Q A'VG��%�d0�"&�2�ot﯇y�^���{����P]>
�ٯ�rŌ���F+��+	�<
E�.AB�u9�2;�v��('��'Pz@d�r�K_�ɣB�g�2}�)	PR�����[��$���
�IN+�I�k�ȝ¦y&0|�0��И�p=!�P�7��"-(�"Q���pB�&��q���0���NGw��VM|�`��]Ko\�eb�Jvp.��6~% ���AaV[��g�~��{eO�'��HS��_뫜�~�������o��蹿�Y2-��|F�@�<SO
�P.�|v��u�3�b�׆<J������#c+�R�[��W��C��k�>.TB0w�N_���fw{'}�2�@��"�߻�T�GLL��z_�����\b����w-u?�'���F�-��S��zʂ�`	j��� 
�V䬨�3΁,O{cMe;W,5�5Ai'g�Ş�d��u��ڎas�R�H�A��w�ų�s���I�E����?v&�'Aq��T��@=>�Y.���3�Q�c�l������Ƨ���F���I%Ddf�_�1�Zm<i��;$�j��LdK���{�K���2!֝�KE�K�����lӦ���>�f%:_��oʠ۩�bCm`_��Xmѐ���:P��( ���eR�-z�Q��t���yN��*$�V�;����ʗ:b��zx	�dz��}���B���x0 �ζ���Ɉ�q�,k��)�۳U��l`e]��]g���[�8ز�EV�e�}�|	lN�>L��5���ۘH���vL���9(?�m*�'2���I��!Cb�f�S#�̘ź���*��}�r I��)%�G��h�Xz���M�c�냖�w�#����P�=����'�pe�C�k�SHa�w��3�Y>�p�DjYsY�sc/Rfe�t�h��,m����hǗ�2m����eo���waIͮ��6��/ɡ���E�ށK��ϹpN��	
U��1�t�D.\�W��A�#`��O��Km]�.���ǐ���G�k�+&n�Z�<���c�%��S�3�]m�
�o��n�����r��9�'���n���g�4;p3Qۓ�"��x�>��*R���u��w'a���C��>�W:m�x�"����#�W�.�a@a0+u�<���M ���oT��A����T\sU�G��1 G�TԏL�;��(Y,u��<b_���g]��[�i�.W/�8�~?Q�#',nR)0�s������K�}V�O,�ӱ]��g�ՖLY;&�
04A8�3��9$�o��\d��I�e΢G*�3���H"�aD�݄��(1А�s�5u܏?\rՏ�D�p������
�Wq��s���f�ѨS���:5X�ѝ�3A�����氧��l��ɝ�~��{��}\WXS�b�_���2Y��<�h�v日�4�43.�flWb����!����_��}�s�Sy�knh�&F$��d���%.�W �d�%�,K��z�3��ʑI�XhtftӕM�^�������~%޳=~�^^�F�9�<FW"BYOK|�Jp���t�[�|P���p��R	ժ:l��4�%k���2��*�VB���(&������鮓����!�%朗
�rb�[�p����}Y$�:���i_B�}�ج
+�6M�?��A�6S�4�?�A)TgHqӃm;�0p��L%7�h+fޒ���*
�x��@} ��!�u_
�u��vee�w��ſ�֫ �}ԅ	�B��$Q���j���Lt�rjtx�Eȿ�L���^l� ��O�zW[y�}�
R<߉a��o������ǄŰh����h���|ިS�}E�}��sΎ�Q�Η���V�]���v6��s5�^:�GT��"����^`ADf�`vu�Ҩ�[��^����O{�(����@�6�^vm��o<�� F8�8M�r͍@���z��� ^M쌮#�s�;�oxo���Q��ê�VDm�n]��jd�ej�Q	�V5��\�WJ:=������Н�4�/*Fq`o�R?b�]sV��5�7b��V	�˽?�;M �h�h�5��1�Oetu�F㙳�"�)�?尤y3O�n�wz�u������B��5J}�g{:G��z|%��qH>��CQG�]c�>a.׹v�i�m�����:��:��=�͉N{��ف�d'{2�_w��Ƙ��6d�(�6��OF�4�mF��X��j�q�˂�-u�ś��6iXb3�N�Y3���f�