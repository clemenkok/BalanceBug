��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�F���U�C��SC��63�Qg��ͼ��F
c��ô�T$ ��i�s�c��F�����#�gF�K#�UL�b@�����;���Aբ��p��|��X�了�z$M�zu��A�s��N_MIm�/,3�z�i��,��3��K�z�Ѯ���Zׁ�$ ����R�׻�h���J��f�|Ck��ݟ&������o4M^e8�7���q����OXh �i�� c�[�[�>2�ZDʻN���:��Z�ԡy�#�
�2M��nI6��'�ՠ� 6�6b��E9���s��rWpzG��ݐ�I��7�,���,�:��O͡��i�CI���b����M_ �{c��t�͠'��M������7�=���A�԰'�2(��'= sI�#�t��tcq��s\T<azĈ/�ϐ�Ӻ��x��x��5���-�n����.� ���x��Cј�^�ɏu�#�$��q4� ~�+�dUd�q��9�Fb�4�}�_,2r�o�;?�&N'��I+�2��Z��Z��kt�*qm��k�׶�iǏq�vx�Ё��_�qI��{Mh�"6xm��@��Z3�v�����*��VU�@��!N��R�=�gaV	"v��:P�F���o��pׅ�$J$�i�&LN��/wmX��=ǭ�vM�ɥ�Ib���ߖ7�P���'U%�ſy�b�0�`B�{��ߠ���$�L�,��{i��n������\�z�R뗼��������Kk��u,�yn���ד<ᷤ�L�m͸���}O�3�fh��H3N׵�c6���9t�_�e���$
�-�����c|�V�B�M�8|�@q��G�>��m!��^0^����[9/r�yAn�g���߸ϵ�{T����X�ah��K�� �ʧQi��9/VCK�=TAf+f�g1�E�����﫷���Y�e�X+�(�A���$%#Y�f���pN�l��y䬑G�_P��Ú�.C�ɐ]ٷ���5�����]jr]03���a=\�y�3�L���~1a��k7��Ad�M�{�rX��֌�D�n���c��/7��y��P,�O��
W���fJ�L%��^G�K�[��?QM�WC^��grEŃ�FR�U��ah���3/�}@�6�\������UC�c/=gqJ��n�O%O}�����~ǋ�°�`P������oӢ���Naj���������2ZK��L�s��+?���C���=��0EvgϕѨ����Ş��r�0�YF��5��~��q�T��A��n�]�o7]w��F�n����A��(�sb��6Vw�N���Ӈn���-O��馝�S�	Rd�A��vs�X<�ܰO��"M :M �Z��s�]Ǹo�c4?ޛKS2���7KZ ꬽ�Io��<�^�\{��fH:Ѝ~�F�4�S��H�r2���O]u��6�v[�;.Ӿ(@'[]Z�{1TBłp
D�=��{����]���OD9>_�K6�����} �>������V��GD�%(dJ.��X�kO�(���2_����ox�(� �_��o� ��H}C��,}����߀�����ɹ*���[�ͣ��k�M+҈�:C� �`��GH���v�;����^D�O<�~��Yp�1?0��[���C�w�(����X��C����Ii��\�gP���.9a�di�a*�^ޞ�Yn��۞��l��b�����gL{?���&�YCc�6cZF��*���c�A�<�D/ZU�Ĉ'2� (\�$����=.��}H�vA��(��������͝;�Vv2|�0\���^[�Vp��0i�|����ɘ��(����7�t�����߈W�jK��ae�ܵ�Q����Om�K5k��D����+�B���([=��4�<26���YH�݇�{��{����q7B�b<�wM���b
V7��"��ڣ���%г�T�b���a��?x򗍷�%�n��[�����&B\G`�B�,s{<Z�����{�gl�f�u��(�*su����A�� 'Q�塅�۞�g�5��$@�pb�t��Y0��Q��һ���q���O?�c���6�Lǈ�շoQUr��.'���#?�?��qe�Nr��ڪ���m/D��f�?�i�&k����[���x.]�|���?�\/{
���SÇ��E��Ն���TC1��-�,?�(v��]�q���ԏ|�"�a;�Q�ǎv��6�u�Y��0kl���\����G���U>X����W���w°VD�Mw�����R��E���,.K>�(�(�h��$Hb��)����Ǎ=�&K!��������L�Ë�����Zilfn]Py}M�!G�ߡ�Nw�p+i�Bzf�5fi�f�bq��	Lih3я��Y%#;�A�����q�yz�Ƒ�*�� ��-J_8���g���v�>I賢l�R�<�P9�,��ALPh9a+
>���h�j�z��O�h�	��+�( ��+,���~9uG��&z��oipU!�r}�����0-��8	����g'��|ڨS�L�x�i$"�Gcgm|28�NE�&�9|+���삚�o�_�;.C+�	g�e�5ۑ�p�P������O,��kD-n(ƒ]]3E� ��]��rvB�t�7�q�ºi�K�2,@1��IŽ|G�7�:�A]D0��b{�-��_ӝM����l-]�{<�o��Z�[�;PNz*R?���	��ztJ|)��_ '"��1���0k$m<��k��"\K���ʷO�%�@H���ς$�4�x�S���"��:�}� !��У�Q����.VH2�e�@��1~����rw�2*j��mPX`�n�����u#�m.�Hݡ��j �u�J�ã�};*�X�b{\������}�s�.���O�"|7�@p�N����~ta�l6�ƅ��R	�u./z��!;�#L�-OboG�R�&���'��E^�D5ƉE�L��zK���2z,."/����!O�B|Ӄ�_j�Kp�������iMI:~.4w��Ngdܱ�O"l)�f�>�6���%ਟ\3G���!�x:�`c��겘��R&>`�[���g' �tʉ̛�h������_��Z�HV\�h�-��`?�S� @�����Na���@T�c̬�a��a�ޙ����+1E�,c�c��1t�Ó�|��Y�?�%5�&/�]�ޥ'#�#�D:z-��Ŋ��|>�br2�C_P-�i}��&��+h"�e�D!���*���{�����2{1U��B��+5�u<��3%�7F+�{�yI4�Q�N�Ʈ��(D��	ߑ��]�O��ܗ��)Z�36X��v;B��0^��;������ �0�ۧ�l�	��>5݅RN:��h��}��c8��ZxV�Jz5=��pmA����n}�t�s6�[@���с�M��������DѨ_H�K�n2q��;z*.��%]�UK�s:��@�\U'4�'\�`|����9A'I��Z'���/�1���wB������R,9u�45� ����I����yE���vMM0G>�5�f������;��i�RH��Ί�+��#�h��Ir͟�0Y���7����}�'t�3f��Q$/��d�'6����덁ˮ��|��L/��'��6-a�{ݳ�/��R�ˈu�����sk��Y=����m2/�/�f_��Q	�=0/�,�A�/��2$ի f�]�$�_���z�F�!���<*����J�س}�K	_GcM
>6Y�F^�O%��_�P���o�}���`����y�	!�*����G�oi��gBCg�Y�ו�zW��=yt�eud�\]L�z!�aL^$ ���ѷeHy�Vі�QdƧ���
��r>�.�Ȁ8U�]	p2��]:�70e��aUC�j�)�_0�}������	0>��: KB�G���"Hވk'�g/��I�_�u95ڽ��л�^B�f�W��]�A��1't����+%6�L����N��JI�x�>iX3:�_�U0���ә-=���`�n����p�� �ۺI�#r��H�A�����m_Mф��E@�������db�����	�0Tz<�	��J�?�ŉb2�x,̰B�(/��
���O	��n2��D.�@'	���n�������RT3�ԗ��mp��@q~��Yh��s(R{�#�&�4����i�m2?oPh �ҴX`�̠�ȫ#�~�}�.�����֑����;��F�cf��E6�ݵ��h����wޜQy�CGA����>�Kas̛ͅ-�Fa�T��q:~2R�N<��AO�N׫ҪaQ�(8|Y��:m��Q z���V]m��eC!OW4R0{}�U[�\8ٺ�;�L(eOX*NIq[�m2�q�-K7K�c��ר�M�vv\Y��!�G/��X?5SЭۏ����a� &q|��z���J�d�M�F�����ڲ�(������]�M�P�m�,)^�����,��Y؃N�G�ƅ�q�������H��a�J����#��(e�n�X����I��H�,p�Bד�N�j�����i_��u�lW�|��A�#���ѝ.&�F�J둇R�1���$(�x�O�c�A�A�b�ڪ�B$�Bk�?%����o} �����p���1�RC�f���W�/�Q����	��	�3�}�9�e���=&�5����ײ����f@���p�u�.R�O�o|�>�[^��De�r��ʅ���f����t4srQ��vo����U�8%w�!x�"�O�0������D�S�V��.�e)�:���\����/Zȧ���<��@����Ϣ%}G��s�?Ig-71e������U��	0���Y�̔f�<ȩ��N�M�ŀ�'����9�΍���g� �-�2f-W�K�w_3�� ����%��{�,䖪j�;]��+ϲ>�̯�p�A�#|�5��=� '^��Bh�a��)x_�"|�~��<*�2�Z��e������<��Pz�4m�`���Q�6��O�D�W)��ٱ��W�VM;�Wf�q��PG�HUmK��Z%lF��Y�Ok�U��[�^ɤ�k�xk��V��d��n�p	�Gt%��p�0�z��'��8��-A����^��J��D�N݊�{�oz��\Q%BH�������c�^�ur ��4KԀ%Uھt�o�O�(g ����n�� �%���0�L�l{��Brzj���)���1��*�?T@p}��Ìdz�h�X}��������b@���S7Fj�Xw����$x�`��?�X�/'�j�P�^��
^��Le�`��M�n�{�M5�[΂8����#�Q�u���P�3򊢺�����C9$a��u-��u��<ܮ1A�YM<��i�����F=]�PG��c��9�huzm��C������C9�]r&���U�ʲ��6��v� �e�Y-Ht�q;M�c�`��m���&;�������A��Z:���8����$�M;�7ܽ�Ӫ�lhg!)���vZ����{*���o��b8E��R�]���c��jن��g��T�h��� Q���FʎW��~C�p��U`�B{��ֈ�җ5!�b�h�8e�ɳbkRҬ���1���Y������4LZ� +���0}���6~��>
�+���rҕ�H3?�j�yJ��w�{�{H.�E�t��L�[r��#��L�D&�[�E+P.�Ri��Ts_L����@$�Z�d�����fd�0�;�tjד�@�]	j�척vw�ExNL0����g�ya��o�pc$9��۶&=wk�쀢�Pv
��Q��5�@� ��~����O,��,��@i#������J��4V`!����H	�-�ѕK��"ݓ��y��]=0�:�קE){��ۛs�����u�M]XW��g�4 
1� �zh�R�-mw�b�8}��օ�k�A���M֢,� �8�#��%���ˋ �-����=gN�:Sz ޠ�����Lq�(�cղ�@m��HdC�J��G
cGrk σ��K��4���
�l�~,��9�V���!(@�F6LM���H�ϸ��1C�Gx��1�ɱ[���A�(�:����(���u���؁nGL�1w0r�	 �����Ҩ#-ÒyXN_u[���ih+5qJp���BaNL+�z� G��=	�KL0�`��R�+s�QvV���-{��60vafɪ�<z����`�P��_$�E�׮�PO��|ԃRR�
��������z|�>��3�jE���?x�]ST�4����E��ǱQ��y�2J��y^1ί·��?�H�~�_�p�C��'��>]�z.n�XP���P��:MZ�ߵ;N�s����]�
����&̬\�\$)��?;��� Y`=^�Г0៱u��2�y��S��NX%���#O�����������c�)�Y��l��@�����\�<V��=2�����@�I��r�_S�&�@7��r�Ǳ�M��A9[̀���K�������E�Ư*�e�dN��cG*M����4�"ߵ	��~:����l����䮩�d�_�ɉ�YH�p�k����<�:8!S��<��,��sP�iLA:꺚�a�� !��.�=��JN��<�	���K#�b�Zo �哫YTۂdM!���U�]9vi~;ZD	�n�Ҹg�c>����Q��C����d�`�w�Kq�]AF��(�rm�B�B)��PE��/�����jd�[��~\1[o��n��{����\�����XX{Ӛ�s�hW��ptM)!Tt&%)z�@C��� u&��m���Y
�Y�P\>ɉ29��{�y�ϵ�ֿ�lǕ��&I�D�"GK����R3Q�ꄆz5o`�܌%�D��8(&T��o
��*:5	L��.��ص���?��%edXV?(Y����lF���aS����?�H7�D�Ʋ?̺h�d���������T�����`���c��TCX?Q)�e��!��m�;wߣ
8��_�جܖ��XH�ǧ���q�5\e�T?����Rxx�^-�������Qz�wxj�Q�UdOG<+V�2�N�D�,f��̲�Wg�l7!+ʆ��:ǰ}��R�$j�Ҏ�{u\�l��(�~���D��)C�4����d�J�K����	GR�yJ�rt�F��_ ��!|�]�4l�7KX�(eV�-���mč������zd�__tN��3����#��3��~����#���>��pQ�hp�}c\ 7-��0���i��	���ʍ&ӸL}踀>�p�왱[��.�wxa�$?[f�Ez%@/�y[��bw@�P��zÇZ1�'
tQ��,�Z���/ʫ��-��e)��c���P�[}����A�*XV{��<�р��Tj�gD� C�R�������8ّ�\2] .qD��]/R��I��L
���hb��#m)�}$�+i�~��ۃ�v�u�	_^���b��-���]=,	��G>���q�g	�fI���j	���E��_���
�/���V8��Ij����@>�꾃�`|.�	��nt�P�L��yxR�C�u��^5΄�&��;��DA�����I�H�=zU����V�!�(1y5� �%-���|����#�V0�a�/<��X5�1g���c/��K���'�k��n�S\��tY�_�����TRϘe1aj=/.H�7^|�*�����i���	�1�I\���79�f�	��[dq��U�G}Дkan2H1� ��6z�w��e/Wi��q������(-��睒IO�����Y���"��;��z�A�91ub��< �|"�삝�����	Ƨ���K8�$١��8�}hF_!����	��4�Da�{Lx�5DC%�	N�b�8݁D�u�{��~ �NT�&��/xd#�J�qQ����ST,��
�r�t��8N#�&&�f��o-]�����j�*/IƮ���&# E�T���s�L�e�j�眾�/�hGCe��+�d2a�}K����k
1w텵/[C��-�٩��3i�A/vgI���4��_���MI�Y��=����>=O�/���qr�e����$*x�����;SAzv���
����O�~ȯk?�_����7T3��r>&z�v�ڔHf��GW�#�W�����.i�RbRRE����$
�`�:�l��&�]�����m-�G'�Q��3$C�H�"E���}�ޯ.��"�O�2Gs�Ol-W�ؽ�S�Rm�p�����?X"!ڽ�
T_���� �MY���*�A! ��E�U~�|������<B)�N"�c��fA�r����	6^DXzbSf5X<�(�QWɂl"�y�,��Si$j�&���٪��5�z��6�V���_ls���������}��fz�eW\f7|�������@h��p�]�g�Â�[��n���=�]Ԡ�^����z}�$���E*]:I5o�aNO�m�闘�����0i/̈́���E��`��v�������z�I%�� ��c�j�XeͿ��MO�`�bc&$�� (Ǐ�v�^n �{�����v����ֵS�r�����I\��^.zr�'l��G!q�3����5�|w��j�����V���4r�'��f�]�d��T�7�./�f;f|��~�G�'�SƶV
�~�h�Yebs.p>]�Zr;9��/\��{q�Pb��8��Eo�9ӈ9l��
����-;�������~�����)�ę�þ�b����fp7�2�y#盹Y[vVJ���A�
��������N����@�2^`�նJ�� �J��v�D�s��E��%"L�2+��Ĥ��ɼZ�$�pl��ګW>��9�fr�O'^�i���Г�<�h�<��N�#p�*a��A�3ei~�Y�2���Ym�ft#R�t��S��n`��c|��xW����oȗ�-%���ט���3j�8���\o@/�/eMw� ��c+qkq������c�Ne,���D;�čO���r����Q�"� 0�y�(�ӑ!�rw�h��T�5��:�11oY1K:�ů������u6-^���pUH������ *HA��Ȳo�J�meA�|X�!5�
���U� 1�앙%$�P���=��U��x��Q@����=z
�6����XUu������[�����́lJ��3��3M��͠�bFk7���(���>�� �Dt�q�J\O.]Qh�f ��ذ�~�m�A��Ñ4=4',�+$�t'�Z���9�ݫ
H�E�C표5�=El(D�Lx:��YCë�_F�~:`{Q�O)��,���c�DG��ъ��Ŭ	�V�#9��C}�N�+�ؚ�L�k���}��5�
f�;��`��1nqCN߶0:)�YJ��ogPZ��#��ZB&"ֺ5�`G��
���kޓ�%P�s���CFI�22�!��<v�2k��{c�ZgB�(�r,)yٝX�ō����O�����R#���Tp�'BO:+2��~��U�_rr�6�����v�|:V�x�"�冄�=u����#еr���NF8�&a�)+�'����A갸��=Y�E���\�s�J�*_S"	e4'ǎ���H&���R�Q�>�����H/!�aO�N0��w�L,7�z�ɯ�U��)��s�p��&�T:x)`�1�ܛ��_�gK��6�s~Q6x�|2Ǎ�ڡt*ĴMju�s��e
��� ��`�i���Ճ��a%�er�(hf֛_��q��������ʠ*�n�	�F-��ly����P/_�s���������hf���JA�~��b�g�QSS���.>�� �=5"�ڮ�
��.�7���[+w����=���f�Mhv	:��d �ڠ��{��ij�;E��*/M��:��a�:"�7pS�E�!�;�xL�0N�ߢ�����?�&�_��n��˦z�s�L.Z��g����~�e9�|)��/��:�@��a�!����C�;OC�	��F	�7j�׎V��N	UR���B�$IV�Y��x�H&m�U`���w�f��6+v�c���F�����N�au:�x0��'��2kG�#L��O[���M(Ej��Ha�:D�i��)#n|�|���K�t������jȳ��&�(݀#�^��A�x�*��+���O��B��EV�Ñ����Ҁ����d���a0��DT���s�M�aj!1�T��\K�kpr�C�⽑BK�L��o�06�}�̹gg�{|z8�
�|]�ET�?E�bP;]V�D�޲9�n���%��2�Z�7E$�c�c�}��d��_;�Uru�&#�-0q5���ށ�sL$c7�F����T`���Ug��A�{�aA3^N�.!���f�8�c�B���;��.દ�!.��������i�oﺬD��
<�w�\>Ǻ�}XË����� J��o���討����۫q>�g����nЇx2D��Mtuc�X���L}3��t&��R@�F�}��?�;^�. $ýVS}г�_�i*����sS�����7���.@.���0�ခ�I%a}��X����n������+b 6u�V���lM��$4��۪�{k��c��~� wˎ�[N�w��\��h����>�$~IT�H� �i���Y��o�G�� �����%�zS��|&��z���lt�Y�������%}����zC��/��'_o_]W�p^;L��JϦ@���e(����
I	��1������g��z��z��:�-��5H�ȭ�A8�"̆����\�ο���?�>t�DӔ2���lg8�0.R�.f'*���s/0���]G�ۢ�Bxr��8��(a�u+�Am<��O�Ѕ�b���`Z����T,JQ�J,	�H�b�Z_���hJ���GG�+�Dğ5��y���N��'�G��R�t���M��z hz��&��'_�G�2
T�^��=��Rq����^۽�U;��R��_�hS�/�"H(=���s>BǶcR���y�Z��A���=l,��Nt��sPK�\�ؚ�/jH���y����`�cG��;�/�c��_����p.��c�_}w����"�k+����-]ĹQ�k��}�����9!�3�7�d���+�[����_��Vvgr��^"�r�,�pO���3��K�3w݀3v�`*�7��=�u����7�d��U�Q�J輧&bA|5�'�NG!{%�]J�J��#Mq.aѪ�?p$J�@ɘ�ړ���I��}��	�b�����M�2@�s�Qk@�d���N�;$1��,�,΅�V7W3���/�����kZ�֩6i�8�2��n4��v���۰mʦ�����D�'�*���&�If����w@�l!�s��NR��d�%!��uUp�a��斀P����3��`���'n��ă��`�`��x�`�ʴ�� c��0����Hv��9���l�BW���S=�Ǭ�G�m� �)5��4��ĕ��6������\J�M�b^3�VC����o��Qe�@��V�( ���Pd�<�Oυ�"	��{zPJ�@f5H��[�i��*~T[�,#V�iA��6$����!FľL���yg��=�LN�?Y¶y4���J�<66?>'&���F@�p�@�w׭"��9�ٳU��i�w�71�Dwp�̀��.'� @oًZ]�0§UM#x���X���/y|�I��򉗧~�c�U�O��Y�,$\I�o߬�"6��'�[[ۄ�gʰ�x���ɬ�ƫ�%��sU1�Mq,����E������m�|�{'�?'���E@��@��湣���t���<�l�u�W�����`�΁t���k0|��4]|���@�M9|Wq�"�U&6����@I�{@|���|��@s�WI.mИhC&�W �B�/ G]��!*n��W�����L���\ �0#�/�0��lY>��cM.����Oe����7�� �d���?��Ï�R�3F�XRo�I���$N�'pX���qot@H�y{���a�k���M��kc�pu�ux�o,��hBFN�Қc@�4˃�V�H+Ӟ�C��]Iv$ǖ��'�`X�:�L8��D���i�Avbkud��s��Z��k��}#$$�
�X��W��	A���)�m�r���[�Y�A��>Q����,��Y�$I�?6��������0~��r�Ty�;����� �JO���^�61I���ʎM�?d�i�*P�{���eIO{H%ԇҌ�]����Za=�T:/��cר��w!4�d����"�.;?�D�ԑ�0f�&�`Q�v���w�E�i��i�o%�E�����9r��JM��5hep��a�н��1�)���?���$O�qkɥj6D�	{9�1S$u8j��q !Oqf�*N�|%T�����9K�b��As�$��#j�aS�D`G�=�
���&��2�����DM��.$�+�Q�B��f�Ձ�\��4����d��N����������Tצ���!/�L+�5.�0��Y�S�gC�����T�	���	][p�ʖ��K�Ta� 0��;�E�,SS��
���+du[�p�@V�ӹ�k>�W\ �tm�:�n#4O���SnT(���n�г�8/�<�25�:x�r7{E.�j�Q�B��ᦑG0ӻ�=<�`�f�6�Jx�8m�UP��S;R��)���\������G2S�G�������
\����m�)hZJ"��b��QB��`v�鍀i�vi��Ǧ�F��?Dj���V���4�ƿ���E8ޝu�Iz��&�V8���M8(���n�>K4q`�F��9��/g��:G�)ޒw��=N�L����*}�h�"Dr)�t���Gk��~Q"�  :{l?y�H�G���TX,WU�y���l	"5%�d���p�ЭwB���oVŹ�2u��E�	0����x�� 1��hB���eS��s܆�.@�_v�(��l0�|쬍M�2�׈�u�TX�0J�p�����Ywh�e�n�&Q�m�4��[�(�~�d]>��y��	^�/x���o$���Z���޺�a�W.\��qn��}4��֔���������w�i�CyU��g����nn2<�L(�i�?juR�_�(]Ė�D�q~���9�o|��FE̓��W�v(|�F�� K����~� ռ��G�AiÆ��8y����9����W�*V��B�tq�qP0���7�U�i�-Aɂ�Vl��%M\z<Ѐ���vM��x1z�Ҥ�t2o�9�a�|;ɶd� =� �|RI2����^���>�U!E�*�nms����f��)��N�B�}�l�bb�E�b�-��A�����gӝo�d����!�����*�~�|U׹�����e�C�Nk��<�=� �gh_'�͋_��+9Z��� �ުa�I��*�~�߾�6�Z9�:?#���gk��1l+z���_�nȴ�������RWP�}t����v�:-��B����M���R�[S���	�UU�D��'@QS;/��%�e!���b��b	���L�����V8:T���W7��}�=V\S))J���W_��o��M{j� r=c�ul�G�ى`�{(J�Ҭ�[��W~&o������2�P9����ľ�_�^���K�1"[����X���)A���+E� 5���f.Ze�P� ��c?475�"��I2����@5���+�ʴ�uF4���.����I�g�X���u-*�
C���؍�7��mF�s�\c8�����N������ә�ڣ5(��қ���������V��hj�oz�ΜtB�gbe����̻ՄT�����SW"C��0��T�vw^!��r�W�+ة�ko<{IhZ���t�4(�(8I@��wYZ&���:ST�Nb��4�������ƫ��(�`7��:�R�j��g�a�Z@)FƑ�-��{���Pu�uKU��Τ�q��O��|���)UMz�����ʳz�6E��*��pH�wq!���m8��16����Q<k[��i��� �4�T��m":(h��X�UUg�3�Jvr�=��v�L�ZjG �έr=v<�=t����XB�]�A���kEТ����<�]$����:�x|w�+��e+��§t#�����t��OMU���vF��lnh��o��E��J�����\o:L�L��$�7�ZƬ��<��O����oC�\��m�C�kξS���q�^�����q���c�ZE��o���k�t����e�%�Y[�5��L�)}�Hp�1��k��
ӟ|�
H���n��I������`�bE�X����d��k��Cطr���N#���<��9�Gb%�Y�+i��MsZM��I�江�O���$,n�S����0�R½B���Ԣ�I�pe{�͚��
���z�.1� ���kl�a8��QT���/w�O�#�
��Y:���DF���x/29{%�#�ǐy�)9����U�`t���#g�y�c�����`YR,,�m�V���yX�W@C�#c�*���r���	����O��Eo��&��l
}k� "�LT[�,��P���ϫ���p�v�����)��dz���+���Y�GD�.4̝`}y�3�����/F��1:xT9s���Έ��c�����ƶ�,��C/=� �"��Fi#p�V�k���k�Zu�����MN����|�Q_�H���מg-�S������F��-����O�z�i�י~K�Gioy0>��K�c��2j�� ]��d!�nB�=زUGL�{U���	M�8��;�t��%��u�H��Z�Y&�'�~vuT�l�l_��ۃ���x9�Rm�J,�״jJ��$��������+%�]3���E��;�>��\�(i�(�e�*#���[EvCʱ:�@�଄�:���a���0������Q���K�a�Ҵ�Ф��*����A?N���t�SX���)��A#��U*���n��O\
�CJ�����>�,��mr��->���4�Ձ�;h�-j��{�f���\����#���]2?�6w-}�g�m�D�Mا�]M�-l�Bo���M�8��#��AF�$Z0�<�E�Z�u�&}��Ky�N�YH����w��{�;��?:2Q�o��(��*6�t�E�x5��gq���]�e$�ͫ����9��P����f����r��s�v��>�#�*�_��P��X��{���.}��|�*K�0/���0�,�=����"@�([Q^)<7(��2��}:�����~��z��,/��h?@����seb�N(�I�no��_���{��Z�J����L���Ů����s���/qB.�����:�Fv��c̵ݩY��T��+��;���F� ���jVH��;u����"�a����5�I�`>q���}��O��9�5eH]�/��l�2>(|�I���:LsU}(�*m���0Hq�܍jaKuWO(�kQUW��V��Ї䲖el������pXLi�*ڪ:V�w�v�&91��GY
���a/k��̧E���~p�*e.Դ'3s�ߡ�����A��@�b����a8؎żR�/���^�r�@��`���MsAW��V��K[onX����|� ��:Dh��INIS �9�Yif���Ej�_�KL�"`潥�G=|v�޶�t?�r��� �9���	���ѣ�(^�Ȉ
�*7�����ǒsA�[	n����Ǌ�+�0>�+Q-|OQf18��3�Ι�-�[n}dh=������)�h�a8*����+�2#ITࠩ�N�̊7sK�6ʬ��S٠�d��r��U�q�ft����O���J4�W�P���{=���7��f�!cu�&M8]�>͆z��N�[��f���0�S�Bpv�����+&�G���2���]��%*�ڈ+Z;̰*t0}6�[b%��A�j��CR�:6�[�U]CőA!�,EM>�]NmyW�$9�P�W��Qڶ��Q��~���o] �P��>2_xkt&b�F�1�('"𽿎�D$x�Z�J����x� iP�J-.��?�[�9��V�#�Y��(CK�[>b1}YK�
${�B�F�n<��P��EKL�T��5�~����V��y؆��ں,�2qy>iM���.�F���|{ƌK�����@L���%,ڹ������"�pċ���T�2dg�!N����-9m���~�/U)�G���t`�RϡѸ,B��`_��?7 .�O��é�;�p#M�m)�D�O�����7)�<�{����I�������T&�c���F��>��f�����������]Y��GY�E���d/�U'�δ�;�E���pO���Q�?�d�?�?�<��o:9���< j ��rR�8k3o��D�\X�oM��
�s	���/;Jo%�q�`*1o:{�{2�{x�-�T:h�C�>7������mc�C;-��Ck�?U#Q"��{�$�l��#͈��N/�Nˊ8]�C�O'�y¼oA�`�ߦ&a�0Nbh�ғ��pA`�=�"�e�Z���kzT��h�Ur��u��#�@c c966��C��S�d7���~a.�;��y�:z{�3zK)���G7���ui�sgi�����Nu�k��/�n?����S��q9�2D�I�Gոp)��v~6���f ,�\0����v����ŝj� C���p��V��%��T9�"Jp[��L����>�CI�\PL��A�5C�|j� u,��kO^��1M�&r&+�3H�W�0���ˇH����"�c��N�K��mJ�9�C��f�2]#5�c�ޞ�v>9���/����l<6 �z�[���#�3
���w/����2�I7�����OV��ћ�&%�7��SV�윮����{�)��lAE�)×��R�]�!���K�¥q�~��\EA[�*]n
���IKw�_�'# dM�7Ei ;��O��`l���Z;|��O��T��0�t�e�^���u��&kR��7��31m`�.�q�CBȩQ���C{����͙�&��1E�e�1�>ҟT�y`�:�T1�n�4��Q����.%�_�K���QH�]������Nv޴��-Z�Tn.s���������qZ�V�����$!eSh�$�eRy�sk_I�`U��Uo#�!���j<�FWw����"E�	��E?C���P|��\�Ҟ�4v���TO��J�tЂ���i�Vh�oUS�{E$����v�c�k� �ɿ(�]L�^�b�3lg���XM�C�?�	�^(�NQ8񬷎z�P�r����*+�d�;@�v�XTr-�<�z~�PB�Y<Ǚ�q�2�-����t����#ʍ��T����!Mh;�m���JB`�[��D�P<�ڥqn�*����{�����o#��@*\�l�K!y�\�CQ�63.)^��}-NVtHщ*����=�u�a9�_ó9r��ؗQ[˨0��T�*�u��n��"�0I��`w�u0��n� Fg�Kχ��V��F[H�L���}�au�s�{{�T��ޟ���4TDn�w��$	}n0v��9����4��D]�p�XO&2È���(I��/���Ƅ���L��� �K���n~�"��R�=�IJ���Nzʄ���wm 2S����T�:
�Xb�gq�sn1��&�������0�����N8n��A�'W;�R
��S�p�Oo�
9/���yx8#֭��S%�'$V�S��˾�P@�3�h�j�4u")�GϺ��N�)�;�)+29���>Y�~r�w�$�:rU�w���J,AQ�s�N|���TK$��
1��'�ZB���$���T~�X�z�N�a}���	�j߇����]H���CʩHs�!��$�h3�mŬ�c~��Ù�@�4L��Ȓ�z�0��m蠃�o�i*|r�@ ��q�_[��ݑ�Ӣ����?VZ����v�i�O�i��Dx"϶?� ���k:V���4���]�$�-e#�"E�hjU1����T�`[����6�'_qZ]i�ܯ�t�DT~q�	'D��[��C|���W��+�n&fE��3�������#��0vw���?X�:���"|�$]I#����+�H̨���ٮ�R0�_ks<Qr��f7p��|����#�}���ռ�1�E��cB�h�����\�����|����s����%Ã�O�ϑ1Np���œIb���P-�*��pu9�ʵq���)����Fj֎�r�V�=��X5c�j"6VV����+�;��ޙ��P}H�k"}���vj�3�,F�-����t�7UD�C8�������[C�,�s�=$��y4��zu/��#�S�t2��U�$�²�=��J^ϙ���yU���-(���_�	�+iB���h�1���v��m�{^�ڒ�&�X&d�:�:�p�9��y���������線`�>�^��s�����uÊ�c���A�+�b�*�0h!�����n ���YQ�l�m`)P~/�J�}����)B\���X)��d�&>��p9��r5<۠�=�u��RH$`T;�Ad�ϐ��S�aA\ k"�F��	(e^O(&�s@��'h�V3
A��N�D�A�4
�_��|i�	��o�GN[�#�p�_P	�?؂3�� u��#X� G3�*=��2�LA����2������۷u�{)�@]�V  C~KI�L�����~�b�A~���>��F{�os4ӮĪ�*}�#�}Xǘ}�&�S��9�%���)�\x�w����'M�$�)��n&RO4���֯�(]'3���=�4գ�~���C�\]�ٶ���Y]Mc.I7"�D���w��.���[b�w:�1�����~t���Վg�.��>0���y��U�?6"�ʺ�q�r;<Y[C�h�H'"H����ꯜc9�@�@�1q��O�+�p{� MT[3��c$��N�����f��Xa�h�����^h������1ȁ5$lW�&QcֲI-����-�v�����O�~�3��e��b[��DX��k��[|mޢ^���?��?�a��A����o�I	^�5���6�X���A��as�Ni�J�U�I�Y��2]֐�_tx�fK���;�E/���W�]lqF��G��9�iyu?G0�*�71��Ml���2�І���y�� �Gfԛ�wn���z/RaG+C�h���	��ll�l\a�2�}��2��y&�ӯ�5i�f��w��k2��㸬J�`wM��\�j$Ju9�MA��^^,�a�'�Z@V��g����3�����n�=6�iJ�@oK�hT�q��(Ϸh��D�=@��cX�+�@[
J����q��D��W��I�xn�4�����ھ�O��P>Y��*�aJqwx��|�柰�?
��N()&Q�Z��� �W;��>��:?��?$��za�����z���|e�ZZ�ES�x�S����{X�h
�9+�2�ش�2��G��*���� O<��n�@#|�MG�VHI@�62��!��A�Z������_���q]�?���|�'�{�7߃XA���k���O��c9p%kz}�T1CS18C]x��U�mMa���4�-+�=����*�,S簯|����?e=��l�А����S���72��b~���z��YYn�Sԉ(���R�B�:ۓ`�
��x�ޥ'	ZR�ONpwP���YL�ͮoɦ����dFu�D��=��F�ن�P��TG���.w="��iڸ�l�����&rֻzN��)�P�B&��0�����ʳ����ή�e�� �>��JZ<����u-�!8���^�MyA�5U���
W���d���Up.�(^��S����!�,���� �oK؍G1��𵛹�m��ڜ����̐}�j($���&������	5(.[N��LTi�޲N��%Z�c��B5j��gJb��Kܙ�°Z��N����<�X*�7���Igܛ��;]X���a4j� �0��\N!��"��$e�Eռ�IU�uztN;ɰ��&�|�4יD�fq�-�ނ�<6�M�<�c�5H�o˝ѼO��ɡ�
�1o�D�Eޜ/f/O��8����Jƿ(�l�ˣ��i�a��h'j��2��Oӗ�kA�:��}w�� +r�t9��2���ˎs�F�pu�R�g�(��&X9Sۘ�r��:S�rtIz�����=	Q�{�8�ݠ�*4T[bU�������f�l T�P��yu
9�X�X��t���rid�؍x���
�HغR����}V�09GT�^Z�Y��`��Ąy=����r�5��A��Io6�\[RN���j��.7�=8��5nC
�p�C+g}U<���:#Ycn@�b᧤�����BU�Z�% 
ܧJ��tph���]b!��E�:H� ��~�h�(�'uPZ̭�H-h'��;L+����t8|i^=�q��k4��mzj��i����.��ϑp��Q_�����B.�������K<&�)�g���	�d�F���G�R�)3���):�>A�9tMcDӄ�T{?�ܦS,{�B����S�Z�aZ�3~+2ɹ���P����,O�.�ޱq!^�R�L�d��N�[��u�[��l�;j�h�,�yZ����D��ot`J�B�7@X���&O��ŋ����섛��U�#(3g=upi�Fj_@���ÁM­�A�<�V��g%Q��~6��R�]��f�7fP�)`���ۗ�z���*Ϳ�7��z��E��t�H"YC)�n	{��*�&�$:�։�e�+������ �E��Ž3��_#l,�I�#[���8��m%�^�qrG�>��jO.\��`��J1�׈��>c{s����HeJF�(��O�Y�ސ�[��y'n�`|[:0�R��S]tyc�K����O��!�����/Q�5l�k�RC�m����&;臕ך���+EN-2�xQ-}�J�H��(�|�\2��kV�W8XsKl�ߨ-�@�꘍�+|?4x�/ֻX����-{�����1�����WH����X�����>�o�٦#p�>؜����5��=|0�<h�c_�����&7�zd����������t��s%��2�DzѮ�����0/o�-�@��c�����s�4S^��a	�X��,��@t�g�
�(M��Cd�E�	���F��w���V��+r���u�ޮ�ݙ���H���eGPX��(7�}��En�7լR��-L�F���w���n��$�jMNAoZ�G��M8�W�Qqp��b�13`^Be�w��T=��>�I��*�S��Ǻ�|}�+5}|�_���ꖉ�Ι%	�N�8<���ֹ�����χ�ң[=��r����B�AW�-�� ^�>�q$�$o�n��9+��4M'/���<�3m�����RYG|��h���"�AzWW��Q��dӢ��Ӣ��f���L�f(qh���ђ阐��x���QHU!�j7����L^�)��K� ��?����s`CD<4�!$�
�}�Xm��g��/KMc`Y(�'�h�.��
����فf�>#ꊇᴼ��H/��G�ʋO[A��������uʊ�N�苽=W��De�j%�h���^�s���nO������T�g��se`�/�/�Ϳ�|o�h���ܶ��"����`�s�;��s�iz�T��V^����Y�>��鍑�Vm;�>�/,��Ӄ�Ů���}Kjs���r>(p6'K���ִe��+
7�e]��@%��N�@��Ɵqk�h��J��^m�١��h�9�^��d��K�,�(�f�X����sw?���C�ڽ&]jr"H�׹m���uD�F͐��ڍKV�\~B?B��+dT>6�+nw���KNDLH���+��{� ��G�| t0��y�]����A(BM�r��Rl�eQo]>,� �Ο���多��HMsE+����=��H��U^�����殔7r~�9/-i)|���vG�v:���{��+W�A~6�՘o���1�eK�t	vL(28�[�wػ��E�,w'�]�s$�h�s�}���>�N�����u�t�b1_;�~6� ٨�2��Ir���q�3l���(�i�NC�Bg��i&H�|������r�*� [ô�{�|���5g�T�.�\ty����w<��Y/ ��f��bJ��e�.z���-� �8 ���c��Xs��L�.���C�����U��ο�F!$��9�2c]��H��d)PIX�&n�l�����rɲ.�'��˾'?e*:&��W[rV���/'jYgs��Ŭ�Í�4?}tIY!n�*�)o�Zۜ�H��`�� rK��[��%�?�gZ;��N����?�yTߺg�ƈ���P�(�oU?PO20�`}ڰ�"�������4�ei=�W��Z� ��J�����A]�!���cw����Kv�Ƹ��q�h��)���]:�}Y����E�%��E�YHa&�2"80��4p��>D����l�f��Ţ�.��h�.�RT~��"����%1g��˳g��ف�jă.#0��?B򢃝��<��;TK�`�Cv�Q���r!�5 ��#Zw�1��or/�x-�z�f���L������䆾��#CE��%����Ay]��v��t�;V��?ڢ�nq��l�,�a�n�f�u�θ^_Z�1����@�+�)Im�GC�+rq@Y	"[ ���;���P���z	����w<%�B�,*���w1��Q��g,�a�I�!���c<�U�0��D�,�ՠPkM�p�㻶IIŹCX7�I���*�$B�#]o@��U^{�jo[�S1�`��*��sT6R~nLR ��K2���LM)�ޟ�N���NEb�����o��y>�9������������� ��8�U�������>vI0��1�>X�G\����� �i�����Z �HUt=��*��/8*`�q���q��v_��J�5�R��l���b}fp�yy����L������O���/�UTj+^�L
��5�`�q���{E����y��(�U(��E���
����ٯ*�k�7 I/�k���s��:XU�(B4=J�JZ���*�W[�_xQ��C��q�-X0���X�]vp=+������cA�F����?����ܪ"d�Nշ��BEm�Z3��'�$(?���zn��~&�]��My����TF��7�4=3h�2Eu�ժ�º�{������ܯ�Sj`�\T������w>�ơ�������W����u�f����3��(��*骘�D-e�i��=ee��iu��B�\��f���-oɔ.�(��n9
�=ܳ��0�*�ǿ��2Y�$�����w��C�j�l1���<�Z�Ի�B���(H���E=�]����'I�H����6^�K�TaE��a$��
l�mM����'�	O������g�]���lU�`0K��;���$����n8l�Me�Q��)�t r�O�+���5�^�h��?6��M�ObF�����9�:�O"��qq|?ǘ��Q��\m(KZbHÔ�).H��y> ��WΦ����!��)O�0�jZ�3��?2\ރ_7�&��O����f�Re\V����i!J]*y����^��?;tr����O��p�Rx���H�v���zڨ-B�B�'�Ď�=���OJW9H}����,��b���=e]+Σ+�H@Oi��H�O�4�4Q�cTtO����OT�����=|��Ei���Oi�A����hJB�h�Ч�<jo�[��*'o��\�� ���@����븆V� ���ɼW��_��I�,S��w�e~��XKΜ�o/m�Xh�jf`ׅ잣R���S:��=����;JE�sʗ*���	;�G���!��t�w�I�Ӌ~�º(~ҕy��h�O�!�Ȅ�6�q��o�ݗ���Ũ�]*�����@j�s�z��TK:�J��^E�3�w�1<�}~�S��~�����D�j���R�UIp5�I~�kB�>댘澲���K��g�U��(c��u����횊�O�7�B
����_'����`!���F�<�~�U�ߣ#{�Z���b����siZ5��"�OߺFOق�������!�qx��jk$~
G�*���!��yV�7eR�Γe�#��[�)�����i�i"��Ǆ��\vEI�>�}�g�Ք!����⠌Qs��U�����|��%h�u�5�����(�P�rGꦵKf�,eS"zE�Fa�?-Q����C�ef*���EcI5?��Sc�(O8���p���E_�Y"�Xc�Hv�]���A�9��.�v�<�����=��N��ر1��Ǹc���c��S��1�Amsh�G�O $+17��X�܃�柍ȹ�5�-�)8���L{�_jgUڹ�׭��Ra������&^���_�k�.������e�b�}c9 �1���Ĝ�T������p�d:��*��{�e\�����`�� 
�*�(f:�}[2� }`k>��$�"U�*LA��_����Sl�e�����;W)l2o<_�|��3��g��C%뻍��2- YCV����x��Ųn>Y�0u8xc>tL�9�Sئ[鳠���8��%U�`_!R|g���`���ƗW/�e�\��պE9���" 呵��	�Ｔ'Y�����_Y�p�.&�o��G#��8j�)�5�.�2��t���m��m8+��p�T/,���2N��m4uh�P��,�q歶�R��U�!��D��r��M�YDg���z&�rK%���b��?�v�g�6��⭤lG��m]��8�_���-P��:�2��ւ�Y!g_��W�!0��oMt1#!�6�Ҳ��\;�g6v�r
��:�n{��4^���g����ACߚI�����/��/���A8��:"+�.}j���!Z���x3�9�S��U7cIك(����љ�u��D�V���_up&�_jz�)t�+����s���)U���.e������J,��Ն�j�ǣ���{���O|�M�#�f���W���1���[VhP�0/�dbu�4��-�r�N��V�믥�=���L�@-g^������@��<����9��D�t�3�
K ��YZX�8��w�"`���$���<UR�.Y� ��o��������,�&=&]�8��,?��tU�"c@��⾙��0_ZI�Q�/O���	�fceM�a�[U״���J\�x���{������q�T�ɼ�A֢���f'�/�Z��)7���@˕4��g]r�7�	�c�^�`�31
������~����Ζ�e'�������7eF&�v�;�h�
6X�+�<�;�ۇ����^/rR\>ߓu����j*��(F�4ۢJ��H/N@y>��gP�K�8M�YmW��oTn���
������~��d�i)f-Z[7@�ׯR�s7B���Vb�t�N����=m�t��T��~��E��1L��}Gٜz?���^�����>�������n�D����|z�I���(q/C(�nCC��Wb�2�;���פ���^�}viY�^�3��dq���3E�WiqG�TMr&1F��i'kt-�W��$W~�B��#���gUk�Cy��"+ً�T��Sq�)c���:A���W�{�����"�����wB�[�UmQ�d��t<�Xr��&�!,t�J�jQZ���$��	���hƪ��`�HI\����ۧ9�^���]��,��F�ZlLC㇠ɼ���� �҉t�nE��h��O�0A�C~��rі�L�����.�c��m����L��=��̶�<)(�_������y���� `��l�m�p���:�<۲���s�0�l7��s��ɥ�j�T��K�����:
�R�����v����"�?Y�Tl(�;�}P$�~4�	(V{h������ �Z<�_f���f�!�E(�u��x�eKY:�txn�M��dj�H�*��f'�J�1�
@"j�D��@�>�k=-����%��Fΰ��� <��=:�{kx7��aB-$��Y+!Ǫحd�b���nԬX{d�Y���N2�2W�y��a�0��ٗ���-�j����*��j�չƩ��W�ޒ��5aX�	r!l�x�5�Aߖ�\��6�C��ؼ���)�\��B~��L &��q�V�/���~	Χ�	�o��F9̅Ps���5J�I ȕ<g��������x�ժؿK�L��'ڵ ����x���ܒ[C���"�y\��Ѻ�m\��Q|ٰc�0�/5��
�m.��j8[8"2��l�~x.�)	\{�����%ay�����G;�\յ�w�}/Z3��\qx��w��h7�i+��?S��R_~��1�'=�;,K�	�X�yH�ͺj���/v��P?|���Vbf�b�
����S|�7��nҽ��}���� �"A�����'QR��z��n6 0TC���訜Uϔ>1X���0N��Ίk�iU��Km {�)o���rjA
��U#Oy
��@���٭6/.�̓��0*��yf�7Fw�:3�G��������o��d�j�� �ܱ�]���P	��,[t�@0꘱�DB�dOǜj�8�Xr/Ol� ��k�&Q����P��җ��>o�����]��&��Z@'�i�;�+��Q�:�ǥJ�����7o:�^�ٛ�)p4Ɵ�d�����v�;z��0����꾇��b���D-E��U������|?hVV	��a����o���0/������H�5���~n�wu���8B���P[MX�oz,�RR�-2����lg�|�&$g��/n$�h��d:��ޫE��S�q�|��1n�j��Fn;զ��a�Y��6�l3�| z� G<��%�в��R�>��"t9��TD�%q���|�q�ߟ����a7�{u/ZW�<���&Q�	N�9��;a�ppqA�>S�k���<�+�=S�
�JkGp&rR�����'
�;S��w�{�(���k?��/�+�t^�B{.�9g�7��gi[����\�l�l��bA�r@=g?K>_��5�`XX�/*m�9l����I1Y���06j�c��(�A#�r�o�.)W�$Qe~SB?�D�Uȥ��cJg#�Cl��Z�r ;*���|�!��D�t�u�a��m�H�����.�P���Ɖ������qRi�s̳��U�F�{ �3��;L�Qf��P��{�(~-�`�Z8y;&���{].	�/|�� y��<��j�C�
UO!��7��I?C-�c�g��(��g�>�RԁQ����[F��.4(+��3��oo�+�������=`T3��P���A����M�/)�Q���d��}Ӧb
�.��y�Wg��Cd���.|
�Er�M!�rݻ�Y.Q�I_��;e&��}maD	P�(L�ĝ�V��|�~�	��2��,'�K�ܺ�e��3Ǧ���Vb&�%t�Ba)P�%8��Ԓ�0���W-v���͹��Dj��(�����ۙpu�{8�h�Ɔ��0�	��l��_��,٢{�;T96��������|wjl<A#��u$5��Ü7C��b*|n�bA�*�@�T!l,�_�]{�ي���S_�0��bT�h;�M�q�K��h��\�?W�����n�������
7���u������3�3�9�O��U��"f+u����j�V~������y�u"}|��5��Aʸ�F#O�PE􎅥s,���q�+G�����y�}����E����5_fQ �Θ<���B�ص;��P��!����r	�8�^��A��:�*���H��(��i�d4�<[��\n�g��;��.6�Չm'�����2É05��D_�%!��#5V��g�R�x(P���� U���B>Qk&��h7^�bK��R��i�<���}0#j� ���iĬHE}���ansB�gl�aT��l��T2oS�!wY���mB8����Z���g v���0t,���zo���,ڣ���Ǌw5g���"s]�r�NG,C�YgKѩZ72�*��~*z�oԁ��=J��D��� �KV���� P�K$���e�J4�@Kh#�C8F�����}�[��`PC>��`g��S˛o�S�)��ծ��B��|
 ?�#J��Y-&һzz��oV��2�k���Q�>L��k}�<�4��J N�E2�}�/�~s�P��+��7Z�As������8�*��׷=�����MNE�G�I2�!	��OgcJ��S�-Oݢ��%�5C?[�K�-���/ ��޼� hf���h�����������b:U�/�a%�g���G���o5p�K�9g�'�re[8�ko|Ꙛ�	�@3�0n�`R���+�'�}�t^5�U��^Xx��lܕ��`d�d���=��+ǵ�魎Y}cۃ�M��ý�,`?
!�C�΂a"y&��dj�IO�(\z|���2�$�V���2��,%*=�hx� ��&&ꛘ��ő����gۡ&��ʊ�h�������ݷ���� �^�U#%'����܃�@���cl��8��^�b}U�R};䙸�͢|r��)�;�;�ĕ���6B�	̥�	�DA�!x��
�z��Ьh��׼����l��i�o�Ls� Gқ�L̯.�,x%�ca ��Hga~����ԑ�>akz�ח	?��_1n3r\
��}F����z���sEjSN��E:B�� wP�MGu�Ҏ����zJ;_A����,��5��6�! W��{�)�
+����A�����k�6����d�7��.��w�@9�wW�B��4yS&L�;�y��(Yt%Snt,X�9?	-9N��Ke�eȅ/�E�}�X�.��	9q�H8 G�l7�;��e�E�n,�\P�j��#�i��P�3p�y��g1I�J�����Vb��u	�,C|E���� ��E}��?߈i�kE&��t���P�Kβ����G/^B^��'o��n;�B����xk��c-t
�ft�>*K����ʘ5!k�"rJ-��#�`J[0����̧v���[�TWj�4����#��;O�]Ѡ��u#l��J�>k��U�K<o d�k�7b�lx[�#g#B*>B����K������XL7������
68�E����2��4���`��2�_+}�����J�l1FfA����&L X  �\.d���Yp��H~!�����٩e�ƏS�9o�z�[!� ¢�3!$X�<Bv�F���W ����Q7�L����o��|ㅷ� E�i{o��i���ڧM�6i�=}7�|��ݳ3��Gn��)T��BB�{`T�*�;y�����T\�	����Ϭ������@��N��r���S����<��[VV'���)��
'!W�U��$ݣ;����ŗ�@A��l\�O��g�L����y�l���5�a��>9W�QG�'3 6b�;Ҕ���|�0xC�k5.�8���\��F���5M�80OM��d6O� Kܙqz��LGD/������m��ԏ�W��h�	,��N7t6m��d���Uǵ�A�Q&�;��\sN=��"�vW��'�U/^f@@�w`���lT����݃�xܙ��*��>� f8qw0����Bh�R��I�q�?-H,���w�ހf��"6�x�������L$�)ac.�7GA���S��� �L
[ ��S��IJ/�=��?�R�K!q��n���s�;�\���dM+��˭V�sՂ>���pHW_2����ֳ�3�d�S����������	b�8�/=����Q�xP�{wQS��W�u�h **@%��&U�²1 �w$4�E@�?=�����4U�Ch54�ߔ��!FZ[*մUx�M��"h��<wI��'1#w��t��� �K�
�]��(\Bn
�����ܴ֞sջ8/&R��rn5�v�X��FILD�B��4��`��\�rZ�Z�A
"�h;��G7���#92px��\��q�>y��CJ�j{�1>� �h��<py1�)�tF��Դ&[,ȋ{�^�"�o��_�V����9� kw���q�6�w�$��*�-���N�&zY輻΄Y��)�5f�'��X�+��Dw�~��^��r�b?��Φrۈ!7�9D����Vo�C�-�����^`<����-B ��
�<���P�����ۂh�ƺ;<��a�Zh䪭V�@�c=2A��[<E��}�`'�9�'�S�����0�v�מ�q5�G�,8�◝��S�I�/�Գ^���"�k���Uϟ�>�~%MO	�Qy�z?��@�0t��w>8�� ���X���*������2��iP��M� E�τ|d/-6O�ݫFT���1V�d0��U� �1)�b��v�kT�(�4u�T��Rm,:�=�v�<���X�;(t��g~�d�#2���-�q?ЭiͧPg�٤�<<�6��g�3>r<^Wl2��9���{��$L������]�rZ3�C⛾�o��¬}^�G���;,��`����c`�J�w��~ L]�++/>��V�����%��jp�V`��_��}���J;s� mkŘ�Y��#Y���<�cU=��KRO�b�ZQ�)��i�g�#m�~��@�J��SP)�#$���&�Q�?�D��)'�B30 +����u���l����Uu ��-v�C��Ck�_��->ۑ�=��:'S!tPX��D�r!���$� ��ƅ?������%��P$r=�	�]���V����1ʔx�$�rя��T��p
��a���4��]�S�#qiV�L�A�<�O�H75�KY��w-�ɷ*���W�n14ُ�C�fRH�X�ژ��3��wӼݨX�������5����Ѝ��>�A
�V\�]��ɭ;�k���n��z��b��%	i��)`���J]S<R嫁����>c� ;�j��n��&O`xUi㔕�gcg_]� ���E�ݽ_�_������H���3=����fI�V�^�OP^Ҋ6�"����Lw�sq-�H�w���b�/>��[� ��M�CL�4���V���$��B�/g��#�PYܔ�'�t�4Ǭ����ƨyd!���)�1B��x-���{�~^��)�ݒ_*'�i��Xf�?j)пl]�tܕE{[^�H�� 0��-��	�j���U
�X]f.Hl$���)1,��c�w]-�.ܟl�������ײ�������e ��}l���=����d��:�<?_�t���=ӷ�%��3��3q�#�ң�.�E� d�ˍA���A���z�z��j��m�7��k�!�6L�^�%���Y�t���m+��96�H@�a;)��tЪ?#���V��0�=�|+�$y�J!�.�7��#G��������[�&B>��w��HVu#������
ݮ��V�w�: �8���K $���;O��s�� ��ߺ��E����-�2>^<2�A�%"�#+$,s��Z�XM)�T:��`���vNg+ĘN��<R0�!��T>u(��d���@�Ἵ�5�wn�sH)\e@{���If����_��.h�ZШ��)�e]����)��id�`��I)M�����;�1�����t�p���Laʟ;m�����aG���d�c��n7�+ۡ1�9W�7Ċ3���A'��$ɖ�m7�ǼS.�Kh�SɦtmU�r�$Yk�ﮘt�A|F�Ow
�d�)�~LdH6�L���0��(�߯:�k$� &�Η٘�c�E6�����֘% �iP�7�&�i��c��9r��� k���^`f?20��چ��\��}�S&n~!f�?�(�����b�tA¯%�*��+�y���	
QE��:E��>�E��鎷��T�ZwM�l-Wv��Åa�|�v7�C
�^�$�&��9X�9ӄ+�Ε
�W,�)6��%�|%<��m��¥�����&�7Fc�u {�qG��E,yB�e��pI&������[��d�5	D��f�r���;���P�r�'Zτ�@�ڏN���7�`HB�d-k�&�6���{7l����^� 4�4@�m�$V�fΰD���f�_:$	����㩾f����������`\D����Y����\aQ�d�t%g�	"y�)Of�K���/l\8&`Ϩ�<{N�2_��Gy��;M2|a��ؤtR�O���h�q�zk�I�$K�3�����5�R֑���`��X��Y/`&@�����jD����N>Y��Z�m�V��W��������b��f]� ș�)�W%n��@
&����G���Y�����h�w�������d[��=�c�tL� )d_��D��]�4��yh��`1iûm�"g��I�����N&j��o~z̋J��>H� ��A���g'XĤ����i���J.C�RKl��~K�' 0�إ�\���6ɴ`j�a�&�����c�E�.7��=絛6%�L���A �|>D'�ٿϔ�v�V�G"B��Ui~�%�7��w:��E������ O��UO������2����������j�1/|��\�)��+Ҁe��S�Ӈ���A�ޅ�����m��m�M�'���8�>c#m��B_z�-ngj~b���&(�z1���毉�1�R }p�e�7�//�v��ůͫ�� ��˽0ƺ���(lP
co�-�ղ�R��K��V�%�	�0� ��Kh��à�q@U�ᦾ���)s7�����X�Z�v��6`�D�& �ܖ2�.�K��d{+\�@�+�}>NY���kId4�ʋ;��D��1�L5z_�)ײ h�%�R�'�`�B^�Q�MP�,�	oo��@�p�;����,ME��%ץj�<����=u	�U�����&�w���c�跽9��r0���!��44<���A�qNنS��tjY�J�
�G"Ń_B�b��.7�){k NDr�G�������J�4e��d�.*�o��^4�\�<������"���R�8�L��=���Y��W��`�P�z`k>�0�*Ҷ������!��r�d^T�����G�sNل���S��}�����4e���oE48d�� �3�K�.x�w]X*R!|�d�6���7�����Þ  ��p�S&�3�6l�ɛ6_�Wլ���'kv�L5�.��_��/ф�S�_�DJ���)� �% �˞*�"�����΁�qJE p~C�8㭛&�)���!1�ȯX[�2A5�2��K�����T�����LZ�Ku#Ί�&��F�4�߬�z��'�pf:!�}�Bh-)�����I��SR�Y|�
��#3��m'TC/u.]����S�3�V��@�pύK��ސ�D�(-L����J�&�����׽�H�WM�� �ο?f���)HF�w��`CB,Rb��-��K�0il9��S���=g�%�	#=�ۂ�|
��Oq��)���1�͙�5�f!-�ǣMs��Q2�S`��볗W�mG��nON~�JMz��$�NU�dh$�ܒ
GVBWX.g��A�rW�=���(�`� ���^P��e*��\H���CJ�=�;�"�n��!;�Ƀ�i�ߑjv�s|9�R[��1�y� ����4=M@�<|jaK,������L�%���@��gQE��27�-疃+y�φmi� ��]%�l�t�&Hk�*r�׸�^��c <���5��u�P\b�44���z#���06re�@t��ՖI�r���g�;8N�0:e�\�>�7�c��<�d?V�MK@������r<��5�
<�����tm��c��һ�%9x"I��]�
7ĝF�p~���eS��Hc��	�����,n^>,���hҩ���V! ���)n��
�Aa��'�*4�A'�"��p,�82;��1�x��vev��]���R����V�>Qf�ς��=����O¤б]�|�����ˋ:�Z��.!�2�V�T�? oEE��p_��]5V�����*�I{dl�*�խ:Ǥh�	{ě{�r�1��a��Mw�`�g��2��/���#�|�Q�ہ;�� /ru>T��wE�ˡ}����1�XX�c���<�G�{e��lN`���u���%�-��o J�p}9Lo���V�5`�z���u�5����������-]�\���y����R�8U�iܱj*���
,�%�o#Ƭ?Lu ?�72�/ɨ�o�j�o�Ԥ�^���{}=ȗP,v�{.9ͬ΄�k�4�N��t��������5=�TdEK*��l�b-q�	C�`�|,�\fr� ���B��pC�b��)���94&��]_�˫r���GV @���Q�vj�?S��8Z����X���e���ж��S;|�vm�4���$��G9a|ź V�U��O�G�څ�����Ҳ2���a=�ѣ�qu�X����Q�A ջ+eKۮU!�̓����ظR�O	�en�����^|�7�K+=R���`���9u X���X@#w�d.��;����m^��T��ӳi�cH��+�%2��r��ZX�o"H�Ci	��	��I��uE`�P�_�G�����M��6�+�dU�����M�;�m"R������R=�4ka�ɂ
C�1�0m�j�s~L�5O�UƄ��+����,
3O�����t�9�݆�;���o�m̤��(�8����tc�N^I����g�^؂,7����;�f'=�����ӁE�x?ͬ�('����OZ!�BY5��P�=6&?M��`(����"ƻYI�l�:�>�E�MY�3uM5��t���`=m�]F�n f��@炙�<-x#�J �d�,d���f�/��ѯ�M���E�;.$�9�P;��+�(��`����v���p���P�b��	��+m���o��xj֎~�����a���O�h��
��QS���#w���dR�At-��^'�
~'���Sa~�@[�3��_��Dߩ)���G�ˆ��18"Jx���g����^��䍴p�~�S�rR��d��
8������+DC�I5�[���	��Ąbyv��a�Í�w#*}�`W�kŭz����.��A��]�jJ�*��^w��5d����{*�=���`�8���������E�jℐ�@� ��W��\�'�&�Q���{����'�����zx���j��.��n�;Z{ֹ��+�Y���+#�A�5H�Uo?��'��8M*m^F.|�Bx��Km�/Za�jrAS����c1���|���Hj���۔h�z墭2E�NQġg�7����z �T����4IX\��U�4���?�x��'��w�|����oڼ��S�ȁ
���x6��@{��l>�V*U��)�(J�?�4�M�ř��Tb-!���˞-y�y�o�C�6)�d�s�9K��q��Ux8r��qy�t���� =�$U��d�f�4����[�ԾZ�^�m�k��Y�X��@-=e���Z��"+�>**=+��'4aX*������#�H����>�#�����|�d�w�E�pB�D�K���~8��9Z���M�	�$0�Oy�X�h�����lg-�t�Y�|E�F�z'���'��vG�GHjq����bϓ^1��he�]j��X�ڒ|�A���N6$c=hS.!��S��}��������K�x�sR�߷��#�F�gF�|���¤����s�ݔz�Z :�	j��'@+���}S�0q����=ɹU��'�O�L�u��V�|��ZcC���{ϴ��3 �|�4p֙�{�SҲY� ��aR���M�vI[��6C���jڸ���g؅>F����c��n����EG��ηZ�BqW'ً����O��]�>�����~�/^�W�ߚLp����>��p� �����(DN�-��ܨn���c��V}��,�����)��4>.��l��\߲�5��g8E?�m��p�҄��r�(m�B�瞌j�^�: �����Hr(��Rm�����Ii�����l�`[RwHس��Xr�������E��U�� �x֓N�c���L�a��~D����-녃�lv
s+�f�_�*���O|q��!���1�,����1������|���xM�z!Jb���e���s2g�[����!���Jrs��N�_�y� ?=X��t=�LL��(;���E���B�|<��Z�C4�B�_R�v ž���m�N-��Bj�H+iZtJ���,��y��br%�,SPe�w-�"7��(��柁�@��T�[��rKhL]�8
?���#a���/�e{����r`VP���Ի#����Z�U�.��i;�j'N@4�[��X����Y���wt�X��Q��L[��em��P�BD�ܰL��u@o�l��[�V;� ׽��۱�iM,*䯑"]&>o��@����ܪ��b��an#r���X!;g ����3|u���TWv���_X<����J��9Z��G�,�!��Zth���dt.-8
(Cb�I��ri�ŽFs�b�,�Ɯ����0�)��w���\$	��RJ�7��f�׎-`z���R�W�>���7~�HY�Ӑ*�9���¸�!2@��=r%d���^��ڵ]B!#`��f��H���
�1;~�(��˯�_ɣS���Z�W�w�0XU�d���$��:&�nd�?�5��sQ��Bծ@��e�9yʕ	�^a4��E���F��ӂš��<�;��t"1H��8��D��S�����R�I�K�,:�9����9�����V�������t5�v��t ��N���CH�b���պ��,�� C]M;E��
�ƥ}X�L;4�u���2�IVŠ��\~��ïҦ��yx��Zt�ƚ?�؀�����;��ã��N��oph�V�G(}פ�o�c|��Έ�$�I�S�==rs�"94�[�3���!)4��^.��l)9V٣��C47�cӸ�kf��R�F�/��;p~�9�OD�t\4k&���0F�����7�}jn��|��H�M[(�솴U� z�3Ve���C[��r^A`��ٻ��Qr���N$�X�-L7\�)I,��7E'�/��ME�@��L%J�P�,
�=gC�ༀ�Q�Z����q��SqI����^1������]���bgk�Ħ���R%�<*���l�yõ��m����,�D��+CR��y9G#�[�}�`���"7i����_9b���:uZt�KC _��l�ZNҵ����и�?|��a� %������g���w*�z58��̉z�/9�j}�mi g͟���RE��~v�p15����c�����a[jfO�6��o�/,i���Z�.7�L|8,|-�Z�V�W�.������B�2i��eE�L�����
L��K�;�����p�ӹ��}@�?��o�l|fs�_SE4~]��d�񀽛>e5���|�Ga�là��Eu�΃�]��_�~� ��/��� WItq���VJ]�p�n�ܺ���&E! b�����
m߉�s��y���n�d��.jJ�6b���\��i��c�C���_>Ac��Z�D��(��H� �!0��i�%��=�j����jF�����+�SW�o���ā�;���8J�D��xe��
ʹ#���w`g�`��=���f�x�jQ~V�r�0��}���)p�;,�>�ݓm�eT���Ǔ&��5�1���m���bg6n [ߤ���.U��^Ds|���ύi�T����D	X�**�<[.&�E���m(������>8������:Jm���Bֶ�!S��ʰ�_�G���������K�S��\��%g|3@R�f��
�4m+�s���`N��i�#t��Gfԙ0�����~���|G3P�Ţ]=��U���� �Q�v0��~���>g�P:Ԭ߲F9&�o����
�c:uVTYw���9*�:_�R_���.�8�ݮ^^U�+l��T%$��y�3�\q��R�J�9���aӑ�pø�)���)���s/�
)���2}tȓ?��ye-ݎ9Q}�������-�: 7f�͗�� nO��Y��"�%�6%"�ܷF5���5#E)��r�y#���9P���'}If��H��9*������師l��L�Z�����_�
$�b	t�Ar+��!�U[��Z #��*k��ꯝ�W�>]�p�z�
�C��ԯ�E�5���l���=r>�i����o���͗y����7��6�r��nH�jc+��{��&��K�iR����Ik�5��>����^�\���4�<�=R���؜��x^��TgK�B�v37e�K��9�ԭ��m%HpU�j�'l����A����N)8)8Y��@���������-x���cL.(��{�U9
S�ܗ�\�~�ۍ\�Ʀ ������7��w�h�g�װTY���R�A���VKh����xȞ���i� �HNރ ��mJ�W"`ﲒ��=�bUleo��ɖ�l=���j��T�u����ǲs1*�Y��~��^�Ļ�6jJjί�/Ά,0C6���h��Wɐ)K2M��[�x���G� �[���M0&���s櫡b�9J��b�+�:hN��(��<�"sq�����`�_�@���$ï�������9�4I��E>�4H� gkf���X��+q�/D˾���3LÞ��h,�\l4������}�[ރ��"_��+>!?���}
h��"Uo�"� ����)�G�Ukpԛ¼��Ԉ����}��D�;g��rH�v�t/oB�Lh�*�ԉD�57bW&����������}����Gߐv�n�ۏ豼^ҋ�n�ҿ��x�,�(��Ji;������d��<�K������ֺ���de�%OT�}�Vԭ�m1qҞ�,}�#y��/@�+g��nҕ�U��T���ˍ�&a��˿�c���
�\'��:�zl�Kr���H��yz.�r=��~�䁞z�r���%�ΐć7�� ��蚪ީ}r��ᘆ�NAu��cT������u�E�H�r-�2ӕ��p-��gnG���oh@7T���f��2�J^Zd�&��[h��)�\v(�Qk)~��"͡����eqY����Hչ
X[�>^mBűL�M�H��R��5#J�U9��D�
_�>��Sq�EdPUI`�KB�̼C\(���|� �G)Sb��-Jr1Xx5)Ҝ����O����q��w���+A������IOv�X_I�Bg��e1~��ܙn�9�����@��������9�p�7����� ��0�1\��a�n��*a�KT���֭!�4WD��5$2��?X�b��Z������ݟ�������<����H2�hS�� �dfT�j��Ȏ]:�0��-�s|��N���W�+�j��4��1� �_fA|�* P'��
H
H8��OCᮝ~{�� �E=AW�W�]y�À�S7���܁�7>��I��j�x7��X��-Q��ՄQ���ļhhJ�b�o<e�
�	/T,?����^����$M�j�w�.��e@��M,'���,����y�?�������2�E�+P�VY�����R#� ,*b������>�MnœZ���[�6f�_�K<�vk��ONl/ve$�eC�=ֿ>�g����ړ7�#)���L��m��3C��p�˞�[���T҄!��qh�����>۹"G��A�K7D��`�z��T��������u�m̶����A	�s�}��MZ�4r�A�"z6��} ���?ᴇh���:�%[i34�
Mň,I����߬@�l0:��癱��B���%I��:�V�YE�q�7����?0�v�wЬ�$[W�}�ܰ�P�Ě�4!�����K���n���`�!#�AK�\�~I3<���n��.�BvW>��C"z��vM� f�}�����.�Mi�#��|4�����A���Jױ���8���.�w��$���}n���}k��   ��4��w���RX��||h�K���,B&J
o�x���������}�ۨ'�;�O�Q˺�"`�f��O^~����W�ŎV4M�0���N�B�2�!��iYHܰ��q�	}�km�Ob�K�q�#S
�m�>*��g�����U]m[&U��)փ����O�����-����5m���{��?�J0j����Ok�aɶr�-�q-�0���ʂ���f�A�z��&P5���멌��IVd�6���޻:cμr���Л�
�� �u\��c#p_^��8��j���Qm�����c�Q sLc�!��-���m@�s�4�`tW�Uv���c�x����9��'&X����X�C�� �����,,�?�I�mq�����S�sh�q�q�oiDn�X���6wՒt����ЇS6��{厊��(��<�����8��!&��EX?9[�dwY���DQ{�>�k7��{c:�`A�*ǒq�2�e}��kq2��p����]�I��B_�-�L�/���yS��-�y�����HQ9yq4�q0S�/<E��L��j�d<�'G��k�fK�v���<!7��y�~�
$�b���T��QuLҷ���f+�~����T��L���37$nGy#%-���6�V�)J�/(�A���kgI5=�K�P	��5�A0��&�|ЉG�]=��}��4�ހ������*W���Z�ZV��z�<säJM$q~���xd��#���PZMc[����L�U�Mv�S��1Z��-���8�2El�B +�fɂ�1y�K`U���㣎! ��b�Xf��<�����2GPEv2�E�YT]�O)�vpc�#����4�!
��8	2�%�t������o�~����pX����\�lY�H�b�?i���os��B�%Կ��r�5o3\6U:Q�]�� �F��k׆�q������(����7M��ܶ�22�K���0$aM(� s��Zܩ�U��}lNB[��J5U&����br���B�ʛ��hF��,�������!���V����kq �}!(/U9{z/R�+��"���t"OY=��c����quѦr������(�a��ش6����ؔ�h�ƒg�yD�T⯫fl�����kn (��c�����pŁEP�}���G������#|�j�E��R�j�L�_�'���vP[ZY�%����׹ĵ����R����C��7�� 6T\*W}��-5E<��@̐�bZ&����fu�C����j���	���؍��{]�
w��m4Q�1���6�t�SKHz���J�!u���M����)�q=<�xv��֩�8�	�<�dh�gw�"�Ԉ@A�����V���Цw�������̧�<N|}̅����&�q�o	դ"��gʽI�T�A�`{T���+Z��-<3�{��>vP������'�U��Y�����;��총��Z`#�㫕!�3/����<H��(��@�&!�$��5,]�l�	��Qe%��Co�i�5������šG�]���Ici䗓0vp֯2jgh��0�%��Da\��账,�h��:@���bj4r$AؔY��>���Eä�IA�M�+z�H�I��dJ�{5tn��2"UP2֤+7�>|E~�\��өh&/t�Bn}&m�N�C����HeX����\Sc�Y�M�l�#�N7� \��E&%��B��I!��.�%�)`�ۃx��6o��42�>(��Ȣ�L�V��O�µ����̛�$�#����%s���f:�8 �~2���!���/���R"��>'m��)����O��R�#��*H(~����.F�����o�he���$ֶ�m��C�9�	�ޛ���G%�����S-�����s�W[,�֌,^}��"*�`��}�W��V{��s���9�{������ؑW��;t��Ξvt� ��Bn�ృD�i�6+�U��T��v.��FNu�]�\�A_�w19m�q���f�<���6����k�WY9ID8o��3<�G`����]Q֙&)�������@�D�y�h�;ׁ�:4eʦ�"��#b�a��&~�vc;IPv+lV�ak󕟑G��*ܖG7K�����9�9�J�n���L��x�_S�Z)U���cU�=���b���"�h��V���1�̣Ǘ��Rp/"M�k�ť���)~3��(�	Q�{�b�ov��q�!~��������	r�%�&yH�� _:�A��&���vH>&��	EC���f�h�[%���z ���_5�i��%�<6�O��G�31�"%�w�CC�"$`~�<�lNj�>>\�h���P�qRH��
�})�MXh��Zң�3U���4Q�%�|���3P��[OemXN���c*�M��z8��V���tP���r��S=�FIM�̅�C�~B��?�qN��T�U7���pk���V����>��:SNYȗ�T(x��8�^P6����RhN�o&���3.+�X+<�G\G=|�	e�*�l�:����꯺@�Ѡ_���I�N~8��֒U���.=�$e��ܟ��@p��Z��[ՕD� ��;�����/h�J��'KB .}�����R���(��P�����v�%�#�a"��bpD��-J���Ϟ?b�tCB2����c
r��^��<}Y�C��;q��>�0�m��^s��mL�]�(��������;Б;���5]?g~�E��������2Qn�6\�����������<V	(����X,2Me�E/'&��.�I�D׿^][Ը�/�@��+��ڀ��ϖ$�㛖�s����m�����DJ'G�w7�ݨV
N}T�y���`���QeG�H����2;�_�G��M�t���y%����{��Lv2���U`��8!o��"V� m1T'��@Z�g
�J�)o�{)|��v;����V�3[e�NBC��p�����V��/<���hZa%�
�m�(�!�"�[��"�Ԅ��M�C���1���>�syb~��"Ԯ=���S�'�� )��o��Թ�tT�t�2�	q ��Zx�$��[ˮpC���S���Vo]�~�!h��Z�`W@�q�(R�Yt&��M��(�����QGK�كQ� 3��r��p����1ˬ���I��i���U���2� ܆�:=����˛|��[j��&3@��x��T�̲���*�*�8���A/�R��փQs�h�����g�k�E�ڪء�dc�֖�a�H_���6魞Ħ�W�<p���t�-��l����6����(
��N� ��aDD3Kuw>h?]xF���xg��1��M<'����oJjG�oP,2�Ԣ\!�
@�a�&�W��?r����H�<H԰�0��� ��5C�GS�r�9@�j{P⳻���		9�u�maǓ~��X�;-�N��JdL�x$�}V��aW�8�1��f��p�f:E��Ǘ�	-��T�$H\<~Lľܘ|�hأ!?ƞ�T�>��@E;��$��*ϊ 7��p=Y�N�M�Cu�]�ρU��2Ԟ]s�N��n	ɞ�bWD-E���uT�Vc^t�n��՗��+�x�dSG nQ���!�W�,��������������+=x[v*����:���ĕ;����k^�����+3�A���A��V8��W�T6Rc"?�1�
e'���B�l�������1�����K������fyyL��� �1���A~�و3���2S�D��e+3<%���$Z߅z	Ŭ.[�j������鳍i�`�2��
:��फ़����Nb7�mV~@�R��lܪvyi�5�ó|.o�͟w�gFgI��!��*S�����M���h�CP�,c�9_�4��F}�İ���F�,q6٫3���O#�ߟ�ux���.n� ew�<�Rp*.}��N��1�Ѕe�q���"b0&
�"Y��Q��4K��b���ks�[�MZ;���7�A���;1�u�������z&�����3���G�U�U�
�;O9{s�"v�P�&/S�]�P�9s3⥀5_�5Hm;v�$�\9��PϏv���WoY��r8�螄l�z�u GS8�Tp��cH���[���ݐξ]a��G4����I�Z�#���	U�S��"���.����6�N����sk��r�r���NK��i������K����"I����}���[�l`�H��H��18}tX�R1X��@�k�O�
�(q���;M7�ekVt03C#O�V��j����4��n��O:.�w�`C�a��l0O�����D�|�r�~]���T�U�_��7���u�.��q��F�џ!lR|'F;��Y�ga��r��!����!p�2�PC$��.�LU�]yW��E�;f�ܬ�yN��0�/.\��s*�>���Q0G�OJ��W�x�m �X1�A�8l2����՞��ޟAC�b7�BF�M�$�o����xV�J1T������֫"����~����C+�S8h��FWM1��	��~�L��H���C������-�j��1MĂ<��ot]�9�S�w�����'w[�r:s�,���zŹ����
o1�t�����O�y'^p�"�LU'�Fج�����`C~3���"��0G��q��ڼV�1J�+�ױsL�H�쳶�(,���ү��s1��a���I��Z�R�TH��Ӣ=�j��t፭}YC��6Mx�#3	���E�C����ے.�@ђ���$�5�Ǝ�u<��:��xp��m{�v�9��#u��wPo��պ�B��p�1*�������2?>��!�}}�#KJ�9�4�Xvf^"���?
�����Qk4
9Y����*u�@���(v�+N�A��b���6�[V�����?�_��>���^ ф��iЙ��K��EP�,
�E����ˉSb=�x�B!��:�!�j�	�M+����>�"o�]�>X�k�h���dCv6"G5�V�*=����C�Q&>�����X�h�KC���s�zSJ֌�㐣�9A髾L�W�1b������{����v����v &�
�>��f�����>; �NT�Z8D�ʡ
�
��7d�?.NL;tο2�ѩ)�p�Vy���Ӣ��a�",]���8� 98���ɗ��zL*�z!`��f-�����B4�]�yu��-U��k�y��,�U��zҩ�r�_?��y�����Y����bq�l,������s_�h,|ko���ߤtT��X��k��c^�N�?�7�S�ѓ�
��0�b'�&��}��-ԅs��*q�<s �Db�C?0"y�~�s�,C�p,U���o`/�� ����������U�F�|$5@���'��nzT9��t�C=��FT�ä�Q�0��5���u�LQ����2��-���X�x�B��B��l4rƤ�_0t�����I�b���"��ndЌ6��A���O�n7��m$\��z�B|������~�:����ͤ���d��iw�CAO�Ce*�ЬR����\K��Mg����;m�Iy�1#�xZ~O�P����@�e�����	k&r/�<���t�J�[�Ǽǲl{����_���_D�Ⓗ>Ǣw%��P6tWPRO��5��AAVs���_HL��$���sz�c�4H��*�/xC��-��$ ���V��CȄˑ��z�m��3q���k��H%����L�NO�gļ��?��(d�I����EP�9�!��.��}n���.�S�U��i���G������g����o��gP5�e�������Z��|Le����@����ꮵ#���	G����H&�b6������G�+ù|��1�
�V�ɕ>������0��K����*�g�FB`�$ι0��%B��-�#3/���q��C9�Iszá������AYO꓇j�����k�b��i6�����^��K�L�B�N�dɭ��'<f��5� �2hڏ��֗-���@��ݦSʜ�mqG��Gj�8���/���	�t����&�У��G��?�ѹ+z�)/@��}Mp\Ҽr~���iL+������)����-�a4�"�8�h�v�e�˥<й}ε:Ǘ�޴�yJq��S^o�x�|��2v��z�B��p�d�9�168���'Q��(޻���ɁT�.4�<�S���$^��8�mx&�դs��
�X�g�O�&�v2cY���ɎS�)����Wfc�:�Hρ�(��i��ڝ�K�lp��+�jӗ}�#WB��0��El��2[1�������P����g�h0������r�5�.�QN�3xWPF9W�����F�ڻP�X��{��"4����e�
] ���6��1$�ز%~�8�'��s�5�W�Dy�ToF�������;��ؘ���?}A��]d\���l�SB^��eُ��-ш�;���O����?>v�F�$���g�Bd�a����Z�g>�[��DJ��� �43'�X3������'�t	N��\�J��r Fi�5�����8a	��D���.�lZ��=/K䰂w.���̵tϬȱ�<B+�guf�a't�k��"��n��s�+K�p�v��j�O����F�*[�
�{�뇊��:,uۢ�Pp|���/0o���u�8��VV���,ً���5�}�G�/����e�N�{^�����~�i�B_
��R��W�˘����,�*-����$&Z��pQ�]-��.�"<#&*� �}7��9L�0��@��JX8y�9Rъ���<#�,��D�;:j��K}��ڍҪ ZYC����Y*I�Q�?��m)z!�>@���5f�I�Ɨa4W`e
���!94���s�@	Rt2cU�1�#7� �Ӣ��h���� -�x��4-�'�z�]O t����,����sO�Wd�<�l�/̪�)? ��̆�*l���5�DF�!����Ʋ{��l
r��d�~�˫Ю�a�F���d��b������~��s�N�u�?��