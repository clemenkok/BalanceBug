��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�!��
��%Y l�׾�m�F��������2�p�D�����W7��i��ߊ���3�%���,mn�rPp�s\��h�|#%hGd�&@ ������M褏l�#%��[������?m����������;��/qd�Tmm�S|�'��M[��V��=!�l�D���"�c�%%��t��b�"�A�����;����p��Z;�ԙ��{["~���@�
+�Hݢ��cF���,
�Z�I��D��[�#��հ�o1�Ä6��;��~���r�i&��*tVR��tt������:�c)Yk~d���o�g_ quP�9�jt?�� �')��A�Y�ȰD����1��I�Y5�ʅX��T7)���Ɣ��/ա��!���nq$���4��Ҟ�`�@t�l]aj��V٣S��a�ٕ�����Y�T��?AZWߜH�C�^�oz�)Qby�%g��'&9�9 c�@�z�����2�1Vc ����Ry�q7s��Ƞ�2^p���7D*w쉁��%�N����Lp��L��(D�����q�8h�� �|E@;�u㳖��)v	���.�\*#-���a��Z�V�#A�*�$#��:����P���V�)�(�B�ni���!gCU�7��3���Ě�����vx���ݸ��F���*��?�d6	<���Nls	T��n9�mN�L���n��T�xg���S#���	���4nw�hq�5�B�ʡ&�	�m���A���T^��Ku����x�Ͱ)����ɂ=����7��E��D..��	��@Ԛ�"*�wxBe��/�h� l��g�
'%��aӤ�G��H1�}b��8!V�~e�>S#c$���?d�L����p�2�f��|$��&��;9�f��֯3�_�����t�ϐ�3�`8�8��Hŕ�,�E��#;���������O�(�L�7Bw|��ܦ�'��y�,[�M�l)2����u?�/�.
=(��u�,	�s�m����ߒRXۊ�B��<b�7��B̑��3�}Z��/���|h�Z������������!�Jr���r"v\J]���5�qp����i���|���j�z��\�#�o������d8�-��MІ�V6�2<?�l�'M�O^���ʇkZr�w՝���OS�E�����G���Շ�ٽ�����#�"h��xO����dGK�htC��\�-�+\�Usɝl�Ψ_��5\�q��L@�%��Lb���K��oE��¸r��d?$�]Fu��i���E��^ﹶ�+�����KI��� ��4JA�EU��m����x�H�j,ɲY��/�|_�慆]�T3�C~��� Tv"��A�z�P3{ݟ	��`��$�<|� ����k0Vnآ��~qX��ߙ�=˗���M���h���r�%� K�z��I� ��SƎ��+@�V��7���~��
ެ⯊�b&�6�J��er�FSs��)CX�����a�@��*��m����]�&����j;`2"[���P��&�	-��^�i��ie�p�:�:>p!���<���S� ��#�Sd��INR掌��+��[�X�A�ɦj��\�5 8��'s;3n}цݞ�)��#BŒo<���X�&[8����Eݭ1=+��&�W��w�b�»$����
l͇�A������y2r�E�T�Q�����8��$_/�7)п�Xw��6���m��J�m͊����T�D@�+ET�ir&=��p�PC^��e	����W1'��O&��1R���*����:��ZFx�m$ˁa�0d��%ܞ̢�X����֪Ӽ�à�%��f�Q��IH`
B��P��5�89�} �s�����8:x��'#(����'�8�.o��r̢�{|������"t�w8�}mks���q��/nO�A&�$I�f,�f �q�3��λ��eƽm��&DK�b]2s��V`	w'B>�A���dYc�3��i4y0_��}�n�E��RX���Vu�'1m��Q�i7-���M�2��6�=���P����V�@DMA)`�����ʶ;|��z�VK� 9C��Ȳ��RYnhq2���-^[��?z�`:���Z}}="�_����V��ݷ�|f�K�F�<�S{7tw��������뇊�g��
�@m	�փ��xp�����oʋtR����L��ʲ�J�/Wׁ~>�����BީN��g���q�1M�I��s'O���r@�wtJ}��d���ڋ֚�ӲD��%��[�}BT:^x�g����e�[c9�:T��~�7�G{lZC�bW#&-s���u�-"��ܠ�i�},��R�ŪI�1�?�C!����P�Gg���2�T x�0��M�gz?�e I�4���0�=̱���{:RXn�k�wÎ�[�-���c�'P#��)G�7t7�\M�H�!zW�ja3��+��;�p)�R���������DB�@)�W.;~��\����ty��	��P͋&{�H�]��C�BY)ħ�}v*O?�$�Г��<�1P�g�h�9s��$v�?����O���L����tM�ԑ��NZ )���~E�D)D=匔9����x�	a��je16�O�A�SW�(�9_��=ޙ���gL���
N����֔������	�V��0�m�[�꣖������}R�݉�����,�^q#B)���}��$���U�}{�j��7��W�O�pΣR�|S�Ҡ���7��Y�/X�����~�:S�A����#M7a��2ߜx�湒�R�� �q>����9�:����Z��E����ל��~�vTn ���ޘ�~T!��b��/���D0C�O�I�$[;�B�t;E��:��+ۑ�����[J�(`���s�����i~�c�S^��Id�c��c�RM��&qK"�]�5�w�݉�ȴ����n�	@d�{t:,���Y��J"B	x��k�Gq��Ǫ`)�R��3��J�D���1�&i��B��␾�U��|��>]p���'�k����}I�,lg��R.��2�O�);'�!Q���AX|{|���U�Q�#��I���c\ת,{�\�|ϕ��1��_�;�	�>�-�A�ds�G:��x{��!acR�g��씱�|���l$y������D���$��!E��*-�7��veS�]P�����ܬn/��)�Qp;�<kȰ�#���V�q[��Q�c��엗퐲�FP����h�L����l< MaT�3G�ʌ�C"7�@K��'DRh�$�6�KԐt&�OD�*r�;��&2ѐ1N�#,�v����%���ņ'�s��<{Y��Ύ/�����Q�}�����[���3������xqz�W�}�ܑ=�M,��@\b�+$��Au�Z���L��;K���dz�:�KDQz;<�B`8i�(�a1h�����{�Z3-7���j��m���<���[,a�ݱ��~k I���1�m�����l��ғ��4q�[T�i�#Jlذ�Iv/�}��VCjX�OYs�,U?*��+-$d�͉$��q"܇��k��ػ��*��Ьe2c���
y�<�����F@G �U�fᑊ�H9�(������[�yC@�k�#�L�����Gm��Z��慈v�jZ�mR��]^��G.�<�Y��o-B�gȽm-<�r�iXI(ۈ�Ô�P̚�n���\J�1`��m�ē`?(2T~��[G����x��6�*��ڠ�X�l=%�9m�\�n������;H�GD�Z�����7[	�$�ȵ%a� Qۻc&�l�֤�E��fP��¦��*��
��&�	�ˑ5�ߺ�� ~ A�H*������^W��5.xL���FhXF����zȿ����H���F��c	��%j�&����J&����C�UQ�b�5��E_罕=��*�*4F(��W�ê��TY�^�`#(�w&}ǒVLK�2����;�u���C�_��P�;,(bK>��Zw���¯���� l8�2{��נ�Pȓ^e�.s�-=b���|���K�	�ͮX>?�c�
�I������'�kϝ>J�� �3?-��)'�p~j����W⍚!B�'"x�a�ӗ&>a�;U�NZ�A����Q�ډ���˄���)�חۺY��Ә��b}�����JT9w?�%2��`�ُ[�R�RH�n�U�%ޤa�ldr<�H0h�㰉��O�	��?�O@�6;4�L8bV��Nq�w�=�v}2w���3Y���_^�*�=Sھv���`�#��j���'*��?Fp�M���0G}�aKR�/����zs;��W�Y쥦�E��O��P~6,Њ���(��%z3���]5�i�(�P�d,�R�^�[�w@�K�'�ث�,�I�a(�ǲ�t�6W�s�JΎ��pN�	[��E��[FV������\�������A���MFhN��2�J
�.��*aչ�~(���ĠVp�Ô���������Z�����U)N�\ ���X�9Y�n��=I��9;O��pc����|�� ��Of�,�R��B�� T�0۬��g��@���*7��R����
7�F��&����J�G�R��ۖ�y�BT�ך���(��X��Gsf��G�V0���D���
zȨ��I񳀐�JT�ԣ@�ѻ�t�7Q�� r�;��3x�B����x��0�"�3R�o Dnl#&u� �x��E��)��A9�,�O:UDGK�W+za��J:ĻAt�<�[,��Üg5��n��`$���sع�|�E�E�x�������j���P�����HPQ��8f�̇X[�=`9c3rONg�ȸ�B)�nF�e���X���W6����Ć���?�)oB1�����[�&�{���j��a� W�_M�Ia�R�^��l�����H�̾SSN&����r+,Ih�=�Hu��I-�3�|��ꢘ�\A��{�J��Ă)�o�����b�~wl�X�y?�NaW�t`Uc]ܛ_�$��G<�1�tb���9qc0�6+
3��V�����5bC$!խ���QI�)��[&Ee�'���6�u"Ϭq�$9H�3��"}�o�2n����,l�\P��π�L���6��-���c��6�%NL�x�?�g2�f?RP�acX>��+�G�V�쒚8>�bQr_yM�w�OvQ�(W��h��#��n:xhSZE���P��'=,i�c!a�Gu����W�D��$�d'�L5\�_��>K���%��w��C��8���ވ��ߥ�5�����٢^�J"��1*����y%���ln?���� �B<��d���Tј��\��{�g��2Q���x���SV����<�ءx|s5���1eh9���S���pS��͜����Y��¹���&�>�-�\w���|��B���L��1� �OGΑ]�?��]x��	��A�Զm�����i��!^���rΪ�>Ԏ�ƻR�9��&.����@*����I�e�k���WO9�uN�ZȬ�l��6���!xُ��)o�r�4�ء�TZdeq�꼕��? R9���L(e�5��{)G�.1�ft�yN'�����pA+�/�����O��vYr:��� #�2�9�uQQԡ�5Dў+��T�(��	����j���q������&����-�92IM��`��k����Å+�%�c%��qJƂ��g0�:�,�OT��_x���cl�¨�!�0�d�7/�(���$��R��z(G!mLc�r��^H��[A�*<�'��#��;�Dl|""�6QI�/�S�i��os<bҔ�p���X����u���6���I��$�:D����c͒5N��[ϠT��j��Qj��X<6���r��[[�zpd!��y�`X|�rk�?��펮���7�H�%K8��n����/l���`y�F�
eb�Hg�QK��qfX(4�"�yA��hPz�4ޘE�2�=.W
-��Է��6N�M]c�n��Z��84�e����gr�I���"�,Қ^2Y�T��^��G��ՑD2��Z���%k��=w)���nv�r��ᵛ�)Z
��i�(@l����zS=l�)� �0l�9@r.�i�A�F~��V���V;9,1�Ǡ��ǡlz�X}�O|�-��8O?�g��b���8�I�A��H�� �"f��#�[��R�G���\"��t�3��0��1�ZH�8��K�}�	T!T�sW�y?�iٶ���>^E�x�w`U{��=�!;rHЪ}�{~'��I�c�%�!��6����僱z5��
p>��$�hz��%[Jҩ�>l����!��6��3G�G����Z^c<��^��g\�<�X }ROR���).��@/�����)M@R;��I2(sfʉ�<m���"�\�K8��]:(&���bi{n[��E_�c2�K�'��Cl�*��:��G��g����������M.`�̍�	�o�~;��<�!���k̉�i�b����+6W�����sWg<ub�_f$�"ᵁu���4�L"'�D�z�&U��>��p�'��yh��"��7�4������wQ[ȷ��!���l4c̯,Cݓ�?BzU�M��pN
�y�v����Q���\��A�6j%u��FW��W��@W�h�ER�;!2嚅�=�u�|,1K�1)ֻ�jܩy�Ո3���z���	m��z&"Ƙ�L��l���垗t���d�6�x��u,��ba������X��Mع����"��~�')�&D1^�e)���G����ȏ����p��~gzoo�Jcp"J���s<Hd�<}p�q���]��礶�d�Sw��!��d9x����oH�BV0���D���pɔ	e9ۢY���oP�&�d+�ź-�J��ԓkahI�N<\��ex��}� ��؅�{"�o��6�r6���e
-�.�KD�D�{�����-v����ɥ �޾G?��l�;w�g�Ϥ�Ԭ���܀t�lZv����#y�1Ζ��������(��D��6�C�z�o���L�R=�O��>/��&�\��
�"b_YH�����Ty��	��	!����S_��'?��W�r��sQ^PA�?7�Ap;��B��dL??s��}����+$��@��D�v.tƌ�d�Z
�%�����V���GV�>���N��*4�Z��=�Gx���"*ƙ ��.P��Cԛ��=h�`�٣Ze�����z>�ȕ@�"���U�&ڨ��X0�N;���@�:L
a*���b���rI�3��$�?��z�L.4�1/~�~������Y��\�ϟ����P����B
��?�>m4��_��p�����}Q?+ Wd� \����|^�����:|TJ��i�d����x�/g%H��Rb�qS0��o>�=�<.��:DBMPoh���b��}7Ye���rVGy�8ڥ��p�]��*T�d+�֨fX3�֛N�H���%�WO��0^{y^����-�@�k��d7�����0���B}��]���h�3�@���/�ݧ������6ݶ}%*����c��Z�4�9�ѳNr*���T��Hn�����`þ��r��`�Ih�(@�u][�l��1���ܠ��Dm����Y��E�W+p�*�i �ב���_).t�ӧΨ�X�NS�_�@���RCK���0|^�dY�V7��v{�8�U����#e0��勢�G7�y9�Ȏ\5�xC�ȍQϱ�e�f�V�G�������	2[Ƚ+����=�2$.��Qb��-%���= J�!BH˾R�c�>-��t��v�0З����R����$�T�D�Ƕ�.Fup�|�B�����h�ߑ� ���I��\�#|E,���z"�JJ��L��� ����q�3���~�r��)��k�Q�C1f
J�$���*k��P.���d �{_�L�tx`�(�@���!󼰛�����Br���.<^O�G�q��\�p��*��^�.F�o���>!�=uZ
 �v��'��|�&�ӓT���4Hb5�wr�E��J	�e�{�h'��*!~�2�JV�R�&�E>���]�����Ϸ�?���7ĥ���Y����������K�@�[���$
���� �NkN�"�&�!��mT�2xq�Oյ������[�=�t�fY����m\?c�P�5HSy��?�<_1)����'�Z��7y�;�.�rG���=�20�u5iI�Ñ�cok��+,�84Mf�p��=
�(@�: ���ǽss�c8�	//y�7%��1S@Ў����
��\zX<$�L��@��a/��$EC����s0��|S�S�?7����������%t������|�( ߊ;;��bd}ݜ�!���|)�|�p 1W׏�� 0Fr���H�۵��Ȭq���^:�&=#��/̨�.��<��`���6��&* ׀�.�1O��gBJj�g]���3U���n)(�Cҷ(������^����Ӽ���9�#r��g�C�������B����u�{�3e��W�gw�M����.�<��{��2�fa"�ml�1�^�t<ҩ�!)"<ס�Vg����(3[u��3�o(&�|�9�K�1dƝ�N��?�GP�?�@@ն��K���ܔ�ҿ=�#�fF�Mc�U,�U��'�H�>��.����|��'{@y�ܚ��)�����e04���paBzp��Kj��:(���"���`[��q�1ED��$���l��^i�j�|�
�ĴX9�1@S�쇃7�_ab ~�u�L�(&�VXO��`��|��e:��"���!3L0�g�~�Q�	�z����i?͞���Y`�$���&Z�2O���x?����X��G����l�I[2R�Q?�i�4�isw��S)O��-�Y�4�Ȝp�o� �v!k��Z�3mͬV�2`ʂM������
��)�֡��qVJ?��"����|�4M��D���������)�\�e��B�VQpM�$tߗ.,M�(��B(��ү�	�kqWDTMG��Ȍ����@}J�ڲ��;��r��	�.�b��X�}��z91��D��hHQ�8@у�v˺	mX��*���d��n�k�\5ks���1��ϋ��U���@��i�������tn��0.�@�?�T'�i���H:�Z)&3��ES[B���p�t|�%����/��r
������R�`e2w��%J:�Df��	��hL��t�դ:�Ҙ�'*Z��d�a�灾(��5��W�L���o$� 6p8ؒ9������i����U	ƅ�1h�t����՜�il<-߉gq�v:��K�a�`�'���O�%bUNf��$+�\-T+�:n����;>��:"GZc�6ڧ��cJ�>���$X��5��=���Ȁo6D^��I�6i� I���C�:~�4χ���ٸk[N2=_:��UB>�����6�� Y��y���|B�R! �8�L%�K.	˗oX�ysw���5��)=O�Y'>�Sg�O0/q6�u ��C�b�:GI�{눙u|�G����x�8Ţ�ﭽ263clh�����v
dtx��#�]�'ҫ0N����O�<sj�%1Ld�����G/�t%C��H�\i�A3��aaxIN�	A�xV�gW����LA�&����Yl4{޻�����P�E�j������F�G[�'5�Mw�FxH`9w�ｋĳ?�c��Y^�f2��+V�=Ez���(�v�D*W 
рA fg|g���x0���:b���k�i��aO̶G3e����Q�P�6=`�7ݩ·w��d�Md�J�ET�{8Ha��v�����D>Po��QMeь�b&@����ߜVXW�<#���pۮM�GSWJ�4W��F+�d`4]ƹ���aqJ���`��9."q�	D��	��[5	���Vh��b�~���*����]�~]�e�_�������{��^�ihQ����x���Z����x�rTm8|��+ز��Q:��AZ�G�2_�ȓ�7s�L <Ⰳ(�LA(�AmIGʖ���x�6�H��q< q�����9�jU$J ��G��?�;G��&QU�n|�a��ˊ���B�֙�޹/k>��pݬ��^c����jKR@~�C������/�ZX�`*UE4%��M VQ,�w)u܌}��i|}�L�L6��iY��&h������� Q��&�ܚ��d/h������6�1��(<�|zZ��`��0�aR�+�
�O(�B�'#�;�h|J%�.%�� }AM�,�+���Y*�d�
�At�� ����x�#��w�s�ײ}�u���|ͿD#��$��d���-g�0`o�)VĪn����	�ɽ�/�m�����f\��
����5�ƶv�	��-r�'���Zr�=�j5"OF����z��A�ސ����gm!+�MA�Uִ���AC2����)�6�z'�θ�X4a��Jd[�
��B� >�������r*�.��aiib�Ǖ�ĩv��ae���!�s׸��[��Þx�[�*U�U?���S3��i"Ss�{R%+�����`U�`R�8} ����߮����,Ċ���$u��0�W�,���KQ�����/�Aj��{e.A�Q�Q.��X�����S;��i���
��{���1ẖ@�O���i��0�(I�,H!���8���SoD��	�<��A:����͌8z�)���|?J��qN0�~R�/�"U�;FP�$d�ƅ�Q���];
���f=�'���/!R^^��1U�&�eʇ]����N���B4����
��k��ϙC��XW�O?���b��>�܋�X-�����U F�;hY��M��pз8���S�p(e3�]}F�ybb���$�~7 ��>��ǣU@�45�
��?���:�O����^ ����[��֩3�Dx�,g�稜��o3o3�CTQ�^�<l�3e�A<jD��;��דX�Ka�g-���R�L�Ͷ�x�͗�[��m\x�	
��$"O��R�`�g \�z���o���l�/�أ���ZY���0&���ˌe��!��+R�RUe#��.3��"��!������s���d:s6��cO��TPwS���l[�?�l� ѵ�D�Q��4:�l�����5��|��e,3|�*T�)�d��SD�����-�7���)T�OE����HR����b%{v�Q��i^H�}�����y��IN���/�#���֐�-Ҭ%r	��z7��㎥;I�6Q`&�`��&I�)Ҙ�>��s�:�Y�n�an�[鐒h���Z0�8l�t�t�]k���#1���ui_s���hηS�Z�x���Hϑ���r�=�fJ��[5Ѷܔn�e�Mnp��\��T��O�/�y��^D����u�2�����HnxK��p<����F����~ + f�'T�6�Kb��c���-?��o/�a�3DB:��+��)����Cc�SԦ
��Uu�N"y� %�Vw�Iu���e�%N��#{�c��T<0��#:��0Y��t�&�,[���5"r�it���q]�'��Fb�^������{��9���`�=��}|�& Ig��˞a'>,�w��6:�z �5�ю~���z�+���I�p�Ů���J��d(9A�7Gpg!i�/E[CL�U�˝��X��l�zx�̏������!_�+�3V��5k�7hO�V�$zM�_���#�"������-����}/#-�r�E����
?5Kί�b�ɼh��~;#I`j���nW�X�{��:w��'3��R}�}ɜ;�>I��I���]����q�:���0��f\����/.~\��0`3ѵl�'
?���lA��d������)9���㘽��P��z��S/E�H[4-�O�~���ޯv��M�V��7�\�W;�OI�N��-A�0�������)�r$\�ޗ>ˉ���8$Y���7i��b�^��7�)�O�i35!	�C�z��!'3�UE�����ڤ����M�b� w��41_K?�8�G�꽺�%8��Y,��Y��{,(���O�,a7%M��q�p/�0��]Qϗ8��W8�n֪�:��s`c g��� � �!'��|q���6��;ۆx��U��h�N����p�A3!�����!L`�0D������h��q���:ݣ��_el�y�S���r@�~��-BE��}���zL�4�D\�)C;b��U��˽�#��zlG���k�����m�W8��]�-�^�&��� �J���.zc��|/��b4)����I��k�J^}aqߦӰP��X#t� ��V�]_"�}' �4lc^�HC��g}��s��	7l�̭S&��W�j�)�W��y��7�������^��/���@��!ö�Yh���[	]w��!K�k_��3`���X2 T#=�?����3�~o?0��)�ݳP;��m~C'�M�f�~���J�D��e���:W4��g����h����MD�NȺ�&�3��Aa֦��K�xU� ��e8���A�+�G���E��o�\�ʘ<M�ɫ�1�"U /��+�mR�+!-��_�h��C��[,�ق2�*a4�B���C�[��E7����߬�,*}����z�C/��q0�����H�`��.��w�ޕ��b�t!��/�Şg`�����!����X���[�y�|'�ha�;/�%f�M4I������m�W�>������R#��0�����	�di襏#Ǽ�� �i:����kWI���[���5�Eߛ��Z�k�Lk$�[v����Bg�uZ��nW�AIࢬE -oq�z�h��|K/aG�E�K�'�}
��NC�|��?��^���q!��������OZXJ|
�ƨz��r8�:�������u��q�QT�:n�芇��)а�]em�2=��Sl�p>6�C��n��fgݣhBؼwiQ`�@|p��:�}²v�}2IL:g�����P��C%H��$Q�U��
�B�0���:2(���4�B�l,%�4y�H��/lXѹ�-�!��Pc�*W�NÏ��1�:
|�3�&��]g̫��=����Y���u�9ΉO�ͩ��@�ï;5�~S6��X:�ߕ1��5��P�O�������	+�G�&�ia���v�~��e٦�����s=Jgl峡��Vd�����7�~y�
���Xv���d�z���E���*E�ӂ��9o4qf�M�}U�j�M"Ko[��]�D����r�-wNS�\�7O'Ҟ�������ȸ�Ë�]�' b�Xz��kWX��jZ�̥�^L�����l���ḧ́�6�����S:z��Æ�1dW8$T�OiС����J ��5�'Rk��s�ov�$�s0�Ġʁ.�ߵ�-C��L`�e�Q��<�P�H֌�uW�f�!����o/a��n�ǣg�I:HƿL�n�oWƺob���8���V�,zO_��K ��J���/W��#aB��C�� ��:؟1o!�t2��E(:�S�W��Rb7�e�1�8�{�5s�O�o0�ܣ'B;܊X�O}{���W�c�φX��7�\m��D�"}�[�d�����-~sl��I.ז�I~��o�S-���	q� 
��|c�ѹ^/�8��3��J	
m�L�ΐh�ZA���N��j�N�xK3�	S�iߨ֚n�X&�o�_E�L�>K�-m�{}���_d��<y���<�aa��+E�>ُ�L���߅�k�	ˣWIp1�Wy�@߷Co����O�[�w���'.��K'9};��u��1G"����z�Y�	�mC�#�@#0ۙz������{�	m�7���Wpy����
[��4,��
��|�� �6K���(���(�+�N4�=���r�R�_�=�:BI9ljU8����\T�ǳ��K{V"�<�p��+��9l�W`����3*9|J��5o��[e�<-#Ոs���<չ��LQ��?!V�'k�=��|m�:���??3���8=!���L;�&`����FJ;���l��Ś�X���c��d_i��dt���/V����r΄͐�Kkȳ��d�R�a�&>��l}��1Ɖ����[w��G1:<2���&j��kI+5bԸ�4*�\����n+=�&D���>�Oe�OT=k�f�����As@��d5c����*1%Q	�T��vnj�T8���o���O�;��*Yu���D6�'V]��t�DX@�����X���rTǋ����3�v�@|d�B�hH`_e���fP.}2Ɲ�β����9����jN�1b���B\a��n�8O�6˓@�*[R��9}��&U���o�5�C�l�l���4�LxW������i餽�	��:ܾo���kCqD��x�>�*�{�͇m�r��g�V�0~�-���f���>�ݿC��R#��F�+�K${B퍋Z��U���C9�d��&�=1�H'ׅJ�QD0�1vUgj�ny�B[�eu�� ��׹�03b������p%
�-�f��54v����t�i������}bt���i̱�2�O��j �B��*6x��8��F!��i��H�S�޷p�d���sn>�l7>5u�AM�-V��[:�� Q�wP���1�R:��=5��m�[줂�� ��+��O��p���j6�펪
�����9����0�����{�Go\{�Jw��&�UҸ���-e_�(��J�����p��f3�f�-r��̘�Q|JLdR���[#����ti����"-�
�v���j�y�֝C��.�u�Á�;���ɰ�s��)�Oc�|���ַ��>�3�C��;h��֪�\8R�@�T"����>^�P07���Q�Cü�����q���-�,p�W�{2w�Oj@��[&4ˈ�z$��d���\S�B����|��u� k���>q������4qֵ� K/=���O��T��:�P4l_��l�6Cڍ�;uF�qB�z%ɗ�o�D�h������.�o����Z
�d�F��Yv�}��k ���$����y��� ��ir�+���Fs%l,w^f�����L�Us�8��nW��6�KŰ���o���m��3Ld���-��f�G��ݨ�]Ŵ�]/�2�78���I�5�G�ArM,��k?��rOZ�Ř���o�͟�O_��0чF�@/�65���0_�ޑJ$<�!�/N���2�`I��Ǯ�����߫ں��#I�MB��\~��:5�f��-��(̯�=�ޞ��h(Bx{=6��#qz���
�6Φ���!V�=e�'*�^^!��+;���Z�l�/�Hd���&�?tc��~�6���tq`ԙw�c@�b!;{n�Ra�P����J�{���O�z�\�2�Iϟr^G%���|��e����X���L�y���h9���]Ll1Q��"B�>.�B`?�n���H{/К.բ�P|Rr������H�?��F��W��`~�H�Ug����7�Ki	s;��l�B�5�ux/��7+<��o[��,�C�dw�/�#��ᬒՓ��I���Z�/,4�����ĸ�h1�ΛpA]l�D]�z�0��hl�y�U��_y��C���~ڍU�Tԭj��f���F���[��iOBuX�gO�.��pl�%W�O��s�=�u�`]��:��O7^/`���P���7�t��{~�����ܸ��, QJ�Y1�膏uò�8
��[
�Q�pk�+�d� =���!fE��c���T/ ��M=�R�g�۸��	�]���o����sf�jЌe�O���Z�����6��8�7�ie]�q�~H�0!���X��.7� ��$���hQw�|7e�:ӘI��Y��?M��J(FX��w�V�l����`_cO�c7A�W�)t0?����4��ۉi���Q���������Ϙ���c�č�L�QI)(��A}u�s�w�XʋGn.�1y���b���R���7��߉A>aCρx� �}Y���w��\(�/�~cI߅�%UV���J{���hVM������#���Ԓ�R����"B�5o��x�o)Փҭ��ts��}UH�B�C1����=IA��x�fK#�AS�d���KF�2��5��>~0�0�+ÄmO���̚L�y��+ *m�!����Ot{�(�� d�tk6�QE4qsnX>�֥#��E�=	#�(�G�L:�������;Gzp�)p7��߾<=RE�e0�5B�Ҡ��Ϊ$�h>�8!��d��kV@�~K��r�L�<��g�s�W�����4�F�&v~ut<��¹Ƙ���;+����Bg��ၩ��@O���R��u�G�{�Y�!��+��e՛�:O�y��#Y��{Ht]9��Tq�Ɉ��;�R�����+�$��qP5���Z�,m𪋖�/j�i.����TF����8/f/�n�]�2|�}��
f\�0��21��"r���D��&!�م���J��`�y;$*��!=�؊��Ζ�6 V�1����R����f3<��i��{�L�7�R$�8V��?@�%�n�\AV�YU�]�'��`�w����d2�!��K�Ư��F��W{��=}ڥ�
����9VL(F�(�բ�d5��Q�hӆ��(�X0���z��E����U��(Z��R'�_�j���],?�����3�,1�?9Ҵu��*K����V�u`X��G���R��`�<@�!Jv���a�qq���/#�u��L~}bo�%��'>?���i�J�+��M	/���8�?n�5��4HN��{�Ճ�%�*�hq��ھ@�bT�r=���6?r���i�oʥ Wpe��̰p��n��i��ω���@��um���`֢��M��%!���ND�C���s�s?�����V�~0LKs &$2	C�W��^�
{*ϵ���fw'����$?��	�Y�nb�,^螟���?�Ԏ�$ �%!�r�=i�V�$�g��{���䀾�����V	��=�솜�6j�?�e෮'�)Jq峟O!θ;E(��/"���-���`�Y�Š"� ��`���x��,��#]l7�P���Qo��'>���R�����~�[7KMW�#�ě���>H��ܬҗ���
��&��n\$�f��S�c�Bu`%�q�{�����@�/�ϊՄ��ѐ���U�7�ҴPX� 䳑 O�����3�<��|У����EBSZ���	��1�-˜6t�(���vҵ�,t����E�X1UTD�#'�;~A��r�</����aj���<4��7�����:Ҩ�8�p�-��{�5`0�3�-Y�~rf��	m�-�{��M���{ѶA��� m?A�tz)U �-���U��O�fkD�Z�~���@�����7'�Er����X���֨�a�����2nB�@�xu^���X�v���@��]~V
"U����=�vw;J���m+Pu�D7��?^��م�Ts�V�R�������~LV,�A�E�~����3�����n�Dp�/T�gBq��4�,�!���Z��8�`�R@4� =���W�Fw�6�CRTܴ�!�yL��4�� ��B���rD���Ŗ��j�Y�܈�����"װ-'b�uO����~�n����AC�bAuV�od��ͧhN "�EW&�� }���&ʾb�!n�x]���S`b����0ݲc��f���yǬ؋��|;�����:�����X�8OQ�Iy{A_��`�r�C#�~r��)��IY�	M
t�ʷ�R���p�ď�m��7�Y����qVůgD$F�y�� �ץ�N䨤�l����p��-�9��tU�e�IQ�Z���+�PB$��y���L��7]��u
҉n2��L$|�
A1<�M7@��b��fk'#�\�aK��ب�Yƀ�R�Z�E���a�8��(��Mb��m���H����|�T���nT9�m��D���qݏ�
&�z͝׵�wh��A�Iʀ���ޙ�J�ei��cWFr�*|t�@��65����y���pXs�N�oCrM_�-sv�gV��-I�/9z��w�����T�%)i_�s��z���{��
	MM4��H�i7a8a��ap���7g�ceB��ƽzP`2U�"��_�K>}xz�LZ�M�5d!�Kר���P�/c%�̽R�FR�/襮��j���GLM�	@���M�ؕ7��6����k���)���!^�x���Q9�(on�W�r8���eh����IC��/��
�џK��^�B��(~>l���ƚ�(I��z���ѱԋ+.Ǆ�D�+�#}��J�I���z��11M�쵤�KbR��)՚�v��xoK��l�b_�xB����M%!q|��x�ܢؗ���[F�2d�+$m�ަf��u~x�t�I����J��/ѹ�O���bXYej��1��:d�+O����ȋ���~���~Ʃ���H�NP/����pQ�l�f(�].��G�o�={�m-[��G��X�^�����/C�/�/��c����b5�Q�2�kc���0�pFX�C��}T.�(��o�L����{�����g��Rn!�<�C�'a<�f2V+!6}��Or��/�_�Z��č���O1����T�A�_���$|�
oV
u�����*�>6���)$?\��U"�3"�8��̳�oRg]�)�> ��eJ,gN�6�{r�lĬt|���!�
w�X��n�U����Vs�3�|<����?Vy�lwV�u��X�=�m?(���fv�:z��=(����������w�� ΂q
e��rG�v�Y�q'�A;��t���� {�'�/f$���y�oJ8KD����Di��jJ;O���X7�y�3���1a'�T(K���A�< tr�H�ߢ��D�l�I���c���G4Q���c�l��� k��K#
�"n*V���
@�Ap�����r�H�V�,;����r��p'QLX!�@ۡ��$�qe���f�m��7�F�nV(©��!8��L�w�z�9C��[�k7�J�̳,�,ZE�9z�q�R�'��F�)���727��B}i����n
���v�.q�{�)qE0��Zұ�%��$~�D�B5���_,����_Z&c��H?�qFdyj"�&������6�~S���q�JJ�fjA�z�)Dg7�UT/fdF�ȡ\��ߴ5��=�ft�QO�����P�}��Ez�m��^�'a-�%(Y��1Td��&>���3T��CY~5[�u�j7����N9��'�A�$��j����m��@���J(�H��MI;����F�=��N *Ħ�HK�f0��K-�n�p�b��U���<7T��ћu��e������|�~ed��~\����gLxĹSW����x��)'x�ȡ���+Ʃ�9�K��c���)ӥp�5���ذ��:�m�{��C��.J�?;�m[��3�leH�����Py��N�K'��T�(�/�E���yËj�ݞHG!	��޻n��a�ې���s��R�tR��z��rL3&U��۸�V�u�{��5�]�]�:`x��yZ����p��g�a�oU������:`Q<�\f��f[��n$�DI݌[��?���v)��?�?��lGhު�ZFelR{Qvέb�A��|kR�S�i=�|�A	��S2E�[�O>K��_���B��>3��Bd�k���I<�瑏����xz&�a���
�%�H�i����9���O�nm��pgA����Z�/;q��IC�%n���vg�a����'����r���˴�핧-ٷ��,�0A#�3{���A�ؐ�9h-"r��1m����_u���3ƪ��]�EŶY�Y���5��#�+E��Y�#�@�m����d���|.vG`�ȓ���G.S�����BB��p��1�/b\yށWAIO�ȚV"4��>Ĺ]F�+��}"Ec�|�-�Qc�ӕ;JN;̌Nn"�P(O�'��SQ��k­S�l%%����a3��#9�=�:�t�(��VZ�݅�͟&ak/䋾t�M�H�T��Re`kk[e��1#�(W��%��e�3�t�/�!��J��β�!�J.g�BiM�5r���>�K�)��sr�x�hB�Ѡ%A�;���:_Aa�O��0�r2�E|;jV���+@���E�y��e��bDP��B�d�E���x�7B������#�$�7YN�=P����ՠg����Yb�{��1�`������e��sgE��w���UV�7Vϼs2VF"�LSs���4�u��� ���"�9�s�+g{���A��M�lo���6ۡH�����u1΋���3K���iV�#�l�k�*0���BI��8Y�,�ˠ�x�0�ဓJ�s��L�B'�9�P�'�JW;j���|���ѐvI�"8��>����4/fS����@��n�Bc����=����i�jҩ�p@dgm6h��_N
#l�ɩ�I%&�J�Ӣ`��i��V�{�� y;�:�~�Dt��HA|�Z&�o0��� �y�mzGk��pK<u��g��`p�
�Exb�f��w�T�-FsI�k�R��(��O�Dp�	��Jջ�8Ϳ���=��B�k�g��B-���.Ә��?��Q�x��H v[q�	[j���~d�L�
�
�a]���_趔�>��R�h�:^�dl0�̜�Zn��}�!X@D��r�'�~f���@�zi9i�L��r?$������
G��q0�d���,�%(�������.�?5
�}�?������~���=��r��OQ��O��s��h�6s���bY_5�u��_�V),��9���|Y �ȁ��L��A/v������ f�����=Y#�488�W����,)�5�즮ʤ����$�*9��&�NO�g]�*)��_��.pR-[��M�^~p��F/�#�aDe�04]� j��p��� ��ZT�aK"񈏔A�l���M����qK?�!��Z��6����Z2�q���B�[��q���-�Q��94����-�;���_����,���Y]]��;��ukR-�`ے�{�S�W�*�ԨxRD�G���5CM�y�e7�����按��\OĠ%u��T����9�|b��,'�э þ�x<��K�%)OP�48Y�*x;n�\{h�����R ��%v~z�iC�P�WM9���a8�{�<:@ڌs��!��YNs�&��c%�>�_x���9ґ�8��)	�?�eB-J��uu���~�f�l�����Q|,�yPh��O��4�=�t�����ԧ�zˉ�/�n3�Ρ!������T����8�y�f��X�mZa5�*����q�lnd[���V�3����|ט$Fl�@��-�|�s\�`p�Xw�x挭L5JF>đd����dh�6h������Dٔ3�w���ݐ��`Bx@�yy\�2g�V���@���Y�����h	�xJ=�\�~@{����uV�E��9R��#(��­��&w0&pP�3����1�����]L���T�s�py� ���!�-#C�+���rO�����,}�1���u7a�Tg��,�P���Ǆ��j�� o���5Fwf�À�e�Oja�j*0�h.)�>:�4>"�_�*�ZEh/W�]t���@�g�٘�Y�lYT�VC�t.���;�e"G�wv^z�'��?��K*���|T_�)3�k;�U@���L�ҩ���?�@�q�X:���~��l|;Ӈ����I}�W=R��-ۧ�Y9���a��[��Z�y�K��6�>Hx	;�@:�����2��gT�§C��5�`�	H7چEܾ�xJ4�Ϝ�|߸�rU���D�T���-U�Bw�u5��Ǆ����h��D�UD@r4��kh��:y?Sy?�ϟ�󙬔#_�T��GlX$5TA៫R@U"M�ǸE&�/�ف]�Ԯ��^*c�I�S�T�'��!�6��.�;X|Ҵ��nr�Z��1�� ;�w�=�}�åC��봸v5�(�2�$A���(��Ma���6���>ۘNC��8o#�Z�x�m�ns��c,6h��P�	R��Ûz�ƹ%%m� D�Aqb���!#a���j��Ȃ#�㭵�*d�-��:�"G���>�G-�=�_�oз2�}3�a��6O�P\�r1R�ٔhu��>����e�A� 4^&�-f��n�_���������8��Co����i�A���-���ʛ�	q�]��>�\�]*��s�*�{e;��j�TCR|it�C�V�aCˀ!�<�<����X�[��2t�2�.���Y���&D�󹧪-�Zw�̗L����6��J����:k��m{�S�Њ+�?o9-��풁u�S�4}s,�o�Д}� ��2�N�+��d`�j�3�G��ƉU� gy.��ub�*P�'lT�E&�z��b�)1]�Y�$��8`�k��k@��W����Rw`��/�Mc5��jk�@^"ҩ� �A6?V����(���+��N���B��gvK��[,�?�d�r��[b��ƛسz����N��J*�Y{�����bw(���^K|s�9����W�����"�L��T�.�s���Ah3fF�Ú�°~zj@����u���$M2{l��a53�b6ζ=�VS�6þZ;��2��L	��"�|e�i�e9�]"��*�l|��7�?(]�������"��. ��o��QS�0��Ѐo>����R��mT��x�EO�h��x����os�a�b�r����|m������䵉�nK9�!�a妣���WQK:CL������^a��[;lm�&W�ߚ�g������[����՚#�`�l�G�I��~��w�����y����R�Tm��k
��A;u�bm=�2�}1]T������1����\�ef��ʁn��[�:@h�_}�#o���0� �Ȧ�򔙉zb��Ɯ�l���������Ikh�x���U�@��p.t��<��v0�Rܓ�4ܔ�A�1k�ߠ��O��.v����u�c��&��������Б��1C�$|���O>�!z���o�����e,U-H�x�lB���7r�頚I���#"]�@K'�y�y�IF�S���p��Zgg�������b'��=q�"�;�%����v(ؘd+ϣzמ�4��!"T$G
c-Rߛٸ�lռl֏�GhNm�0����i
��tCE�ZF���Y�{>}��\�2�N6�ae%�I=�;�k��Pb2��æXٟ�i�Kkfִ���w��`�׹K<h\�<��c�q��������5$:�(^��.,$l�@D4�B|$Vj&��r��x]a�����7�.H����Z�2Fq��{$�{s)�+�4�[�"+]�8#چ�xݦ��R�Ԅ��0�M�0���̰�"���|�yn����ȸ��!0I����Hh�~P�i}���� ^�a�0�q��j���l��8p9��j����V�<�����7���ަ���n�9$IC� ��ߵ��ƣ$=������f��#&��o��dⰿ+_�z�G��-�dEKK��r�8����Y� �gQnE��W�(8�� )��\u��̑��e��(�X��6�ק��W�~Yqj;wg%q����
�l���R9ؙ$�M՟���)J�W�n�����E����3II��O��d������k�����V���?J4#��x-vG�el3-7��R-s��Z'���߾v�e��t�B-'�s�s_�c7p�kT���Z<�7��,_fk�+���:���p�^�J��j��s�:E�
x��7��#m2��pi�#�y9ΙK�wI�#�FB�Џp��j� V�cL,\\\�l��ˈ��A,��[�d\d���7Y<X]@~���-uԷ��!82�����n1 ����DZ�����}$?
nI�5��|'�áܤOIϳ�Y�IrM��i/����`�{U
�NkU��Ci�9@ˈ����{΃4)��N��â3�(�u�)52�@�:������7K�� (��{1������(z��0������������2�k5�;e����l�}��#`t�l@ջ,�N��%c��;�;bг\����.! _AE�os��]����ɭr_�h�^;����W��_���"NE�훊6�!f�����ɞB����;R�R{��O�K��^�|F�M��b�n��Ѡ�����'s���注��e�����	�v=0�P[z1[Y��b��J�#M�O ��z%��iiڨR�?�q���][k.Z�
N*���]�أ�!S�.����C�d���I�g��;��U��:τRA�Z�/�p���A�+z�%�IGG.����ke6����(�
N���aV6e����<̹���ϰ��hJi�dB����Q�4�
%�Få��mRgZe?~��m7�x�VCL \�G]BPQ���Q�g՛�<����M؛�{Ҵ[1}���j�t|��I_r��E҆�I�s%z%�
�e�A��7hQ)ƿυ-+8��܎�f�~��k�������.�!�9��k��;��O�854*�9��*w���Ċt�uz�R4#�C0���Q�MW	�>�E��D��E?�feEj�k����ܟ�r�̰j ��\�Yq��O$M�;[l~�چ�D3ϵ9V,=j�Z?r�J�k_���T�v&�=�?;�*+�j�
��=_���.�Z��j�5E��	1��,�63��Ʌ%+X��U^�Y���sJ*)��̸k�S?��T^te�m�_�ꂚl4�D�Zd�N�VwZ=@�[���f�Fy���v^�.�|L�Ĉ_-���`)"�"h� �b]B�c�T�?62�)�Tk���JJ'����+�n�&�٫��(l�r��L��wb�Az�w]������8wx�������@12��"���ݍ���=�����[����r�F���b�2�t龳���/>��Q��C!�yǥ��@��F���s�dĿ�ai}y誼���߯P��|Bs6�G�=E�'�.I���4ķn�#��3���l6~�:��\m(����j�9\p��Ce��J���w�$l4uҪ+���D��4#��Y�c��i�����_���6"�3�6��T��);I~�'�G����G�P�O%���sCz�N9Ғ&�����?SoM����FH*�cy��Z���D�Md0_4e"�d���zx���9�ڠ�	�d(�r�x���=���ɟQ�8,AG�s$��%ڝ�y���~FU����C��P��Iʣ@�K�ڳ�]��|��K��i�3�AAmk7}(Ɲ B����)�ă��y#����9�;
R>�4�D!扜g>�V�%��Ʌ�Ƹ�D�>�_v�E���/��wOh���bJ2��}vCJ�E|~o^Q�ȅ?���e��hi�t8�Vg� �9�e��!��m�E�f%t8�=�*Η~T-H<�ޏ�+���Hb
k|v�8E1!r�t���F�����`����Hj&9��(SaZ{�@8l����n׍���P��Ú��R���%�W�n�WN��^�� �(��Y5�k$3`���H��`�i�D-���Kb@�Ⲧ��d<�z��P�/S�S��1��A��Z�{/����u�\�GO�/�%��P���aN$<T���S6.�A�Ue�C�D��%��K	��
<��,ה��*v|��Ո#=)�4v�:�Z��+��DN�]0e�@�u#��>p�}ڗ)i�)��gA�f�F���@��V����L�ov�����_�O��ޚ0:���O:3�"d �|ݱq�Da[ǨV[ܴbz�<���`ߑs����Jڇ�ۉ1U�v��ѠdΗd֕G7�c�Ɣ�d_�2��SXz��/&���Zl�EB��[��X1mط��(s#���5��MR&�n��tъ:��U@2���t�@���M��HK3�xNᦖ\�?�5hø�~iӣOЎ���l��J���X���yC�f��/��
�s�I.���g+1��9|HxX��Z�����4]t��-���Щ��-��D�65�2<�6-:7��6�vy�ڠ� %J�:�/�Agɟ�d�n�n7���1u��_I0+�f��ғPq��o�`�y4�Y�M�,d9֓�ڀ���~���X�D�j��ԑm8!�1G|m*�;��mw���b�C��'��n��`k�+j4�1,�9���H�s�1��6��ܣ���W�B���ct#�9�͜KX��+l�{�hx���Н�I"$�ە~��uk®�����Mǝ[G��bw�ʻ0<�����!j�])�ȶQ(T�(d��[�aR�1�d������Z��~i67]>2�Z�Y�S'f��,=/ms�C>g����Y�񏼪L_�������/��+{"�����gy���!�a��U=-�$4��WxYH�'3| �-+5�� ���A�ә�*�g�����m�4���1��4��q
�U��AZ��g���f�^e�pS��u����ke�P�������5�JZ��=?� ��?� 	:໰xk���?��J+_v�Բ�ui^w,O(�5�������O$�����!��|1�Y[�iP��aPW�_����O��ٝ��ع�v��۹���i������,k��u�Y�y�Fx1�Yj-�N>CU��f8���w���+��m�
�C���J�N��3?q�Z��[����8�'홳.:�{����Eh]	�Hm:I�:���A�HZb$���r�