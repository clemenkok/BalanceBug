��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�!��
��%Y l�׾����|R�bD�E���y"��O3�xs�XX�~��ς^���o���M�+Ϡ�����,�:"�-p�^��#��m���1�i�h�ӏ���Ó��M.�K��B,�W�x-7���[S��v/ 
�;(BX�Ec���*���ߠU���B yʇu��z}gE��iE�|
�� �a�a��g?����ȔJ�2\��-%�VS�r�܍�NG�`���OjÉxu�ʿVHL{µ�U+�L�чJ�?�9C=E��}�"����z�jy9�c����,�aj�D�����sK����a2�!`��zc��ByS{+��{� ������2���ўXޥ��x�r�,&��t�����m�he�<%
�����?s�?�W����BڰJ�K����-�����2ù�Af�N�H���01����ɇ�}h�	q��1z���7�j�=����V=����Eҳ22E�&�[fM��eZ��j���}G~!���(��t:$�15�fo�0�w�F�YT'�	 �UGUC��2�1RxFo��sL�"�� ��h=Q�N~��V9[r��"��*{��6��#��}�1�
��5*�kh��d�Jj.�7�!�]#R�1�����hqs�Z6��>�Ј~��
$р�ZGX�w�]��?��Q��r+�RI�g��(S���	�[�0����_�s�nr��B"��X��6N����zY�&U�V��m��sy2F9�m(.3�n�����t�=��*j�4��X)�ofAGM��/��8�i<U}�3�Oa+f����0�ڦ9묉bA�۵�ŝ�|p��+�:B`3Vom*=�
���s���p ��G��!H�X�،�;��߃.���N���H.	z}�^�:����[S�zƺ��������a,3�+�ź�ޤ"��ƪ5��6���bA{��i.�5烝��-���Ǌ�J�LFU��gd����R��p�`�OWtv�*� �fսQ�;P�I�A��UC?{�|�P���=��/�:�m���3�c�aԲ���X�����������I�A���Q���+��_!'9��Ը� �N��.�w�_���z�O+��K�M3��'��/CJ���'iv�h��yӿ8b��`m�b��E��v@ ���I�X�	�_,&������/�e׫�W�|\L��d.�,��ʅ��������F�#���I9�f��T����m���E$6!���R $9����E���@��!h4���'a$����q�0��r]j>�9�q�Eq�ӥ"f��f���+O��lz���8m̑z<j�]��78�Z�=At}-�wip0��B��L.=���^�Ö�Q�M�P�_G<�hBA���M��B��_VB4m_��(ؤ� :�ª���5r2ݎ����@���g���{�������!'�"L�=�FY�?PA@��qCPX��>2U7Nx��XA%À��ަ�,6����?I���'������Ɩ���1����Z��c���J���^Ĺ�u&�����A�,���˓�c�N���SrU�S�
wL�=
����_�1��g�.j��&�֑���8���V�:�+^	�j\[�dvu���|��!���~�s�mj@�SHeʓ��"���z�2�3i�Tp��(�O��Ot��u*��P� |�q�L,��~)m�F з�s�	-� �4�p���j�	n� Afg{w����I[�?ɧ��o���Bp�G�����#���z���V9�(�UC�k�J�h�P^h�5�]�����k.�mž�o�wh*x�kF��%ڈYfD��]�č�f*q�0P��My�}C�����6��65@�U=�"��f e�V5��j����� =��:�����
��V�1���n�#9,���|(�n+O��܏�Ľ�XY�)"%����,w�G_�*���\DZ �$K�u�������t�����!���"!�\��%� i�����TX�GF8j�vr����=9��d!�ֈ���c�Bg5#��,����c��	��z��JN�Vk�5To���Fe��
���z��:�>�$�a���k�u�ӴO��آ|
Q��뉚�W�k�Fl`���<��iAG�	͏��o%)!�D�)�S�g�H�E~� #Og��-��=r�?x����Q �$aH�5/�4�gcw�'�>�AW�~��U[�:|����kr��T:�m����NrRM�8��UB�9�4���.�F����8�LvUˀ�8ü̫�)ͣ7LO�jg �Tz�]�jR)�14����V�c x��j&�א�ia�O��Ĥ�a��$�J�,�L٣��}�%/v�4�n�ю:͡֎���p���M2b�j�qcAI�;S��R�ڽ[��K�E����"�����\kj��#*��%O7�%{��j��_\�1$P��:עP�Aqz٧������Z�?��������؆����\��E����?i�4vg��&+��Μ7���e�n�lE�]W]�"@��+�T��j�C����#�:�24�;4�8�9OKw��`A*��oԗc�e�E�'��g�2��E��/��]�u����~�I	#��}=����YO5B� �X>(��"5��
6��a�����c¿̳?�ޏ4U���]g�S�@�~��؏�yA��5'b|�5(�����6��OR�+�I'�^�S�Y�\�&i�1��L+�r"CW�gw�ΏÊHRJ�s�����?p��!(��P��J�H�\�S��� Ԫ� *���R��N1�k��'{����K�t����WA�&ש�*&V���@��B\���q�Q溏Q#6(Bฯ�5��ի���]���^ ى��\�Ok�N��L�5�*4�<.y& ���+f�ض���7�>�}j�ʱ��"[�$�7��I���z�+��u��D"G	0��&ԝu��c��ҧ_�ED~l�ۚ,~Z��ҥ���/m�/W�
j��,�Q���M}�����ťܶ&��k'�e�vn�ڻsi{JLv;i�
���sΐ�Q��j,�L�Ea>NXW��в��v&�)��p�.���w��Hۂ�`n��{ ������[���cP"3:ɑ�7a�l"\U�{&}/�e�i��O �\`�~�u�ؒE�*�B]#L�	��~Z��J������4h���=�ϳ5��z3����KM�ZF�]���{�]"���U�~%�XI#��eL��.�ԇr��I;u#R!�1����9㨛�f� Lۍܛ�B�����G�Ns2pm��䎞����o�x�M���� �ihV�)�c� ����胹��A⦂Z�Nά����J���s6�9a��1r��!r��L}���_����d�˄��SJ�I3��,��2�]�\H���O=�vo��+�3����S��p������j�i�v�h�1ݛ�,�9���v�t/w������ɭ�9y^�~��~�J<{�D�`ǩ�wJ&������9��_ �}��LU_���qU��#�������7�T�x�:8,�ٌ�J_�0�c�E>e�즂ߎ�>g��ø��+7�bP/m�~�Y�S�+v'[v�F$Fo���XE��g��Q'�3uŶ�|s�]w4*��"�Pa0ԣ