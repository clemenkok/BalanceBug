��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�!��
��%Y l�׾�kqDL���K��1�`� q'Ni$7�rbV��N�l��ǚڊe�����/�V�(F^c"�w��㥻�4���#"�ʷ���=Ypl\s4��>�1Fx\$���l�m^����~��,�yg]Lw�%���)ě)xU�	��0��N��u+�3�vu�aJ���S^8��\ʵ8�a��>�ƪ��%W\+˷کzH}Y�pK��y�%�.3e]��R�@��y6X��Jm���3�Tr�./���6�'9A#��s�rH#�M)2`�[����ޟj ��OT��R�M�%����������F���>o�%xK�,��T��Cݏb���k�^��[g�:�k�ATCf&�ML�J��	m�oZ�l?3�x>=�&a������>�M���ASt65�$9�%҄�� 
i�J�g��l�/|�	�&p�)���'T*��¸�W���la����e�Z�Z�*��c�,����[Vg9l~0���f�z-S$L�Pob����{s�,ݞԪ�uKr(��4�:=���$D��x��9�JƆs���2����m�#���o���Vˎ�Y��&�v��X������F h�/�!��Ь6�|��a8����*Z"�զ���8�����~b��	U7�u�:*��&����㞵];j�P�Xg0�}�Z�hlr2;؅�)��M;\�'�5�d4��Tb�Q�HG��6e*Kb����Ҝ��7N����C����5�Qi���*�(�zM2Mh#P�2 y#�(��%�gv<��T]�M�r����_+��ܗmx�f��ay\s���N��WcZ�7'�q
C���UΡ����p����MW��3 me�,�a8��HPn�|��k��������`G��N~	�3����v�������},���A�.T��k�Q�
�G���Z�j�t�44pK�����zX\tAK�,��E�-���Z�	�
�����}mnY�
��l@$�*C�V2{X�g�k���}��|��R�%Cfn��j��q�\�'4�Mi�yɴD`:��ަ!]�����CǨdgJ;}�|h��z��(�}>�#����c�DlU(H��W=JI�����g������#!uO�vJ����F�m=���P�����W�;$���}�b�>e�-X�4��K���ɨծ���:Pv��E?��'��jʃg�~7�,�=������G��mG�;Rb/�c0�6��؅�,�ݫ��%�;G~%���ʢG�]�A���Z�v�A-?�?����|����u�b\u�Y�T"�K}�B�YA��N$T�T��=*���ծ�S1�`I#��֐uzhq��*�����`̓DK���K�nX݌o~g�`Λ���nQ�_#a����]�м�;�*�UtJ�@��(��	�5�kc'6Fvvu�S&�osV�M\s�˓CAq���g&�x�Ot�ד���[��g��8,�����QZZ��
Q��E��!���ʫ�=J�o޿��W�xZ��r�E(���{�:|6	�0�-}j,[��Fџ5c�������vF��I7zŎ�u&�����̸mbc���.GE0���0>����N���m}J���X��)U���Ό�I#�K���c���Op�XT��{8�@*m�a'q ��hپFp�L����Ր0]mq5���dm�l��JP��B�>�y]Ae���Q��u��"��g�+.��QK2��#��(����!s�w� �Y��8?pi����6��/��.;F��чx*����ր븆J����ǎn
�%\X	Xҋ��#B1�TXB����X�/�Ֆ��w�{P��������W9@p.wv�{17[���sE�_Ǝ��~IG�O�RQ���M�����I����kL�������\�g���m�]��Q��Y�ǖ�-��^З/�ض�eh]Œ���U0
'��o��_�B��e���۬gx�KZ �AP%��}S��o�O	8<�>؎���7��9�pۭr�Er��w��*�qk���
,a�/hKY)��Uk\[��Օ
O�D��W�Y�����-��.��P�"z�}β-!�����_��6"�R�������Pk�&�J��]��4<B� ]_��+P�μ�r�(ᒊ���V�b��~B\C�'y:�}�Ĩ)V־F:��i�mڋ�Dq�:�PGq�Z�UOQ.�w3A�f_{�W�S��N����}��t ���yhaWم�CnM��%�,a��ej5Vt�fİx��~IeR��Uv��
s��7U���7]����lW���%����;�yG�|}�� il�2m��ac�MA<�H��5��??Q.C�^���e���t������c_4 Z!�8iQd�8@B+�!��37%��HP�5�n�Nعj{o](�]t�a$���]/-���%QOe%z�`�z�wAb[4��Ǖ	E��ܲ��6��a1�A�e�\X�c�K>��z �8s�U��p��ރ���k_G
C�qE���@I��gڅ�k�8ziӃSL�OGQ�yD܆`�h7�Լ#^��Q��
�<�X��.s҆��?�ķ�@,Y�����TiWy����8����r����h�u��6��1�R��NLE��.ODՙ��`z5�a��K!!/���,�4H&��U_Jׅ�t��y=�<'��C��c��8�L�c�P��*�%��C����)�4���I�4��o5g�ˈ�r�7�����z�4����%$�A
�m4�W�1����w��2;&#Wr�R��1o����b�t4G��M ��=�(}Q���	�����H���^3{&����[�3���v�����,�+�E9�v6Wao�����\�eӝ�q����#�CWOBrv�<=����s�/P���N�6S��i�����{Pt(;��ըD(q-����br;WM���`���;b��<��7���O��@d#h�R	�3� +���׬����7*c��jL̆��'xޣa�珡Fq$������x�[wi�P��H��δի:0x��#�M���}G!����p&<{�O'V�ɞؕ��G�n�#�=p�=����<�q�_��I�%���Y��ѡ U��M����
g~͊^|�?+4�?d3�oo�� �1:LV�>r�ڑ`����G��e��gE��V>�A�����4��S�H2Y)�6�����S���<- ����;(C�$������ڣ�k9��1��X� O�b�bg���΍���D��4\*�e�6=w����mltK�jJ�1����vC�E^՛ǀ�s�9��\Gcl�^#su�p�wSƚ�|��V[k����Ӡ^`J����;8(�#-8Ϯia���"!@��آB�B֒����LA�S�MPѰ[�2XSW��.��υ'=v�,�SJ��C�ѿ��[�څ��^�yx�T����i�܊t}�U��-��B'Y�kK�9���0]Ot+�:��2��A�<�
��#s���������ޓ��$�T��G$�~H��5�)�(�o}�ˊ�S��v�A٭Ŷ�
����=,٧��V0US����S,�Z����fl:DႽV�25\�z�ׁ��Z�r-����P�!CPL���
����{�aS$]EQ���sk%�r�R���/�G6e�!0�ݥ��=&�o�;�o�0,=#$�]�|����m���xS�_zY�2�R:Z���*�M���il �ή�Ó�� ߄d���M~��OP���]�c����vC��������{�0��x����(Q;��ͭ�<p���߷r�� ��q���g�%!7�S�/g��H�e�!<M*�_����8�3V샛z�D��$�L���F�b!W}И�����*��z��K�Vm����^�oj�u��ǁD� Re�P�"�i�-�i��
��9�����|��S*3R/��g)z����rG��g�S�"	�B{�B[z$ge!@c\$yk�7�j\�n��=�{F�)�o}~�I3�
��G�(*�ZoK��?^/��
@��4�׺��G҉�ùO��z��t���P� �"��E��z�W������ˤ��eMP��A]�AqN��>���#����6>�>h:h�;5C�[��~ iͩ�:u�0X8<��U2�Δ�'�C2b�[�}���d� D��=��)���
h෬VX��D��4[��=M2q4H�*�\���s20�H����������CwG��q��|X���7�2�C�8�j�G��
�6�h�	C%PP�9F��ݠ$)�</
t�H��b@�C�u���eJ������o��NI� K��&u�}�Ɨ4�k��u�x>>��_yӕQ���ٲJL"kW��p����r8�د�*]�9EN���� 9�7��I�aod�lT̞�#�FB&4s�}�����Ϙ.Ku�U#cM�.8;3�nV�"e���t�`�E/l�U!�i��W�Jfr�/��"T/�%��]'K��h�T��wh�<2y߁}�&fو��^��`<���j�F��C	����_�Ï�jU�-ѯ_��XD~��V�ŽS�2Y�c�[�ܗ�2�ݬT�#���f�0�F%�i�r���HGc	�=y.6����5�?N�۾�Wd���8b��[��;\�C��_#�2�?��k�����Ŷ,Yݕv ��N��,#��F���$�e!���ܴ�6����7u�C.*���1~����տP�j��Y�1�]��O�_(h� l~˽+�$�Tq�'�R�`���@��{�",[KO��w!�e��7׍��6���A�P�?��M��,��v��kW��jk��`	-C`}�	-.sq��f&$�
�l0y��;0�fʬP���Oz2s����E�N=�����D���EPC>��p�@O�~A�u��p����kq��è�
w��/Җ�5.�{RQ��U#�k�u�)�BMp���/M׌d�5ޒ$�-Y����� _�� ���;6�E��'-�� �r��o$GǕ�1�F�{C�j(�f�:�y�7v|�q�/�bG�O.6��$Z'��g�UN���L�Y�]�#,a�i�LU���|9���ph�%\�^�܄����v���*;e��E�h5��ʼx���P�#�_Kl�z�H��}1dT��
�X4��,�eֽ����Y4B��'��������Wos��6Z&�EP�l�����}8/�|l�+��d�������.%�
���i9���h�.>S`W�R�%8�{�.�o�Rj��c�������x���lmT��sG�5���э*FL�B#�8,�K����S� ��	Dc%o�V�N1��;џ�z�Y0�y�\Iʅ��7ܴ�+�����5Ο>�N@��?/�%+�wbSAr&��-FN QXi�O�dj�o������!�@sY��p5�S�l���`s�MyM�o�{�Y�0���)�oU[��� {��C�\w���s��d>\2½7�&?��1t������P���_�de���߁�&����t���IuB,�Z��/�}X(�E��j�?�Zc����i�- m���m~�8��p��2��8eC�`��d��wR$m�oڠ��a(&��]zޣ�#�E�<$�sѱT�.n���v$�om%��03@�[h(����o����������GM�y���p��������֒��e��2>eS�/�=H?�4���N0$����_���"k��n?+`�ݭ�9tJN�TS��K�i#}1��R�h�7�-h�-���1��JεAR�mc���8�
�@��*��}BQU�A�(�>��7�Z�|�E�/��v�4Y������c�W���s��J�N���O��W^�<8�	�$�6m.� ��)�uw����^}���=)��V��F�;��x�E9��[��e�U~��|�Eߌ/0���bY�`��[쌘)T��a���o?�%֎z� ��W���~3�bJ8ʨB�t�%����x<�t���ơ�9q�ˎ���K]����	�_@X�eO� ���a����lPT��$[��.&	K�˨��QY�O����y��È�<�Ol�o��O��d���(�8U�a:�`E�f=�س�I~�$	K�}�<IY�UZ5�W��I������Љ d�wA�q�Q�����1Ғ��v��ccqL8�2�_�(n��Y���Aׇ���oO;�����'�摫������q��X~
�	��.��,����O̾��T�h�#y tj+�\��y"�grr�Ѡw}ۃ���s�@v$��2�)��8��-j'>�A���ר�.�Ui���B�ã��C@)�y�w�N��ڄ�O)�
?b���+�����	�$��~�d��I�&��:s}��tyK�gj
�E���q��,���ܛ�-�� ��b�F��O�֩�4��*'�R�T�G�fovh�/=���;W� �6�3K�K�a)�� MS��[>�C�?Gg2SS{����B �y#��H˼�8Ǩ�1�M�.%N��8��r�*�{��z��v�^�o�b��~^}YpZ|�o<g�ӝ<��9��(����M�\!z�)y���Q?j�r�t����.N�"\�ژY�+���cc8�$+e��OȊ�%j�Un`p��i��4ʔ,�1 � Ql������h]���ߧ�(���L��'���II��q���d6�bi�gZ��Q��2Ⱥ�c7�?!��4���C��g �yNX������\>��������9*`I��y��T�t8L|}!�l��4.�B���<-ð��ĭ�o�6֊��E��r�[6��K��}hr�y�:�r*�F�휀����@>P���
]�՟͎���dN�E`Խ�}tSP��,N��b��R�q����JǾp3z����76�8-�^��ާ��|D�����rr-�p�f	z�\/�Ot�ք����+��<2��
����J����s%�Y�,��N��/�);�81�q�B����L�I��2ژ�&�錝އ��'�@�C�����C�tc����=.6����t����h��m}�Z���+j��T��x��� ����y\����+@h�;���kP���@���K�q�sET�����g�e�r��ߛ�6�2�1�&pi[\��l� .���"#Y�oHjM�W���LS���I��Ym9 ��`rHx���-C;j&6��	���b~�0���x�Vbx`eؗr"T�HstL��7^X-�O1��,E��X}�A��^:�8}�x�X%E��M�qM��	}���^�����A�b{�`&�iU�[��"��!�<�YHM�c�r�/�I�n�%d�m[I��вgO�Ya���~g�MF� �i����OyU��Űf�El��t\9�S���n��_Uz>�a����=M$#�����D�/����`č�E�c�
R���S�v�@���ɁE���b�e��ς�v���Q+�N�K��T)/���`�n��ƪ�:�70�[ �-)^��僐V��E�E�����Z	��&(�,��f�U}�*�ڧf��k����(��D~��Xm}��P�p�?����s,5���=��鉭n�l\)�ƪ��͞��'0�k����eSk��l�O��	`?-����bX>"Iwĕ_a(1Y/=Ҵ[�g��_,ӊ����8��ܶ���o���b�:�|�v�@!��Z{V�	!PDJ�5��h����H(<�r:T���O2Y�Xw�2����̔�H�!E��y��郞�ߐ�1>qf\>�mx]G����E���%8���I`b�[���	�P,�6���pMJ���D(��4�F��a�)-"��Ī��3Յ���ǳ~����6*dX	��7�e�a�{���ޖ�RP��w�.����`�RM�*��A����Pی>s7u�[�t����C�E-h��xFc^M��uò�P�7Y8o�Ha��e��F:H�8z��������?.Z4�-���զ�2?.�U�at�o���<��ޖrFv�{�9�R���w���	�ɧ�V���[�F8��0s�?����B7LOKj����
{�����nO���������F=L��&�dxI�Gj���v�܋�����y�}��kžNΪ��La���},��kN�sG�ibi������x����]+��3�$�m�L�;+���i�#���SZ�0�h�m�U0��E9����6~��p{o�� �E�u�h:*9���넬��@�n�toǙ�3$6�[C����������%=-;62�~?.Sg��	y=���ָ���K���L�a��F��ߏ�F��
B��1�2 �Vj[�V�g�T���3��/Zx��C	p������RD$M�̊��E��/m�z�d�����֨�>|�P�wdݢ�������X0���^�:٩dåY#�t�آA�"?��H(�M�_%	��lj���xx�"�U�NLVG؛�D����)�Tp?��ӭ�o�B鯞(e)���e�k�?��_�~��/��}H?3ko��H������F\�0��:W�KPn�nh�0��ˠs�	lW(���wd��<,B�/>22~�<JH,Z�m�ETEƂp�R�f��y��o�e�b���!�!�U/� j��Q�h3_�x+����]D0���&u��NGm�c��TO�z�&������2�z2靃��������X�!�zY"s���|\��4$����g����-�GnA�C�j����8�90^��V�B�2�сE���╘@L��_�I�>9X�8E�Fv��p���)�����nj�7�����W��E�y�nu����ڔ��[���y����#C���u�A�_\��_L}��Y�*���[�3-�9{S>�������iJ��Aȼ��p9Ooi�Mx��U��VS��{�D�j��3}�Aj�='�{�9��j�������ʇ�>0Hb�hZВ/���%6"7C+�I�I�>�/�pF�����x��iZ�Gރ�����-��ͨ�$����I|B�xD��04�� �S^�ŉ,Z��Y��M��Ah3���ce@�����ۥA���T��&*rER�e�.&��]�p��ܰ��M�K�2ҝi�-`'�O��>(�r��`���_��O�;�P��q�(U�9CA�u%o(��}��>h�Ygv�����a�9�B�\�'��0��2�$� :ޘk;]QH��_�%"OA��3����pD�;D�=�͞b���qj�˕j��o��#��~ѣ�P57��Al�#�a�=ժ%���UQb���! d�0�(b*�����Μ�D�\��%�3M�P,�z�S\�4!6qWMvu���7�s�<���������l��G�(�_P_EZ��-��(RVπ�؍����T.��.k3�\�@NHZ,X���;Q���kAv�h/*X/��xK�z$f���\q7��c�瀁��?���%t�C�V���L�yT$����YS����2�=T��l��~���ADT;����(y�CsA�³��w�/U7�58�4@�`�%������K��/Ab��	����7�h� &4�ȉ#�&5r��%i��Mx���\��^,R�0��d==�Ξ@sb�vɐ�J_�9��	����f�l�/�����o�rJE�d�Y�3h���" $/��@��RG81���p-���3+�ߦ~��r�=�?ϑp�x7�2k�SXn��G�<��/���^�/�lM��
�$�(X@s�q���W}[�/6��x������b�<ڇ�ؾ:��׹�
��I ��XF�&��$V:�?�	��W f�lH��+B��251�
�^��2�9�d��}H��}EJ#�nK�t�n@8%Wj��T ��B�-����Q7G�.�-L�C� �5��&�����H𒝎xee6�PMk�4�r �pC��^V���6�Ve' )�m�\�N��|w����;`�&d����z��%���f*�t�f ��+ĥ
!s�~\�w��멄���!�9z�[���B� �1eO���X�r���p��m�#(��[[�V�:O�f.�U
��FQx�r'�_��dfFM��F)�<��t^^B��-{�nhj�`}��_,��9�!wIg�u�w�䢜*��	AO6y9}��t����7�g�F�A��h�o�x!f���:��F!E�?g�e�'Zt4�g�Pӥ�^}��C�\����N��e��g���5g����*�w���Z��n�{�*����$��!�L�
��� ��_�ޏ�op�;��@�?6ƝQ�����Q�g��ࢾ��e�6�:�S�*�ش�k,�MR���82^\�w6����T%�AG��314mBl��U zM�b�m�O>I�e�qD?4�#�(�<z\F]v��do�H[|3�5>��?��5���.=DJ"�3���#yp�´[�77�'�aIՉ� ����8ʥ5����[T�G/N��?ғ�Y`��u =Aw��KLҠ�1�� �ǲ���qa�eJ&�ppw���p���8�y�(�&<$�(��#����Pg��*rE�８�^�	��U%zuFL�si�c��9V��0�e��Κs砵�%[M56�
���y�U�0:�i�^���0�KU��S�{NnD�މ9�Bwhoqb�s) #�|׀�t��^v��L'aۑ0�A�:����YK�t��{qPL�s(�&����u�/Pl������z]�Q�C��@�$��2�����_�B3Y�nО��ć��K]���O���DNɷ����̺�k�;�U?W1HL�ڄ�����`��Į�Λ`�}����=��r�B ���Nf��F�QRd�u�X���;�B�v���7������1%-��!�Wv����aW.��l֊~�k_��[^$�"6�+	��aZ͕s����ʥ�A����K7�y"�?*�q����ƣ'oZ)ߦ�T�hا����<=���5��;���2��{̾���{��X'5� ��r���K��$K}z���@8`Dv���~}R!�J@���2h�Ȗ�Xd{������9qU˒H��F_�&�#t`~m��4Y֊��j�]�_���z,u�o�b��f˰��C5��x$M�6�>�e�uhcG`���������W�G�zЅ������w����}���بT�L�nz����"���Q/���/�I�Ѭf�jR�7����G^�D؂�q�d�m_Q�c�g>���w��^���hw� � q�\�_@���-���<r0YFd���u���TV��9�&���iM�}���_XTJT����t�8��^��7�K�q�)!?��zڨ�Fj������ra�ղ���h��nh$Pu�C�92�:I�3>׫P2���)��j��!�^?�d<���1w���"`�Rk��������B��]  4 ��-��3�u(�nC��e�-qO�7๴z/u*�7<����L�X���g��O@*o��槃p�q	'�����1՟ҟ�4ˡF��Tg$��#�}�t�ȕFG(��d�k�rn
\j��[��yS_�
ɰ5�ߖ(�HC,�9h%F�Q.���1J4��t R��&��LU���車�kjz���:sWۋ�$��
�������|A7�������E�}���?�m&��t����sv�\$���d�t����G�`���.N��Cߏ�P��rNA~pb���)������	a�6����ɰ�@���n��A ��a��S$��R��:�qX���^/�j� ���Kz\(G�c�!���t�ɐ� �ăm���s�"��]�	]�glP�<�A,1��
���.q�_�����sN.���r��]�ͱ�*�ё����l��{Z1�x:�nx$1��|}�f�zW(6I�"����O�أZ��8����l��21�$�:�3�^�$I~��.e$��{�}5��������Yn�Xj�^���t��j��+|�kڑl�|})��}�:��^I�A�ǾL����Gh{3��FzN�Â�GŊ�QE*���5�V���x+[�Y�D�?���2\-�m�Ď�1�}.�� V ��7깻�7#@�m����kJ>~Mk��O�V����A�	��h<��\�܃L.j��!`ѿ������f�������(���;�VW8">!��nZ-_n!�D�W��pW���C�~a�
�P��ɶ�
��	�&����U���'���p��@�֮� �`��'�uO�����j��|I�|��J0d-j�ʮK��6��}ޡ"�=�>���_@��':�r&s�ՋY��K+�q���p��4���/˰�B��9�or*pB�t�g銤���5zֲƛGL��s��u���e�-C�t�O��1CϠ�̛�^�,�̊w@ �f-���x�V˘�r����P��Ͻ��́�6q���;,½?c��:����o�l�RLvWC��
aG)���]N�P>�wi�k�����zS��L%}�Y�U��wY#%�ON_��zl�����D����=U��aD����Lp
���_�j[��S�?�����]"�/���׍�C[��Cٝ��۬@=��w�lO�vO~W~1}D�K���M�G��q�6<k���6����M��� ��OH�޹�iQ� ��b!�#�Gڟ*�l�3���nލیH;`F�*E<�P�B_)��G���W��K���"A����l!A�C|��*!R1ܘ��e�˜߿A���{�]�ʤؐ1;�`>r�ׄeJ��Q���v�Qr��6�;r$�~Q�$�wu��M#�A[�̃�t�v@��ceA�P�z�w�e�"��w��٣,\o�c(���@�l�d�t�x����ѵ�@/RJ(v���������@%�@;;C�P���!��'4�ZB���EꜴo����k��Q�d=�ol�98�����M*�(Qʍ�L�����G��x�`8��u[���-I0����J��_�l����qV��u��S�� �*�(,L2�;ֲ�Imة��V���'�ٰ`��צ�C��MN�?�i�����*�����C���{[���W�00��\��s���E}AK��J�&�V2eП�'��<�q���+T���s8���o�5/��Syf1�A9�������Q�K_��b�\���t�`]Rm�N�i�,�;���]�S�����FZ?�� �w��:Շ ݐ���>D��ư���l��~�|��� ������v満G��:��]p�֯p�.�g�)$�m�՘5ӝ �2Lx*\��Dۍu�ω9�ğ/��V�.6z{b�S����BV
�_�<~�5���v�n�i{���֗���z�.����ԵS��j�7Z0�������/7�Qn��H�Y�% =k�T��f_sTg#�Ԡ�;�������hF����	6����稓�SB�oyl U�U�_Ue��b����o'�}
��Ǝ=@S�HЪ�l����`�XEf��s�6X��=�s�J�����V~��������d��ֹV����!"(EG
���_�H!��2���+��0ZYk��Rqϕ�"͖9.�/40����V۷�rÈ9��B���
È�'R��҇��h�c�L辰DVY򇮚j:�7�;�x���B@3BM�f6~	q�0z8k�Ƕ �i��fQ,�fs:�9���d�Hd֕�<�@��NXBߝ{�#*��e�d�ʣ�3R�>�B�*;���e��	҃v3�ًt�P�ӑz���&�g��a����bxъ"ݝ�g �O�:���y�-�&��dɜY���ØEs�#�w��h��0ن���Pl4y�G����� 	s̎7Q����@Ղ�Su��%>��|���g0�w��j7��޿&��,���GdH�(�W��U?w 빘���v�����
h���"CvL�_�FO����~�q%l���š{s�,ӵ/�ܮ�s�i_ar`U�80��'Ƌ�L΄W[>=ih@�d��P���#��A��Ia�;o�4r����@�9\�����
�b�:٘�J��s웳���=�ߡj����۔�f�����W���ﱐ�(�R�3�����|�cAs�m��ں�BTa;��'���l��$.+�e;��:�\MʗT�>�%I��^��7����Z<��:�y�������G/�Qڸ��Υ��.[�p�f��B�\نl��g�e�V`0s�Yr��p�R��fk~Z5�ɵ8)oO:a ǂ���h&����ѓ20�:n��;�c(;i!h]�L"%.�%�	Оu�D�˲��5��Q��5u���#���K�#���d	e����2�;jr�j��a�b�u4�$AGR>ʖi�)���N�R��s��{��G�g"}#���_@Qg���Z�>g�O��j�6���U�j�2�;O%v�����@[�U�5����cݤ.c]����(Z{��^�"-��з6b`����	Z�;q�����\p�� ��%%2"��@���Qd��r1MR6芫5`�{˄;�qN��@tӞ.fF�)��*	�!���� ����:���N��UD+%��V�>��#�=�5��zǹ���</��?��s}���xV�F����o%2xK� �p�~Ⴡ~�W�(��5�HM�$�Xd*"~����/���2M��Mx;�2�-]RE�3���ˁ�+�zm`)CWM�F�GZ:U�`퍡�[[iս��Bړ��,�G�}��ި������?�#t�%)�"�i� $\=� {58"4������3w��6=�H��?=|��)���3�}��|�gO䧎cP���j�	!,�=�Sg���dI9�O��/a��Q"��~���(�#�X����w�-���G��9p�.�8���� �f췯��������$~���XJ�K��{.� �Z�޼���p�_�ȠC ���*����%Mx�@�k�Mx>�� ��O�+�~6��$�[�]#�N���.�-�)z����$�^�������w`k3խq�,|��j�L2hUύm��ǣ�*��p�6��1��Ṁ:n����Xx��&��*E/K���ޭ�IB0ay�։KZz�9��<)1��� d�����-�p(4u�d���@Rc����TgN<��0�q� �9P<4-�vW� �*�|Hک la�F5U{f�b�KG{��Q����g�±@�;�C���og���\)6T�>�w1�L�#V��u���̼I^���춘l7��OvBJ�(E@�m�60C	�V�
JKB~�׌<i=��`q�QHyp��4����ܨOyJN�p�
̉v:D��
�����d����lr�y	�*o KK$W`�y�h1۽z=%��$0��x\���J�}E|\T�@9�������6-��rl4�ԍy	6lˍi���}�G�v�ى��4�LaT��G�q�1���+g����U��'��ߎ\�����=,�3}(|����}g����#؂|ε޽�*6Nx�͒�I���t��ވ�q-)4�POl*%lB�2V���1|�b6��@7s����>��~�ؖ`���2��L�r��mL<��\�a�#	$�����Yן���5�B��d�ݴ8WL��w�{X��Tz��_�Qw8 �zY��=T� :�S�%¢w�>Ѵϵ9U}����)�5�b%�~��ɜf:�!p����`N�Sh����dv=��EC���7֜>g9|���Z�禤��zr[/����sJf�g��e��q���	@�J�!;��̃����0CLQ5��R�1�0�(�O�1g��h�7���|�к�/�ǚI���ki9��v���`.�y�76gJ���:	B�����b�sk@7
��Fb��Ϣ��J�l�d�ئ��]�;g ����Ϡ�o�@UL�Y��������R���{Ko�Ǟ����;��Rp�-&lH���Z��d�R�S��4��4IA�����		!ʳZ�i�����.F���u�o#�V8Ou�26L?�`�]+R�~x�}�ɃVvP�~Ӎ��A�?�����yG�Q2���(��e#�QPYx+�`��t_˫��@��ۍy�%N�Yli�q�ڑr���bx\C����u`x����s�:SV� =�n�wpH�/8��4	A��ؘ��~Lۺ[@���\jvij���r��a�,*�=��R�R/�R�0���c���QI�v���+��L��H��P8��Z���+��n�Kz�n֜y*��a6���+�Q�����H'�Z���K 7���Fe`#l�>��L����)�#�~�������񈞶��?~�ɳ����wAWjyk���s$X�&��N���ƪ~&�]l�)�R��{��H��U�Ǵ��!�Y������F2*�v��-��3�&N�ӄd{&�-O�e��ՍdTw^���0�%�Δ� �R�d���;t2�l��oW��9dʝ 4a<�x�ONX��sH�s7�R�x��^u���iC\u�g
�co�A���2������ �x�ϩg[|���@#4&��<��gZ�@!=��r� ���� W�4��R��펙�%5�bz����8��WX�*���ؔ��=���0��u:tSJD�o>G��*dc��;$�O�7��T�N��D*3�E��S���[?6ҋF&�s�>x
�������?��{˃��+p�=r�A���facv<
����W��b�� �F��|����$6r� ��P�#}_e�l0�o[J�Ϊc��I½3
st�~2pLM����#�L�*z��N�ɾZ�,����9�4JJs=�VhjG~�=G���o5��e�����9%5���M�v�һ!���h�i��xg�h�#(m��� ��}�i%������O���ɾ�qi]��#���F4�-:�F	�5��0����]��*�Շk�6��n�i��B_�۠��Ќ!��ya�	�0�\#1B�����W��������1
��9KL05�BT�,�.�9	���%=����zB�M5�t�fǄ<�H �A�0aq��ކ��}ˑ��.�>�1���l���BVdq�T�~bVQe땲�ß������ ��Os�Ap�>���|c�XmB� 
�a<21�c�D��#+���������X.v�
	4����5ۭ��J⺌*���T�$����W�B�A��f�7���{�݆��t�"�ge��Qt�Ęl��4V� ��9����M��!���H�yB@��7b~o����EU�7��,�g"���S�8���7�+� #݋�/���iad��A�(��x+<JY�
H��@a�����D|gnY�	��7��>y�5��j ͒�2���fT�A>�N��v�h�QY[��΁�K.y���Ngwd�΅�꒲�Ny�M|,Vķ|�b��܂Ǹ\�/2�v&]���A����>�4��HC7�$�F΀�+��%��(Nu(�>\��DRz�(�9����k2� ��i�0ZDP�D`c���[�U)O�KEN⁤�<��;ڷ�j�
���ekt� �k���K�[�l����W��.�1��u(0���~�g*���
40��B�(?5�~�D{�Z+]m�vC.`���^]�5�6�����k���K�Lw����}[.I��1w�Q�묊T�A)�a��U/�΄����1�X�sEE)��V �n�@;y�����+��%~/餴��w;�]��:J�7&8�{�+T�7H�=�N���-��� R�$�>Z��2.��N ���k:wB�����j�Ѫ`v�b����ř�
ȃ�4\��&'i1ih�d���_��t[��װ�̒b��h�b��Dw
-�+Hw���2<�ߠS}��I3[�zX�HIp�k�������|峭�=$�sl��kt���u
����3���N�`�S7c�X��V�.��zKr�x�+RQ3���j�����Vq���Z���2˜���!��{I��%k���5� �T�mً��[��*I��黒B����'Ž4�A#7�*Ze)���y|,Uak���_������dWR��rA��3qma�����%�a`7+D9�n� 1�G:�3�t
�x�(f{���6��1#iL�N��p�7}�a��i�>>;�b&h#��a�ɓ,�G����i�����������"��4�E�*�؍w-�W�S\2aQ�}s� �s��6p��4~�o|ۜ���BHޮ5�n�4����/'���,�J���h�m9�vQ|u lkxE#���Jr���qֈ
�W�@ ��@&�Ћi���dT���Če����v�>Fo�J鷃�ߜp2�%�eg�f�"uS[�b���D�yIɵ'��fZ��Jhp��X�?EG���׷�k%/I��4S�!_<J_n�`���'=�y1a2�A��'i�.�^S��`{20����+��5�}p��r�F�yy#$�7$���GN�[܊��R����%���|�#��.���K��S�<'f�]�� i\�����1D�(��_U��UDg-�Ob�����E�Jx=�ٷ�>�*�A��D#��"�6�ѳ{ud�k�
��oi��s�c�z$9�|��5#u|V,�/��s�E�\���M�o�.�<f��|����/˞t/Ufq�[�� �#8m�t�������ݍ-ǒz�BĲ*��M,�.=G ��9���%af��a��Zh\ցo�L2*�K��������0&/0�ɵ���}t��Vu�������p�������"#o
߭W�|��b؅�zy\E� |G[����Y�$i���<�Ws�r�LT��YqN�*k�:�X�i�S�p"�_1bb�,�!�DNx��Ef۴l�{��i�޳fu�����β�J��Vq����Z�^�������T^^�'�.�ʠ�`��K ^�+��`���F�K��C��fWkg�R��A�]�d3��6���=��$�CV�v7�w���U:��6ڞoڴ�?8>;+��R�ɾ�o�R�� bX
,�<[�	\�t�R�+��۸�����m���R�*�<�s
�z�	Ļ�5s|t6����Z���	(�-�J�[A�K-��p�U�ލp�6��$�I	F/�-�x.R�-v��^�����Z�h��g�͊Єj����ބ�k�Ou͓�7q�0��'�E͂"p���U�tx��>׉�m�i��,Y+q��8#]j��"� a:��OE �'���"|�YH�,,i$%m��߱X�l��D�r�����f��Q���"�W2�xp��SǠ�f+���Fq� �/.k��-Ce5���Q����Lv���E$�Q�w���'�ՠu������n�n��6q�E!��𱋂��pA��vi6���Ȯ7��������X�i�F��2{h��H'�QMn�m�@���ZcW���j�[u�V�D�?�w���q��)[��cz� �� ����间%77��L���UMPU�EH`���#{'��D�bH7���y�J�~	6!�?6��酴J��T�]��3�����R����)�ܞb�!�*q?��4॓X���h� ��d�B��(���{����y/69�a	�VN���2���=���p���obU�t�,���nK|�C�;���}~�u,�>�� dͰ�:������F����g�{W���5:�SIX]�ck��BN�d�,~q�0Q��5k�y�L#ם����9k�U��ӗ�}S���Mܫ����\��Ŵ��ij���Vx�n�8]���~�u;DlD4j02V2���NVqT	4���K����]1��F扖x\-â~j�5GI��@��vk�S����| �H&�q��� w	]<ѣ� �%��|��`J�Ŵ�4O��.�zH�%��2A�x*̭�"�hv�2Zڐf�O�SEc�<8�g~�_G���d-�P��b:,�c�����CۘV[D����ʽ����
�~W4�a�&*<n�C5�B{`ѳ&�.�W@�mT��`{{�J�Cȡ�#/k�ԅ^�7��T^n���/��PiI��ܽ�ćD��1x#���h��Ǹ�kzZT#�P�r��.>�C2��[��8f����y���H9?��v|r��4A�	�h�����@0��x
[�c���g�L���0�b5s�@��-N=;��ގ�>ȕ*�mUFJ��v{D`9����炭�`�����׬��zCh=�Y���'�UK�,����$D�xV��j��{/��[>� q�z�����ğ�Ъ/N���i�w��>���hO�!!R`��]n�.W�0�}&\���8��ߛ�oF�*}i�/��{Hͭ&k�Xq^��G6����
�l�L�W'ֱ��>�+T�Ȗ$��Y��]����
)A�=
Ə��*2M`8*�WVtB�, ��V��~1MV6�ƛ:��=E�5����4'��J����%�w?#�>�%�SI��2���J�BV��24�¨�?*U��%��d���,���rZ��"��`&�hI+P��JU*�u>��:�hg��ζM�������B�"�h�gL��'P[�AQ�v��o�!Q� "�64���\eN���>�Gz�;��2�.��ϔ<�,+�m(��r\g�E|�w�K�C��1�ec]	�$5�rv��L}0D�.�'�0���]v�k6#��Ј|���Mc��d�6�����I<v�w+�7MEj}|�����h�X]l��8���L}�A����@���T	%��CTؒ�R���t>Ƅ����z��n��Ds
���＃j��l{xX���n��r�H��L�iu�r��2��w| {���]z�7��n��>y6�"�z5���{�nu8�>AE���������/���.Вя�H����f��Ӗ��He��"�<	un"+�g�Ʌ�i��|T�<i\Bd=z�X���%`�Z�q�G=5S;hB�i/��@P nm�����R��}�\��I"b�Ikoi"o�9��j�O;�x�����q�;91��Y����o�������L88@}>�U��~u��!Ey0g�9% Z�!���#	1���<�>s�J�[���������p�y�#[af��9�ks�G"͚ꭔ�Gӳ["d�̑%�L_f�&�~���"�^1f�]��R�vI��\^#�,��ɋ�[>�)L�����i�!p������������P��X���A!w���(�U�e�>n4�z�����s�i�]����E�^��?!������!���:�O'\�rW�P�j�����䱹mzʐ��]JY=F�U��0������{����Jc_�r�D��6=��7�U�æ�h'kY#g�$�>�jo��a�PN�y���D��=�mT7�����`y���dN���ۗ0��ݪ��U%�׽]�)�
)��a�!N���<>1=f�����H`���G�)rb6�q�w{��I�]���:��,��-�V�َEt��	7�MBf,\��/����)[���'땋��i�����U{ګ�+�	�}�hw�����#��˩*�d:�x�e����%eTA�k~#�v��[�7�CZ_���~�HL�\A��.��N�y�/2ԣ�g`(��	`c�s�\��c���Q��9]��|0a�M#-�so�M'�o�D@Hbh�nd/��n�pr�ͼ�1f��{�h����L��dE�{�MAo��/�l���y6ⵛ��V�Cδ�"l�).�X��#���P��5wg5v�i��O���8҈Y��~L ��K��� x3��������6)2�8)�M[���� ?����H
��ZW�oKHP�v��t��j>�y=�i���S-c�Hj8al�nlF�J�>�m� "P�y��-e�њ��zD���S��:#��(�F�N�c~5�0����wp��Z��}�a����[c�z�}$M�NǬO���0_[�}��c��}qFl����i����Z����C*��+�(�S�=&\ii�32T�{P��7��]�&���:/CƖAb�*WSE��
��<t�s��r8Q�i0{�9�ضׇ��;�C���b�0x�k�wu��GF턟���.H!�~��߶�����+c���	r���)��"̣I]��R�\�6��( �H���˒Z8�" m����O!� w��.(�_l�˙��g�M�J�sMg`��7�:�Ȉ-����WȐ��A�3$���y�'������$\�u�}���D"pE���|�K�y EH�r��hQ�|�vC̂ZD�yrI��`-��9�}�'[�Rd��� �X4"�˂���d�[���;�v7���Jv ��x�Pr�0���Y!�R�����Xx�h=�N�gH��P�6T �譨+���e��)���;]2�J��4=$_���Jċ?��`�E�.N�ҽMU�(�f� گ�8pO�QNfa�`� D�A+������!�� !@��h�e'��d4v1�����I�� T9x�(�9]�!��X�5�ޚ��+�/�S�����|U���ıy����ռHL%���`6j��om�����k;��ض��Ê��f<�W\^8(�'0/�!Ϋ��Ai7\�B��v�]��&��s�RB�'r��d٤6��(cۗ{\w����)�&"���x0<�K %���`g��`��Z2��V{�F ~ÌcP$�:�t����H�1��Dڳ���w�|���7\
�{�f�:DY";�N~Ag��	�r���]�TЏ|�$��Ә�hlh
2�DD�A�zZeuь�\�2]�0iF^�1&���i����J�h�޲C <�9����m��(T����ݎX�x5�;�S#F,�$�M��{V��Pp^<�75�S�p�T�X��P@�܅Bʟ�3���)~(`j�vޔ&����8�k�uz�Z���d�5.U'��L�ֵ ���y%>+���yv(��_m0��P�r�7�(��C~��Ȕ�"�j&�?��p�ٟ��Sg��xUTW�/t��F+�?o�
�,���Qئx|%�0��7\n��h��ڂ4�*Q}�+�}!����˞�\2T<rS��WB��,kή@�KȮ��S9XN�G�\T����FѰ���¤ƥ�|"j][;l�����O)�!���8�
���P(����b�,(�ycF���ɵ�\x��;o|�k���oӄ=h�8�����#Iɵ�S���q8y�l���۲����W��e��t��	Jxy^&u=��ռ���a�7�R�рrh|<�T���)q3{$�acdm�h9w�ҝ;9��e�~�j���*Y����� ��s�;��-c����R���#v
���o-gpW�A�R�o������a����W2#C�c��W����9\/�z<���D�!]�v�@��x�%Bmt�"_}ZhM�	�Π�Y`|�S4�]��nm������8�g�����?!��A��Ȟ�~�m��ZFV�}U�#n/�n��C �cןpc�p�{�M��A�Q^�w<����IB���.u"Аt�s��"u��a�g��V	O��5١Z��ġ��z�!�zbX�5��C����7�Ib�V��E1��t�2P<�au���8��M�K��~��Q/?Lt�m��YO�V��V	  �9c���T{��1����_^��=(j�>I�8B���^������'�k���xO:�e���k@'ha�.�?��s���d!�a��w�s���܂�?��Ǆ����m�#�Do�h�iڧz	߄��(ޛ�Mov�0R���������o�^�(DfE{���GU�J,@��[� p�,a�_�ۨ�J�)��T�H&����tQ�گ�g�|d��~�� ~�]�&[�V��J��t7��3j�:�T�BV����X�YXQ���C,���������VM��bG]�~�^�?���`���҂�3��]mX�4V��(�K���{��T��KO���soM�G�ĈZ���
D��B� ��������C����>�',��B.=ߒGvfb��8Ưd7�)�ǋ�:�Gw���K�cы�p1q�Z���|FY7�q�w��b�$O�gq���3?��y���� ���l2���gn�T����
]��o��ϸ�>��K�H!a�__�P���)��������Wۚ����U�K~�nU������ѕ�N)F�u�h�vh 1���y��n�7Q�^�J���ԔLm������D49G��~����ߚD����z�a	�p�n�·�F�X	��+8:FM�)ZhY+e��W����\�Kis��>vN_{����xb�{��"x��*Q"�P�-G�4�t�� d'��E�I��@��6" ��]�GՖ
_cW��G$�qw���!+�鹽!?��4TV�Kо9{�!*[_R��=��7Fв�;^��>d�T�8yW�6�9/v�p`n/�Q�ՍZ�4�����Jh.�~����CՇ���>w\`εi�����
G�j���&��_vp.��]���@�x���A��A�y/����e�_�>�q�r:�y���4_��rJ���6���@�|Xcc���X�N�]���?���	<P�+h@��'�5t�un|��X��1�fkq!�!�Y���)$t���V� �*O0���FP\6{\f��jr9���娷��/ƀ��m�#��6I��03F��L�k�F�',�٭sl�L:T�D"|�jo���c*靏��+ؓV�jdх�xQ!�On6�6��)�w�^K
T��A�h ni���� �#%��,������>���A���=�-��#kv���y&�ڦ�/w�T�K=fi�ɗ[Sc�����5���f���/��`���֪�E��Ƭ�'@G���U�c��Y���ͪH�=�N�G��E=��!V�4�o@N���bK�����xV��z۾,ጽ3�'Iƣ�@k��P,,��U_��`HZ�c��n�[���V&��;b�k���U�+Y��[�J�G-�O���G�l�3�H��4�aovH��(����o��k�?���4�W�/�#~P�32?�Ɣ�3!��a'���:02^�*���6I���B�͝d�)��H�L����K�<z+du��m���H��COU���ෑ
��s�H�k�)��n�;�~��%n�iTJ0���$=�4�y�M�z/X�������#��u�[\���n�J��n�k��=���o����Mlx��=�ӄ!��o��Cg�/*��7��9�"������00�O{���x! @�Iݨ��bz%��K!ת����ԎV
s�Ɵ�H�t-�갏}��ע��㚬4�j��B�Y�9~�=d���c� ���օ����|#�������I�'"��C��*
1JW� �l�D籈d��^*��([�C�vrL�V��A���}�q��e�Cqm����U�?�ר��C1]�� <��L�FW%A�^~��&��G����_W�}�;\~�8��A��J����x~��y�<�$�����D��u�G�dÁ^
&���f!��{��	S	�sP�g����X�ج�-�h�z���ߺ�r^	�O��sX�B��u#�қ>��ڐ���n��;(���������.7�N���E�����&� /�<_�^��G��8^�g$��=�B=3�}�b����BaF04B�Ύ�9R1��y�3˒"�����<��
�s"�q5�=-�efl�u��ɟ �#|�1��BT(��+�-�ˎ	@s⃼mgB^�׌԰��h�{?��J��)��)&���9���S�-p��y0�b��}:6u�e⣈W���xo4���4h�� ��Op����?S�ʢ��NE�t�Rn1��؍�m���1(�m���=HZ��!�����P�_��h-$4l�no���Z��{e��, H�&�8g��>���o9O��ب6x�"�̮����h���#��U��0�5��ٜ�6������/*Vw^�C:t�z+W����T_��Iy����+���2k��ð]!M��ͧCU�u@L��K���ӌ).�����G/�YVNq�R����!��የj�k��M?�yL PU�w �J�[��$h$�x���	d��Ε�Y�n�`\��)ѬBe�)�'I�Y��y�ـ�ii��j�����$9.
f�Wu|��,#OP����ϛ�B����9�Y����NsE�J��IQS�c8�͝��9ۺ�ǔ.����6��e-��Ǽ���of�����w��ڹp(Cf��"� ��]��%������P=_[d��*����*H
�B��x�ڰ5H�_��{ �5�g�5)��Mkόw��q�����و�Q����Q�O��LztM��#��c�.�iY6���@�k�&��2F�Z;@�M?hї��H�L�\��2|xl`p(��|֜���d\�h�jʔ�6���%./9�ln���̈́׀8m(s�2�r-1��=X�P�܅� Q��sm��c ��-�K�ɶ��yu�CZho �\�*~����O�ۊtp��+b�����m����"���p��\�%ԡ�;x!穾��zC�"?��.��A����!��!A�+�Ixh#=ϐq�������ִZ�w`$|�c��.<���a�*N�J�s-.��n�s�Sۖ{;�m�Q���\	��c���A�D���$AA`�o�ŋ
Q>x��"_��1q�L�2�͛��f��z�3f
UNl$�-�_��J��J]"�J��~�JJ�x)�ǵh��X�WG�,١ڙ����S�$Y*7�rnWe0��Q�m����zʥx��K<�����H�ܵw�����0-RR�q��dw"`[�$_Ҏ�~�~�okDkN���� �o�[�<�gV���\TE�Ҋ�����̱��#���CaT=H?�υX��B"A�Yw�L�Q��)�	���
��]����価}�g`������\���_.�Y�Q;t�X�fq�Y�z���v�(,���mT!\e=K�Qcef9�%m�R�@?�O/�O�\���(9sP�9�Ӽ��ʑ�2L��.��|�}�2'ƸOva$nԏ<M�ҷ)�^������l��0J����R�_j��Ab�ڼ�.QD�;�	�+��A����q�vy��+�W<�PT+Q�Ι�����I>��;����h�8lQb�p��Ѧ��+3�s����V�C���'qD�j-*�_z%���!�x�R�>�S�q������>O��z/���o�0����Ug]�3���5�j��$ ��zK8�GeI1��k��_���B�HG!K S@I��o��X��<�d���Sl���<Z�#���pA�ϸ�yN�D�ġ�{��ۖw��;�{��P��K˕3�.2,��9��6��U�<�I�γ>��-O�Ŧ��nz�[3�@3�e���82������4���࣒n��	~"� j%�}�U�dE\�/"1ǇL #/b>�o���SgJ;%I|��0�g�,�~lR�I�%J9B(��y��1�șVw��[5��Tʱo��%R���t�ĐH[�P�*/6�D�&Vq"4#�bG�/�P'}������Vz�c� ���, ����sr*<����7R�68N�*>ǋ�F���X���r�4���yXQ�{�s�;e�v��K���D.b�Oo6�s�B�O��I*z9��\��p�~4�4�3�[�����X- qS��Fv��*�v��@�{T�$G��ݔ�4���4����7w�G�YS��!R³�6�Wg~�ҩ>a��x�p4<w�I�f�� 8���������rq�`#��F���w>�f���.����>𐜌
�1Y��Z����5�����ܾK[3��O��G�g�%L�PQA�ۡ��=�*=�X��Y���$���|G~�ʗ�z�7��T�в�P��G�Wz��x�(t�=�e7�����l�g{]:\D��d�-Cp���
އ,���<ʒ<Ț����$$��կ�Cw�=j��lhG��I}�E0��U�[�a�\Dm ��o���<"ۿ�fY,	���0 Jю�掾I������@��������ݟ���/�k@��ε�CE���V�x�����xn0�O�U)gdD���T)��_�ϛ�V��E�ͽ����Z��:O�I<����e���*�����LY{Ж�#�O�R|�>H��aN��v3�����-||؁c�uy�,;�yIPu����el@/d�-�@��J����|Pi�β��~&k�>%�ˈ:ފ".c�B�Y5"�t�ī�3#�TS����g��8�dD����Ak�<�X�?�\�}���V��a�v���-��1��ʀ��R>O��d�����:zhMA��'� �4�,