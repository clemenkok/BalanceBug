��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�!��
��%Y l�׾����|R�bD�E���y"��C[�ϱ�5�O���h\�F@�l*8�H�E-j�|�&�@�D�G�q�3ZV-��Yڴ�a�Zn�N�E	��xSIkG�����3��M�~���MgNO���ҩ2�_5ëDH%��᠈̽'�;���4͐K��t��&ڢ�*]u��� s,���Sj�<9�\��#n��^�
���؊t�Ӆ��R#��L�i
�@6F����lu�xu����B�ŇՈ�u�=��~���&�
�s�l)<��{��u���0� ��{k��|ql����'~�R�}���qq ����F#�J�L{vT�6��$�{q4�@��ʬ	̓�,`RzL��4髓�b���-o��x�[���*vD�F��hj�)�w�G���R�؂%�E�?�C	������{��@<;'�Z���aߔ9��%�wDYa16ו��R��3p��SW�Y�-���R T~Z�S�� �5JT)o�Ƙ*6��S�&��V���ێ��^֕�+&���K��)G�֬��݂:��;ǲ|�P�w��(}/�iH��|JC���pe�]�+�nJ+���=����mu���'n�U���5V,f�8�
I\���\�!ٔ�]K�/�"�j,T��:��۱�$J?I��e��c��	���_F���G�[�<��:�a�q��{),MW&�o@��u���Y�	H�w/q[B-�ɥV�B�����μ�)�|`"���.�z&�U	/�Y��16m#����Mԝyi�H0��C��mN���l���ܟ�C�f���g^h�׭������7aX3�ym�����.�{�����v2�r�%�űm5o��9'
}�h������4_z�w�hw`u-�F�����d]���=����T&�RV`�����@CIrP��vY���IK�1<|�����_�,~2�H0<j��� Zӗ���_�DԢ���v��Tb,���
�AA�-�	��N1��68��e2\h��Naw�K�Hi�CP�X�~^��/�0����1g��iX�}��%������J�����'�%��_�	�?-��a5!+�a�2u""� ��'� 9L/��
:�H�{�U�����-կ�	��b&�G��l�8P�b'{�s�Ă�q���6跗�a��֚��֧n=�ұF�􏍭��u0�r�hRyG�3��D��ޥ0 �#�~1̫��ޒcD��$³�̬Z��XV�N�f��
����4�n�N �r��g�ia3!`j1.�58�\go=��oux�#?z�o���T=���ܻ"p�]�����,��hC�}��S����ӡM��w�xt���SWu���9� 9��'���J_ '?b�
aU��+�|���2�{x0A�������VӜ ,O��X,��.SPMnqB���Y���V2uu��?c�[�E�YW�h����9����'�C��sn����P�,�"ϝsܸ�_��6��Um�$�,�r�a�B�$$�Xࠬ�9�`�[�Y���^�1B��\w�X#L��Pq9"4 ��y��|�����ES7$�v�Ox��6`�ņ~������Ng�R�聉���Tzl@9ϰGı�Ssр��7[���Y&'�&P}�>�ӆc��$���~�bKe<PP�A<��lY����!���ñ�^���h��Îy�q1��9��j��m�|��m4X��Ok�\�nv����.�k�Z��ᰓ�Cޔ�z�J����zJ��;��Fale�{V�D�.\��Fx֟A�6��A�$�1+!φEw��RE�����+-�T��������#���X%/C�vm����L�kLW����Og�d�Sꩥ���:{� \@�ӯ��
��u�(6 ��ȉ%�k�����䵞������o�G\���M�:��PW@rft���.\���T_��(R��C��@'����w;Rc�}�^ч���!�@��/���ؒ>g�J�0 ox�i��>XV����	6"�s[�"ӗF���ϳ����G�_D���D_�˵��Vbu�!-;#�?.�J@�G'�&�^Y�
hֺ�1�� ���2�?�y���&���
��=��Ä.��4�WX�
�&�%���	z�����|�(�O&�J��Q�@�_��O��je���gN�{|1V23��5���DJ	�W�J&Fd�,Ua�#j?;���"����!fB��;�,�lJ� ��b����<'����w֮�������렑$i�j�![�E6�!(1�h�t4=���$��?nR��e��� y���}a�æm�I�p�-�3���XVhY<��3����&�5R�/E�[��r- ��}q�)��$��Z"��%�p�VJda��*�ً�=q�>����6Y�-��@� m�6����HnR�t�9O�Sx�K>�8�l���^�-����;`a������c҆�}Hȧ�wp7�'��� /���'�d~�\����ch��Qt�X���X:�	�;nlCl���OC#���dD��o�;�hFc�<l�;;�k9ҒoM����!������FJ��]c�Ar8�R"5Tv����@�N�����R����_�U	���P��j�H �
YJ��cGX���9Kz�T�?��������������e�| ���� ��˴�iǠx�Z�tt� ���7�`�W��KU m$馓����@d!���@�c�¯�0��v;���������9+xQ׶E�� �x�5������
+|����4a��(��]� h�t��~�Ӛ�6�����IU����/��fm��Q��p���]Ggwl^9��[���F�="G
��0v8���Ba�*sy� s�s���o-����5�Rȼ�$��~�e8�U��oA��$ϴ�9���O���|�gy:�<"�,��=�����Z���'hr�M)!�+�;��K�*Yom���=H��@���:�Ҁ�@�߿�{��#�Rp���n�>Vq�r(8�6V&9�f�	A�5a)F��a+~-��<�i"���{��70U�<���n���8�����f ,���@�g^F�:������@�$c��H)�@���RW~�3)I5O\�7kg^t�,%����l+d�g2��iG��+6{K��%]:�ɗ��m�E[�G2��@L )��M@���9+&�sv�A&$�'7Fs�P�2�����3s�o��١^��]��ف>�tg	���e��yq1�r��gW��	�I	yx�?+<�	�<�RIw����ȴO&�j�<^���
������]^~��NP�"�A���%�x���TL��� #�
n��=s;�y��e����uf'Qk�7��X;RK�ۿ?m�
���0;j� �Whu���$�R�N+_��Oz�\9\�MY� ��su޺�շ�1��w���XG��{��l�8M?��<5�_���	s�7���Dꭧ!�Q�
��\��8.��e��������	�n�{'���D� �km�;����b���
��;74uw��{#F�,X�a�c�)a֮ %�Wz�mI��^�q`�`S�^��g2���ɧ�s}�اnfn���eq�|�)���QROω���~�d�n�R`��,�n[9g��R��D��F*�RM$��aﲁ���⼼��������da��9L���8�nc�$�Ap}d�i�;�r�~Ɲ�S|����$��yYA;���{v��]Q��h�?�<��q�N���eg���E��r����c7�߿��3ꙈA���w�>�`2��ض:�Sk�ʣ����q�C�q��������^vj���}&���dߥ�_�m�P:m���hut�>Ǔ��;S�,~#>^�B&����P�״j"]"�k�n�'	���&�;�%�����ԑԑ����C[��l�E�;;�+,m���@/;W��_�g�t��<|e���p��Ց�"���/���3L�\S'�W����n
5�'ט�tv2(z��fAy�HK��1����ݚ��Z��(嵂Z#a�B�ɇ����9��_� R��"S&|D�Qd�J-z�B$F-A+�4DX?���'���A!|6�L��o�M�4͌�E��M���IS���Q>vi����:#��:��_2w�r"{��v����۵�\Fp�%�ic����?��n�-"��$c�d�a��ob�ʯ��K����.�>A�搮�������>0��>$�GS���^L^&cr;�2��"����d_��b"�^��*�p=�o�˕���7f3�U�4�������p�.��]�h�S�G�6c���:���p�z�-&��Q�es-Ȏ 3�m^[�]𢼄/�Zz�u(g��������׸������^���1e�?1��d뗜�.,���\?�175]u)�\�r;jP�8lW��W�a7����`.ǭ]��yӏ�펭�Sf��JOc�����Ysf�[pD�}�e��͉~��*f7�Y�߿��b���yH%Z���V��~1��S/\��C?IĠ��ݘ�P'��A{!\{a���S��ԂKɕ� G��{�h��|���89��T��R��V$��L0�ܟ.2� -?�T��6#���� FN?�� ��T��[p���Fh�4?�\i�q���{�y������1�>�@�ڲ�����jb��q�6[��R���D�_'�+�Z�2;^��ǑP�p��|8�<S��:aȲ��M�S[���#s���}]�f��ܛ�F���Ro4<rYLa�W�D��~ȳ'r��c{
]�ޣ���I�6��|�|�cJ��D/?��kQ*geD��X���5��k��?��I�_l��ZIB���'K�!BI{>lo����$:i���.��R�P���ÍW.��K!����&Ov��@�r�����0�U��:1Mf캅B�d*%s�svxJ'�K#�Q�ʵ��jR�1��4�8d��9K7QtG��Ķ7ܭ��[!�b�O�� #��ED�I����-ğ�	�Q���]Q̳�Lr;�8��oN.�r�'�<�#	{��,���ß�`���:�~�O���zL�Ķ�v,��(֌~�j�_%9[�����d�Z�qF�P��E��-g��Xc�%6߲u��â*P�l�7��j%�6�
��gE#c9���p>���7�vf}}�Lq�T��� k���پ�	�%��Bd�%	T�X��g�ƙu��K��ɿ���
�I��%�Z3��)(�ٿ��f:���Cb���_Qq(���P���>
�_F)R	��&|������d$�2��Y8,�&�ɊM�Vz��ջ�pU���� !=�K&ˢ����]����t�y�A�3k�?i�MR�w�a���2��T�T�Y����
�A�d��3H2�Mvd�	�E�]�ɵC6D�,]��%����w�rr�xэ��Fx�֫����k���x��мŅ^�C��&���#x�ƻ5��g��*��t�{Ӌ�o�����+a"f9T� �
�N���rv�����-[��YMЯ�/|�����vU}�߯0����U��`��&6���+"��ly���ۣ��
�?����Tp��}��0�㣋����[����s�=��D�Cϩ�@nf[��3����ϊ�ȗ���ޝ�	��/�Ωk9�YI���H�Ţ��N'ž|

�U��o(��i�4��ᆏI��o��f��Z��>�?Ȱ����dkRL^@��*'gݗ�v�Rx�ς�b�p%���_�����3i��&�5�E
{k�z��R��[��3�d-�-�^b�T��N�ڍ���d�ͬ���A?�u����=,��8�Ͽ�/Kf���v�0tE"�q?,7C��&;I��R�mfn��ڌU��x��zt�[K��ͫM��P��3T��ח@_n�In[�#QeB/C�E�SD3����ok���>j���36Hyg ��R������w_���������T�X����z65R��3�7#�DI^B��6ҳ�*�����2�<_D��X���)�]+g6ݲpX�~����	��ev�j���k@y�O1�<�M�~[�s+�~ĕ�Nqm?*�Yv�ɰ]�f*@��S�B�P�;$DXOA���<��EJU|+���7u�x�V=ȼ��[�`�U7lx^�/EU��+��&(��/�3����v�5!	qvu��m�#��aO�������c�'Z��k
�ߨ�qg������mյ8㑹�#+(��%��@Kt�3�O�r]����z����o��KL�"HHnG�g�������H�a?�x�HҴ:��nL�����0v%�_���-�Kt���{�4*u��ň�x�-�zaEk 3��8ς��G3����&e�}:I=f�E͋��b��ޛُ�=T�]�٠6�W�j���W˸�����Lh֜O/�;E�T(�T��	2��K6��"4d������6xp����V�������ó�h�z#�Z	L%�'V�ZU�7ea��ϳo�+��D%W�� (�;v�0�k�|�i��)����l�$�|�@0VXA�H��̾
�E���!�Ra�E��U���.Ok�6T�H�e��w ��P�âr�C�����ݖB��NP�����ck��p$|�~h�%������_�-#p��)��z�sLWѮ�U����E�l��x�$%��SWO����1f��OO�o�֒��U>�;B6�3Y��D�a*3�N�}���2�bA�ZUk۰,��m�M�A[0�$V�H-���=ؙR3G��aXl6��o���m�P��Rc7d�Ժ˻��#l�קP��m2<o��|����)�8���	���Z�,������/�G萤�9`���@	sK��o�3�5o�)��h�����[Br�j6tf�B��ӇJ�T\�CbT�%��uá�c�qy%e��l��z/�_�L