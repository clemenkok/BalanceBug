��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�!��
��%Y l�׾�NX�0A�J5�02ye3��<�a ��j>��B�q3������h@�J��f��)�d��f���-�!D���xv/�b��+���~�q}S���x�g'n�F9g\��3�O}�L<�@�G#���$$K��w�P�6��2I�ޕd")�W��Ғ|�!0Bmx����DC��%95��X +��,J�[�t�/5͜���?*@'���m_)�M���O��1�Wm�/������c�+��0�,�d8�ŭ�ׁ����~(��m',5�=,fRh@4kG��.�N��A�M�c)p�(�B���&�{��Wi��@m،F�|�����*WqBl���=��@_���[nH캺����]p&����19Px:�5�^)Qlo��%� E��7}�4�� �B�SӅ7��`$�����|����w¬�M\~G.���ړٞx�_0���PLY#<�̦����p��} ����ܕ׾�lM+y��Vb,F��ڃ��}��2���J�	lr^���Yaߦ"Ţ�`sFD�Sv]Vܾ&�����_2g���-�A�tuJɣ��L�R���n_ֱ�	-0B๏��>�ɋYq="�+��qb!�X.�O M6���@�9M!�2���[��!Ex1���f�m&�2[��F���D�>���L.���«����n�oS2��Ǎ�e��[��p՟���W8��W��C��9z2�������l�cE�a�A~f�A�\����eU��3��7�QI�J����|�~�Pv�fPq���M��̂EI�p>���޳�4;�������?�c�GC��"�G$�]�%ڸ�"����ԞOu6s��n̨1����i��4[�9�2wOw�U�@��l�� ��c"��ي�y��U�P���Y�:��4!.�r��������B��A7�y��?>�$��0��s���;R�K��LS��GcG69a���Q�JF��nD�%i����qwǔ�kJs���������?֩��_��Vp��6[1�v��ԭ�K����n�@$ ��h�Bݘ[�G ��
�a������ԅG�ܿ�����HǶ}��ȝGS�j�&�� )6yej����*�=�����������WW)�<р�e�1��6
�rfJ����4�eU�P�*��0LZx�][u���h��͕�j�4ܪfZOE�o~�$3g�S��I^n�ݬ�f��N��K+.)��C!��5B\x7.���;��f�2���Pp���x|zڀN՞`�풂�J��H���!����X'g���[5ʾ{�U{�����Q�)��k�
��ɢ�2b)��F{S"ѭR�&U!�*8��7�J	����o*:��5�]�2�vL&Fx%թ���Z��l?�o+X�u��Du���4���Z�o�V���$�Z�"��67�1\�(	+l��9uC�B��UepÙ�Ya>��">�nZ�m㧾�إ�₨ڀ8:x�Ȩ���%8Tz�-����8����+T����LYW�ț~�q`[v����ܤ2��E��c]��R}䜅=��挦�͈����~%��l:
���e�S�t��mR~J�Ĩ�e�9�P������[�Fv��^\|L|�钦[p&r��
\��E~Ls��}�\�}a�S\/�f������ 	�oV�O�m]�(��Or!j=�ȝ�8���9Y_ܳxq	��b� MEq�t���~H��������	8���Ŏ��2����j�FOO�(Sm��Z3���p�f�{�؎˪�^hʬ&o�D��{	�����
�t��Bfo�YK��vv�mWm��S*�ݶ��2&�wG��[���]F�9��!�}�Z��Fb��QAr��Yy��y�ke�O� �k��J:�=/%v�F��}�A_��?�R�R���!�y�vTKH5�f�k����|��p�oN�����@�B�/Rz�s	��)��#�W��x5�� Y�s��U->�q�G��'}���k,_Gm�,5�D!C����GZ �$�5��|��Cϗk���;��N@�lB��W�Ъ��-��4�L�����]nB�9
 cD�X��������ؓ��oW|��ں�d�Em[(jCO�; �W��o�
w���G���f���!�m��蚣o��m�����ƣ��"��=�"��^� �.%�iO��?������;�r��S��3�P��\���g;�
�s�,R��;8A��	�Ō�s|�u¾'��z�aǱ��� �=4k�������	�Z������b,9�L����b�f�+���)�p�����t�sk�L�7����j�L����޺l���=����)Ir}\,���W���X�#��vD���}l���p��$B�_"�υ��=�a�1m$L,%j|��M"�g�v��'u򈞹=�y�4}ئ�$g����SF��q& �Wp���v�Ÿ�l������:���Z��o��BJE��U97eC�:�pH7b���q��rTZt��Ä�ݰ��H��FWŝ�w�a6q��WA�I	���7�T���y*i��NG����|<ks�l��D�,́��I !/���l�'v��^���K+�
�|`�V���0<�R��^fu��L������ܣ�d�`NE���H�!������?�G �$�"�!f����%�ܗB,�v��e�:�N�~�v�p��������ľ�"�^�XEl��ݗӋC��jŇ(R�i��gØ�WF��I"�枩�=h��~%l�2�1t��Ǽ�}u�ƙ&\��9���R��4��!�,�¹!�;5��ӊ�#6��b96^Z{�0J���x��^M�mf��G�� ����j-L�������Y�:�(<;��QC�0����0p��C��� H�A�'�S6!jo����1���o�r^��GhH�[K	>JS�ma��`��0/�a������kG't�{Z���`�)Ӻ���x?�&k6�%:h������eϱ�7�Zd�`��l�����i��|�x5~o�2�Wjq�u6��;�O�B
��������L�>�N�}��SI�@y��3�q��V?��>���)-E����aMvC<��&�2�2C1���fS���K����9|g��f0(:��v������_r����_����y�*�9��PCߎ��zI�\1������{�e���z�vhA{�p	ټ>w����kK�*J&��"�	���$b����a��4��� ��n�_�tw��K�M������M��X�>�AY�1Rw3>F�y:�WP��<Y��𽵬�@�ň�������g����Ê�9�o����v�\��~���/�`6M��,X7��lm��� �my�ґH�Z3c��*�m�p�$�#*�&W<L,d_r��N|�������L���y:u���f����:�I��4��5�2�G�Ӳ�qR<"��"K���ܗd�p��H�4�H	0#��Z�!g�(-J.��dС��*o�;��_0����2I9�Z�=�]}�.���CV˥<A~��Ǔ���;����Ⲍsu��PN��èe)���HPKB����Ȱ�ay�8��>� ��m���J@�ST�<G���Pe�r��U�] ���Uy��38s�&��l'g}P'4zI��Ma�ʮ�'^�&��k6��b�+}��|�D�fU�Uq��Wx֮�lݢcUe�o�St����6k0S�]s��q��@w*ǱN���� �ErP�`��jgg}���;�j��"����mX%�(�7��-�ira�o����~�쒍�H��a����zL��eu�c�W�j| <���.�ڦ)�k^�crMI�D�\�bgZ��<�������Z�<<ϥ��d�V9C�����b��W�s	�yb�\��\1<���ˉ�E�*j�yMٖL<�>��]�hh���O����Ǣ��=�c�r?x\��Z��Aв�.�O���⻾[���}(L�����-3���IF�d�	U�gx~h����[y��q�;.�W�ò�ɵ�6�-&����k�ኆ)�P��
P�.�ʍ6��P[mvR�.�����l��q�.����V�uGբ��j���Q��yr/���DA�g���ڄ�W1�h��3�4 [�M=�������.�,����}�/�y���gl�7qcYf�Q���	c9f�5��Ȫ	��>]�X�*�!r���X9�0�xr VQ��Y(�^~�8`�7��E�f��Ō��6'zI��Y�\c܁ {������+RY�N���B��>��k�0��1�ď������u�3����&�3=^h)C�h��5�'�d]QY:S�S��"��9s�X֕�N���&��>������zz�|q��-q@��:b�	G��$m�Y�6����b#��_��X��%4��l���c����o\������j�>��5˃��<��w�ƕs�Lb?��m57}��1����=73�*wܐ�)��봯$��Q		�Ũ���Q�+�R�t���q%�^̀��K&�b�)��z�M_g��]V5�%w��ʦ+g�[W@�]s���%�{̠��������4�l܄��[`�S��]�Z�:������Y�$,��ք�����ZE��M2R�ώ�����,�A|�m���S�ܰ�a�^�d侇����B�1 ��6ug�F��_<M���,&K������0"+���-l��Œ�2q����25f��-���:��[Z�P� �bۭ����ZX:��o����VcVZ"0�VH	;glf���E��yxCu<qJ�:��^AOQ[�bh9�h@CX�8䕎·+�����5�Lc���X��Bw���LX$�*��(/%�,��	Is�I�!=AAv����bb�8_Jlz_��Dl��;��L]-Sy�[��`�H��j�ջd���͌����}�Hl^R�/��+���m�s�&�R���=yjw�]4&"����G �R��G��׿ ����ZmZ�����8K�my|��Fs�'7ݟP$`����\�mH ��B�a�1��*{�T�k�����7�En��������+Pam��{� ��U�}e�p�!�����Z,4�j��
��ԕv�v��'��;�ʆ�@~�#n��x�c�Y�E��=$qS>)3���n�?=&/�>� T<~2�2(E���Ϣ6��8�&?�vQo{y��$�h�b=��P��EH-��[J��%���gd��y.�"�n�4%r~�X��]�Kb����ۤ�Ⱦd�'b`�T��4́ƃ_�������AB>�7�$Ɗ�,Ya>��k�N��)b=�y��� 7��:�9�B�al%B��dI1xh���WW�3a���-1;ZaX$��@�+0�B�ݾ�����$ލ�⦬���O�z�#��*��/�(���v�C��*j){5�a[�]n��'��xVs���%;�zZi�7�<(;^�!�_�����'=�!VHO�'l�
@H�u� ��ٿj�w����]j����X�32�-Xa`�Id�X�UY�&���&�Sli)��R�`\{���gV}XP:��?�6��%O���aʷFVNj��f���YN8��D�.Ȱ����=�X'=ǜtb����Ʌn��KU񡡉�LN��GND��ڐn�>A�I�m�W�o_�����ޠ��[8F�Ǫ6��@C�b�A��ݙ�_��i?Q�����:X�c�1
�MDl�[0�t��ȉ1#t�;ޔ�a�|���y�/t`���C��D��Fr��;��z�����O���[(J��˥ T�����I�c�����I�Kg��6��k;ߨ~WyE#���D#<�%��:pZq�/� 镏�_��SEJ� ����[H�/ڳ���m�fm��u�㦉�I����Oѭ��Z`#0���䚂֖2�qo���|r��╢��ƚ��\�8w�ԉZ/wT��5��ki�q���3��f1xG�>�!)��f�z&�#���g_o�N�b�v�DR����m�����]º����Qi����L�ʥ�_��ڀˋ����3W��������0�f=�&蝮�(�B��ppq24f"T�dl��'/G�t���+�`(#�*>c�y�%#�T;����S$��6N�7/	��գ%�F��!�4�ԇM���l�b4�Eu=�G&��օy=[U���'�r�g�W��]
���Y�����nt

%*�u�WCċ},f��.��}ߓK�if��ݿ��q��t���lӴ�62�6({I�����D(}�)���{��7�M�}R2Fr,�����C8ַ^�=�I��dWĿ~S���^߃��LfaMY?_�G�C�n�_T ���
�i��R�Y%��o�;x��(@��f��=U��l?+�f=9�����i�d�b�_�l��8�Lȹ��5�{���!��x=�;܆*���SH��)]�g|��*՚��b�[�Gͪ����c�"˳��q/im%�OX�o��\8��7 ��ĂR���W�mǋ��>N��?�gÖ��c^�k�|D�=�/�6"�v\/1�����`�d�����D�������.�v�^��î/"'J��үb�S�.��:'T�k,����I�ŌoK[\�X����/��1N���E0����z�6*��'�y�wqWݾ��J���B�IY EFµ؀���v�cz6ک��S�U�N�h'��5�Hx&&bz~���I�5�8���e��3���B�n14eJ�lrLs��n���ۯ��3;N�i�ㅽ��Z����l��U�7>n��s��d�(P����Q���H�%�U���2�:ɕ�O��T�#�B��K��e���aDv4�����dw���Ncp�uhT @D�X!ci�E#2r��0Q�'�s�  �_97�j����$,7v39��sz^�p��7~dA͚���r�K�P��\����e�b�Y��� ��(P��߈=�@p������2���~����{�v�̐�O������}.#���N��O?Z���~$�l��.;;E�U�B�ӥF3.$�XŅ���5"�=2cj&*���~�c��j�5�[o��ye�ź!L����|8~q�P�;]�L��ټ��硭���6�\q�ɓD&���F�Me��t�{|��F5xV�A�Y��^yס �paz����H�s�z���*ts��k�''vۨ�c��'����1�X�Ax ��
j�o{n����R��u��O!^j��53FQ�s�����uh.��F�+��Ve�aA�FQ�m3�A�dU��|t��|Ç�� ��|���)��ĭ���g�y��>2��Beޙ��*�2`z���q#R+�@�3M!���R����=�L�v�(4�v
w�s����ZR3���+�1q�'![�cPa6���8[�Gm�����[ۋ��F����C�G�V&M\	���k�_�x��G|���%=	7�E$�Ae��|qׯ��c+>�_9�r*�	V�v^�}�R�sy�c�_�0ι;� 6�Dlt������b�WQ�wڦ��i��ӏ��q��Uմ���]�I}������<�u�v$�l�<<��h:��^~��g�G ��,���h��Y�R>����K�����+ȟY���+[�Z1�0.� ��a��rL�XfJ:?�DFH�Tè�U
kpY���☉��r�NTs�T��,��WBU�R��s�FI*��:��G�Ζ��D�ٶW�U�����4�/���^�Χ
��6x���Wp���:aÕ��@�Y#�|���+0.m��t�>���5�
��@���L�(d���(x	��Z�V��N?���wI�瑣��s��\)}�`����&�J۷-��T����g��j����g���.N&Y�T�7-R��d�m��25�n&����re�aF��D�w;�k�~������̐��6[Ea6�O�D/0̻��(�F3���=,hu���a�	�Aګ�g2�Fb^
G
��Le#5V�X���B��23��wD���2��Z/���TC�l�F9�������GV�SAȠ/�.X�?��2�2�f�����$;�\��¶Z�5�3H�:ĩ���3'��| ��\U����c��*�zh��	�R~��o�w��g�x�\q�1����ͤ�
&Y��[�@�3w����߰y|O
��D;��/�[+ϙx-��h�!��kG�B@!1��ߦ I�����sM��,R����>�O��f��H�4O�T.��� N
�d� .#�p�`�q���<h�����L_Df6m�{�����J��`���_p�I�Պ� Pԫ	�)8.���r<j�军�膱N�1�o�ы���¾u��Y۱}�eݨ[9��↹Hb}eϒód����*��zt���ҝKߘ�����5+�l���J{4eO���cǃ�0%!�L��0��tq��j�:|h�]v��:���d�/�>�ع+�l���V�bp��2�U��%(o<���]mc��c� �[��J�����%:#�U�ď]��VM�A�X`5,@��O�PJN��;*B�s�j�0nS�� ��l�k�v��=��_�p1#cT̸];�Өjd�4ٳ#�4�C�h*0aL��"A�,\�����&�dSǋ��H���?5�.�Fƒ*����_��������y*�xq����
K���TؙuY�=�����P|�\�q��^k��kG�6����H<gM2r�`5hye�_�$X��sLe*Q����p�������y��d4Y�����PU�f��m|��Ll�@:��c*+��wp������}_�[UP?Ƴ>��j��|��,v{!�0�ڼ�mgs�����P�z�D8xͦ���D���(}_3
���P"3]��4����=M�1�V
/�8��yX�r���F�4�_R����B�u	��o*X���_�pM?�p@�䵸�h�&�DlAa8�GVbU�+���W�N<�x�+K��:����Dƴ������'��p�>�U�n���p^�D{Nj�H��q
}ͼ�Z���g�Ni�r]�����G㝫�LV�pa�*�ܘ5��:D��K)�; �lᤏr����*�&M���-�����;U�S5��C��xP���F���P]��lw\Y��ж�)dփA�v�ڏ˫�ZI#���˝9I�B�Iu��^�	�Ҡ��x���c����0��d�r�8�:)�f�-9/���K�x�R�-���`��2�s�&�b⑛jkd�sX�S�s�����R���	1t��KA2�fF�֤UK��;q[�u��:�U�y�u�:O�{�%�e��]��SEb�k\�;�y��i�oh�>CV�]9�Y�(e�<�iON�i��~��[�%����y?|�9����L �f�j]�z�������1��!���q1���Һ�r��,��,�f����B����m���Wk+.5�4ZLl�z�Z�t�+,$o}�6�����m�T�@�&�pm�j}l�&ԔRcCN���뢪��d��r���L@�R/(+�����ȉ�ɝG���|D9d-���������@�{�;+QA��S�x4�j��aK�79�2�#[�u��]u��{9m�MU���^[ �{�Oޡ����xG�]���F%�r)7�0�:^������w�)�Z�O"���W��2�h/�K-��%*�k���NC��������<�Ra�Y��b�>�kqF� �d���WR=��*��[��P�H�1%\o�$.�3���P�P��I~��uA�X']J�B��7��A��A��&4��FO��!�{S̨� %5ƞ��W��;#��0��\Q5`�x\e�}k7�'|Eč���(e�'��@U�Pk��JI�Q$c�Q h��T�N7��el�Y�ₜʻ��U�Y��	JB�G�Xg�)���ji��Ѹ��i5a!�[dN�=a[:*��n}�*�W("��!��~P{�D���d�!�2����%*���)�C=��b/.��%B����jO����qpM���sws�8t\_��m���+�VP�wH��]a�ί�H���@D<΀$�ϣ\ i�&c����;������-��N�]]�I(&?u��RM��	���,��p$&���b�م/H�O2M�5�Z?/���%�9��:��I��7r�O6Q�:�`�?���dS636Y�N�j��CuWq�[ز�Na�9`� =���%W[y�{�Wrˠܜ	Lu��7Y�q]Y3�N#ȯ,oI� r�J���IT�c��p]{P�q4��X��Q��},)Fx0�y�x�X��x�r`�U�؍D~L�.��1W�Re k.h��2�M���ܿ<g|�|�F��C��T#�߶�\�+ܰ����L��d\�������x�Z��3�@XЂ����>r}�~�
N����Z���2��{�@���Q��o���Y�A�x.���:"z�刾�'����V�Y:���r�E��27�w{|Eşg!�ƺ~�5>>������O\v����f>��ο��5�W����.p���8�"����lA3�F�N�F#�n:O�$yFc�u��"�:��d?�B=��'�q��I�1:�R\�4����r�2�IPz[�2kzP}����;�Ȗ%j�a"�BXdC2�m?��I��qW9x�*̎�*�rwOk�B����>GZ�ed�@����U����*��n��l�~]$�6�bV�&�l�y!|���M5<ɸUfC����*@�
�l�D�)�\���ݾ��`T�w���w_�����TϾ?F�������ȹ�Wa���*<%j�u�}�}�E��Bt@a|�ĢD5�8 �f���1�����LC�~?�mɊ��3.,���*
!+�����<u�=}��_��b�N� �i�����+���p��3��e����(�H4�?��e��Z褪�VAO��ħeDސ����'3����(��\�at��'Ì�����%mѲ��F-n����Y�����餐͂�̻�݄v�`��wZ�*�/�����
5^�I�c���S֣����3�fo҂=�,|t���������JJn�A��"�&��SU��V��$�k�d�_�C�5,�&��*��<��}�OC\�WW��@�ݺ�I���k������m���-����[��[�>�H��� �� SYδ[�?���8��ǲ��Pm,Uz��y�*a�/_�D��?v>t�Ƴ�������OV��Ţ/�g�O9�j�Z=�[�?G9��z*�A/B�Zl��>z�p\�i,�wY-f��Ŏ"�5�"�k��R76�iP0��o^�P�0��邡.�|��>�&Rw�5�]2� �l�"�#�r��&!�y[��uTW�	̹�oe�\�蜂��`L5�J��p5a��|��~#v�.EN���i'<��Е�ac �*���h��ɦ��i��s;ՅWmb�޶���=�"p���5��J���^O���A��8���o�e�A��ڐ�"�W��4��\�ިN�{��8��T��I�����&��+ ��j��N�^i%z�bGV�D)�/DtT��{s�ٜ#�n|�'Ҕ�А���������<��ϴt����#@�3��-�'3��f�sxg���Nbbs�P�����`z>��T7�(���w�FEs�P�M� ��G�)x���*+37�p�"S��⬼>��=W�,�s"�q����k(ᩋ�f�i{�k��Qڑ��'ms�(��g��:�1�Ǻ����/K�Ц�e�ӗ�'�h��ˊ.�g��F�w᪠�O��=�z�2 �U����f��Μ��d����0�*fo��$t�}w�}}o�C�F�,�+\�B)>�[�����%�Ƒ��&�ayv.8p�i��DP��vK����$9fD�;7V��\�RفJFH��d��R��V�>��9Օ�r�KL�{�k��5�`�~s��"����q�(�Ck�o�O�F��%��3V�
��^�X���x�����􉗢�^מ�� i&�X#,Ar���V,J��F?¡��z��L�: ������@�6S��w����\�^^��R�/�3����z��t��I5>t����X_����wi"QO�lpb�l���D��e|�g��p��i#P���p"]�R�uyR����{7(:�	�����/귐$�3�
�E����g�]��T��d�SL���gFE=��"���.o�c��J�N�*����#gR�,��o%Y'�O�2��f�aO�7N��&H!���:ߊ�+eG��'Y�%A-�׎�B�� �%���ȤL>q%��ԨH]��5�n7w��M��Zk��=hsz��
�,ˤ����/��-��-&�w��%�v�[���y�D4O�`g�v0�ək>�O��r{�1�p�D.��~�a�k��T��b.X(�7N���?u�GҊ�l��3׿�K����@�<��y�yA���4�{�%T��+v�k,��9�"��LeJ[��������0�~"=��Vpp��h�`��U��e�nWvtd�0ڑw�>K3�qn�DQ���"�[��l> ����Tpb����\�\���tZ��!��4���"A�3ym�c��J�N|y�^�����E+M꯾3�i���K��|-1o�B�Wl@�yݬ���ꑯ� SA��m<�A�����D��M*;�>	dA3ض	`9ʭ�f�?e��G��}��gd:��O��R���KKc j�""5y�(�CvAvE^I�1�7�����2$WŲz��T*�����W�L��n ��T�p��j:�X+0i�o�h]�]��[/��˘�D����r�n���m�����Q�3�!�:�4}7D�ς��3v�3q;}#yu�>	z�[F9�y�h{�:�x*�X�Bp���0�[;X�NЌM�ns7��>|���c���E��g���XF��F��2��+ٞ��?�b��H�¸�]K!W�T����Is.��c,|9�(A�n.�;H�p��9�#����m�dsԕ��6�i*��1�� ��"�����:�|�� &�c�٧�'�ߕ��9����e*����l*��{��;�(#�D����ۓw���������N�f�?1���%�h[���\��o¹ ����iR�c�����r���Ǘ�^5dJ�Dʡ�ܧ�n�A��7���Z6�`� M�=�j����zu��1��S��&Քl'��W�jx�L�@^*¥q�1���mm�b��YMu>�,�8BZĲ0P�bZ�g�R������{��cJ�x�	��ے/z{_��*3�����g�:g������2�5o��ln� S��_ܳ�]���j$�h7֖JG|&fuD����_p�ş��_�lv����֟l�X�꒤�bN>�8Ju<9茦�c������.��*���{��@��U�Ky��NH���ڊ�yC��)x��
K5���!3uߟ��:��Մ[�d��cv�Qs�9p�b^ �cbT�̯�Г-Θ��`���9-��%A���:-�h�K�����!3�,\�#�K�<Gl�ۮ��sr9^�z&�\� �}��SV4�T�뚐���A)�ׂ�ʪ� �?Ϛ������ �� ��hk=��k��́AN��컬*��m����/Q�~ޤ(A=�*���5�x7QX*�1� �;�>D~�C�P>��[
�/?"ƫ�����Q�I�m=�B*Ht�Uw'�3�Q���ޑ�ՁKG C�խ	�i`�$~jh��S{�!/YR�G�+�A{�	�1X�5���W�p����3��Fe1"p�gs�ܬ��)zϭ�s:�B���F�vsU<�uuC��LǇ�*Q6{9v�t����[A�����naR O�q���O�"z�S�6���J,O ���� W<������j���K}}�2�{�}���P�� �w�/�H�\:ˠ�r?���h�"��@=������>��^Iٹs�e�����Y���-M�H�p�0\V�N���U�f;�����)�&3](�ع�����K<m8P|3�U��f����S���ܸti��)�R������~�\��X^-��\�i�9
A�oZ"��!�	��_|�f���E���������v�C*�	�C��ל�.]�D\aŔ2�^���/���e�� ��G������a���Ҁ;�Nj�H{EtC�ֹ_��=��es�?l�ʬ�������� �?m�N��luD���9��b��hۆ���⛹�B�&ѽ1uT��"P`0�DA�����n��OH�>q�$��t\}/���[�e� ��PZ�����������q��,R/��#�3d+�ɩ8:=�5�04�3HNP_E��n7l�k����;- �����Y�l��j�D����}[��r�|�ոg4��"?���L��\~��_!X�̂	��@y���pB��8kmp���E�C��j�Yf�%PrpA2���9���E�	���B���&������w�&{f傒�]�",��r�.�d�;��æ�<����y#У��r�o��h�x�a�Q8�%�{0c� +�\u�E������ߣh������3��@xx�l��Ǳ?hho:� �{:t�G�Ti�gl�c�y'M��}q*ۚ��
c��^fr9.��yV��IXS�E�Ep �.y�(i1]|0��T[ǵ7�d���娎U��(�*�G9z�$<MP_��@��z�W;�{.[�6������}[tk��.�]�F�c�$�Q<M�A�l+G�&�T��w�+3��!V��	��L�G�9p�,4����9��U�Sb�;�0�ښ �U�	�N�����j�>���&��gc�[��9?�-�%�v���lr�;�$��lC�˫��$�|�BK��<v���|%CR��������pV�1HA"V��W�[����f�����C��C/���3�3s�V2���>-T�rm��]I���̌M�?�EoD+��Kx2�HCg�0����VQ��n�>R �<,�J�@,�[g8a�g�R�x*L=p�n֙{�׸*ځ��� %���F����{꿺y&��c&��/��j����u�^�c�&h|����wKrv�G6�ۋ��8 Us1�ka��I��}|��U8�b�";�/Ƨ���| �<�F�B�Җ��J�A��.���g[;Q>._T�L4�=,���c���%dyF��8!�)|�T��4�Yx�� K:�ъ�����O����x�ϑ5�w����D�X�JE2���y蠞��������S��O��#��|C�^�o�w淨w���~��?�y(���`�=.?b��)�=:�Wj���@E�| �!�����!Ywh�߂�a��5��' (uSf����=��n�1"H<�v��Z�j��Ow��u8�I����t3���E���j�dc�R��-�D_b���B���k�:&0�"SY�`i �9XC���G@�������A�o̭��`�_L��>_�~����Z]i��gd���o����Ͱ+鈦S�/2a�Კ�![���iV�� Xo0
�wռ@�]c�k�I1�k�#�F��Ђ��X3$��p��Ne/ЫĴ渃��.��%����vx�9�@92��?JRG�<U��8��V����BÒ9���"�΁Q"����𡭎q0���%�]L���� �MT���|�;���k�ŰG��ہs�����2�$�U��z�&k�D)cZ�i@�/�"��f�����&'�{b��իӅǁ�x�Sr�)�: ��8�ŗ�߮�Y�� 4v�
z|�?Z���e:���(�Ưų�P��.G��4�9��Έ�IAV��XT�Q3�4�]b����8J秽j��r�j5��_`��U��I��l�[�kw_G���۝M�<�k��($�S<o;�:�g�})+��bǾ!*r��e��U��>�\(�NIɻ1��@��R�&�����-��Ă5���x���b=�#����)7N�8��2$��tEk���I�9�B�~&Rn��5F�@��=��2�=��=<F��]Δ����FG���Y6&%�Uf�0��S�={�4��hʽ�ŷ����S�|,�����������oP��r�%Z��^z�=���{5aי�H�u�"�hX����'[�t�W�E��w����o���B���������I'��Ԁ�]�R�Y�� ��0�l�YyS�yE�O8�ķ�s`=�	i�	�싂���R⛏����O�d���=ԇ�-Å~ y�G@��F�_�ioKS%JY_-�`H]�w�����`{$��L�gu����Z^\*�\�(�,�f��į��?Ƙ}֘����˲�}�ZF��s��z��;�6��"<��f�CP;I��7��;)��t�N��c�w�,B�b:<��q@H�C��=�Rk�ED���MF+��@ n���������5�Z�(\I�K�e��d=�ϖ&S"Cs:��Q��m/"5��� X�_c:'��ڱ��ΐ����&��RT��6���ܞZK�B	Aq{S#s<��^�������%LW��s��l%>̒޻ᖟ��/V[�N��Ѓ�P��~����Fv��}�;��c���؟ҁ� jUr�In#�#��y������{"�b����=6A�V-t/a;�q��kn�Q'hY��JI)��y�BD�R�����?�Z[	yg�U�QGz�j:�{�j��3�a�{My2�+��ȍ��k������ �X�X�x�ܝBRqH���9)~"�F����� u��4t����W�[o���=�Yq���h;j��0�G�dL�A�J�Cz�\���[�(IZ{>7�]�-��W�w^~��Ű�W
�б,�ד��R֔�X�J�(e�!�0t����nՋ��tXQ�
;��u��iN��EɰFG8���-�T���I�q�/K��J^�/\����#�Y'̲����kZ��g�*{%��(���4�)C��Ժ�^z��	�ķ$����t��
ߝ�;܉��0�ු�g�t�r�S��6= Ma}+ttHhë9h��zW�q�g)Q�>3٩� �"Z'��AB�&�h��A��!�3�ګ?�,���m�9�)zFR!�&&�j�h�����-�a�u�ɷ���#�Z�m��ۮ3��U�����T�֌���)���R�Bx�葧\�ly4�&�zB[��|�C��F�aB��2�J��P, �P9�?�+��[I��6b���y�R�|�V���2�^��G�:�c���6RQ ��\�N;���6s��w��ޔ�ˉ(�맩��6	�~��j�DÀ����g>3�N+7�Ә@�`�("����1B☆:�J̛�4�2�F���0r!S��6;���'�,VL���+�Zj�{fW��1|݂d�ۛ�H�0��C&�l��l2�9LyG���I���H�P$ǈ���r`
�e�:�Ȥظ�ʻQ�������aǡ��;��0��Y�����ƫ�!��.|��Rݔ��,�u{�d9�g�馑�K�|����wًݱp�j�s�Hֳ@y+���=��\(�t���/�����!(��BP<Cr�@��&rc��{���񡰼P����XYJ�yz��Z�s�U��q����z�y�y�$a ~�DD�?�\�T����L>��զ��2�vcQ��\s��ɪ�������8�@s�6*�(J����ɭݢjF�Dh���'v�r~�p�������H9μ��f�xs[7�1�tЈir`cr��J;K��#����7dC��3��c|�g�u����\�SÚo�0��+����+��G�����|��6���O�ܩ���uG���9���� �;tfM%��7˭��ac�p�'�Eq���u�����g�����у����^aϟ�[yY��u����vc���퀀�b��|��5[�NVn�8�(dn-h��w]���vF�v� �c�����Ȍ�u?:��$H�6���NN,���� %�] ��*�>�7�Z;`4���Cz8!P����Ɔ���
k�Xj����o����y�>-���
����Ty_\�p�9��{RF��]������P�B��$��N�˓tN�5ҽ>�vd�7�� �� ��J�H��D�@?��;Z�dgE�u^�Io>+�����A>��O�D?�_���+�S|�_�׷�� ��CВU�<��׽K�������q�s��'�c��Ug��^�ơM3�|�V^\�TS��Q�Xr=�R�����j��>~,��v�Yi�[g6+�-J���\��e'%DE�l��bV�*�j����ƥ�]��-�;d�<��UA���s}�������f�*%��].Ԗ��a�` ieG��h��y�*�S��5�_�9B|@�b5F[T��f��Jn���R_:�0*�؀'����C�3�}*�@�3��ć���}<lUNG���?Hp����[�ܵ�G-�OP�jW�s�F6Mؑc���H&����s��1��_���_�H�ء���z�P���/'3�E`łE�pE�80m�~�r�o,�3�p��o�6����M�1 ���}G���P'K �%�'%x_��7�b��tN49k�T�׾х���s~<2���
"Sޞ��J�"[m��/�(F�Qo\ܐ�XQ"��z1u���E��^���x�/��A�� .�N��K��S�Y���*$�G��. ,Q'�Ҥ��jb��(|5�Yi̩��]�W{d�����g�אe��
Ϯsr74Yk3ހQN�Tл��IN�7�8I#Zvq
r`�t��P@�0*W���,q��u�9khՙ~gOL�ܚ�ˡC��<�����y<T��i6ΐ�����FI�@����5{��+me���J2�k���;>g]Nm�-�1�zA�~Ŗ"�e�!�Q��
#:󦀏���0�R'㍑���w�<�)�I�������~C��FC�_ĥ1\�HL��-Sz2�I��G�����ˤg����F"�I������4cWlJ�e��EpP?�8�G�S��z[-�c��Y-F6l2츞0**
���M}ƛ��"����2�)�bҺ�{�&I�^`?����Q��v� a�u-V��//[uc�`���%i|=��j�b�ItB/I��� L�W
kL۝���6��	i1��헔�,k���g�<��1���^�}ɥ��՘��B5dI��҅���)�T��&A^�|>G����r Ia+c�w�����v]FC~N^�k����sl� �h��!4u�yhO�8��8|��9��]����E���
]�gb�]+��V����_���v Ψ����Ԃ��D_���L}��rIf�4��L�^���y(i�&�S>�)e���B.�Q�W8ƍ��Jo�n���i�_ij����|�ə!�$�<o_���ħ6�z���*�ڿ��lĩa�&ɵ�'n�O�=�9�2���0���� Tٹܪ��ΛƇ��Ş����XG<:%#��۸:�FJU�4/|�a��du���ڶz`�9vm����D����/Qo����/�����9^����&��p0��ȿZL�R�-NErb��Ӑ�O��B�#���Rf�Ӫ� ��c~z� �we��5�t������?]��C�k���)Fӷ��Y�A�4���ˬDN�A�`a�u���z��D�o|g��kkpr�z�u�K�1F������"��/x�}��qyaC��� ��N�V`:u��B5Bf���ZS
�+�A��[�{d<��G�2��a�F)��f�2�i��52se�m��bM/q����ʤ��?�<��+����J�w���y�Ll�Ogt�S�t���Ly��&�95�:�p�.���J���2\I��f�n�% :L��g�#Bj�X�\�q�ATq6x����@�� ���p������{���4��2͍uL�T���}�Z���#x�<i9�*9��߻,!����������I��b�heP���C.íƳ�S0&��� ���M2jb1��_��6.���� ����?[3�r㡸2���Al�-?޺���]��|�z@�5m0{Z�wM�e
8	d��DDCd#�!��,�@��N|�i�d[�AWL�)����Cv�|��f:>B'�x�l�w�c�.���я�����<i��l��Js����-o%�G���7���?���\�>-w�^��0.T|�a��$	@�fw�Ɉ��LUp`��き8�=������-�΄������D�-�c��t4I{��d��t3E^
��w�",�-����{�k���ԥ-Zh���ֲ����a��������[IM_��W)������qd�Wl/��0Of\)B�0�x�t��4*x�h�G�.[�*�#_��{��y��6"/}���kN`�؀}X �2�Y2>���,2��lEj�&r�"y�� �5{�9Q������h�������p2h*�����d7e����|+��'%�
�vZ��-��Dn�'\��'I��v
�G(�opts̆)偁0W����_��"u�[��)�єE��C���U���Ņ/�Q�_�Cq�q$����*̯�q�'9n�c�MG��"�vo�٩^6�{,(�����yv�4���%Ve�Lt�m�8����A�ڧ�5l	 ��/���WB���|�yWn�N}��N�AYq�}��s��q�P�I�M�f/Iܮ����j:`���{D->�R�H���r(�?�Q�#\=p�E�qC�-��T�26>�B}��7��AI�#qpa����8��Z5V�.�n�32]>w�st�O��Q	�.Į}�'�$Uk�}���@�KǊ�1Vu"��dÙ�a�q��T������Jw��[�gKS*��d6��?/U����%�R����n���U|6~�����bZW0b��o�z f��c�恒N�,s��R*��R�=��̙�Q�4&SKAN�Z�XJ���&��1�1�u�+H��ՄF>;��)�K������,�%�0��4\�*�2ve�`C����M����%i�.�"wrF��$i%4L�w����k��%K�~8E�?2���u�$8�	�sT-����?�f�@�<�l���ʡV�#�R���{�� �����3+ξ6�&$M�S*Z�:~��sP�]�{��Ԋ&�
���0�2�({Fe �{	�}U���`{��=n
��PLY)�B���~ŕ��@�o��_<���ZyzY�J���;��lf8��h0E�>�-��o�>�Q?��rP↦>l�R�JC�d�<��SX:���/3�NsI�
��Z��W��e�g����\K��Q�L��<��n(���M0�Ҋ4:R����W�[+�C#�U^��y�V���&�c^\W�%܇׸�qm�-�����.�6���Uu�����s��;ylS� ���������z;]�;𞝸��u��-�]n�R�������>�s>��p-����/�D�Ī���}���1��C'ȓ���i�] 3K������x����C�=U�yQ���{��1���-2��(W3F㹸�f�9q�I7c��n�rX��x��H;�Ž{`�n3�q^����	���E^�٢�����ܟ9�k>����X�q,����3�4m&�:�N :?'���L"8��u&`.�%e�Id�ٺ�݄����Ĳ�_�("���D��$���]��������\ 7͕�����##0���1xu����d)�!����A�'� Ü���;W�#�q���m��8y��xD�����
"����Yo֧����(�"��2����B�٠2ݛ�OV�~��r��$,J��w��_ʯɠ\K��g��&�{��?� s�����WAvB9�m\+�M�$N��f �JS�� ;����xI�)N��nV`��=ˊ?���E��;gZ���.h��ul@�pŝ�M@#��(�&X;��%5��بP'�yU��c�bO3�*	XӪ�߉��o�׉jf��%8:M���I�RV&�����[���/oH��;���lP@z�7�9?{�:|E���;8�d���c��dGk���Y��ȅ��ٔ�L.QV(�V�	Vg���)Iy�p����q6c�M�n)�DI�I�־b�p�ͲF�8�O��律�9���g7� �[�y��l�~p�%*�[R��&\!����"�j��.iF�{�<�8Z�x��s��d�9���`噣	�w>��+ۣ�M���T�J�yj���=���rH�˺P�
*b���5�S+�8%5�ݟ�`��w߃$@�B;�h��K ΁^�t�a���]{/7>��8���5������4��%����ꏍ��)��ʿ}�k�����������y�;.8W8k�q1�#�0���E�)��*���P3��u�1b���KP���}?Ԅ��9!�e����H~^��T�q����L�2��p�g�#��1�)�?���.�-���ߔ`$��PQ�B�+8T����T���2�*5.a};�C�>�\4����<��zZ���> ~?�Ԥs��l~Î��*3���(�.τ��Z��%ď�R�l��-ƕŚ�	8s��N�_��;H�{��w,$�[��)���3>���o�}��zD��y�D���R��;`��i˫>r.�1H?x-�B��S�<M�sD/<�%c��l�~M:�<]#�xB#��hd�=�,�ɭM�p���> �3N��pǙ�,����7-�����{�
o�:�w�E�$*���{�{5&��_�ƮT��j {n)"݊�מ㠮g1�X���HH��R��]9&%. �ٜ �еУ��7C�E��v��s�%����y��Vcc�I����F�[dӁ���ndJ�;ѱԁ��{�;�@y}�?��a��I��CB*��Ŭ�5(�Ɗ��Y�ׯ� �\ it�4qw����F}4�4JdX����J9�H�`f�U����
j{8O,A�u��XA J:>�#��5,=L5ˋ���7D�$zS�D�~Z���?�yR���C�!����x��-�z�KO����gZ�W��y^��gU��O�6�ˡ���P�+LY��rx �v��R���ݥ��~��{FL�	��of7�C�,[	����o`��k]���$�K�̄����X~~wl�on%�=�YS��M'`����IL�Y�����tPH�;��Cz� �b]�-��� �u�|&'�H�I��e�����9�k��w�V:��e>Ft�z�z���gfߙ���J��%>9"���N��`,̑��Ȳ����5��`&�! _�0��}xƵ��W��yR�z�wbo�,��$���)}���*�@��JR�/y�!����A�g��<��o2Z�+:���r'�I��}5ٍ��:����Jb�!q���Y��e_���г1�����u.#��o�.d���k�ScΩkC��7i��kա��+uZ�~�&FNԾdۏZ~�	�s%����T�
c������'f��q>���SP��*�����7�{`���B���P�WL���Xs p	�Y���j���_)��NiY�b1��׫� w'?�A�p�Z�3��{��O�P�\��?�A��f���M�a�<j�q%`��@����^i�k����u�	\��D�ŀ���hBomAU�[Bzb���]i�Oy�3u��R��]�*��'	=�%�"
zS$rWh�H̯��f@�^�=�5]H�Ƿ�n�Ŧt&t���/����7��
::li���vT��_V`7�E�M�RI�iia��6�c �us_��eU�C�x�%�g����@��t�c`��8j�����?��x�næ�)�l�?r6�sV���>ZF�ݜ�J��"*Ic{��?�V�ՍP r���08B�����2���"�۟��������J��(��3��6�z�?�?vGӺ�喼�����ڈ~����PU��DӞS�x*=W�OV�N�����P�v��yc��2��ꝥ*v�XSZª�0��z�H{8���Z��O�P\x�i���䃪��V�Z<�lg�m���Hd�V+�[��'_»S�ck%��c=B�U�1	��f]��)�X���?\��OG�����#1Ӄ���Z{������3�&�q"?Št�k�E���/,�j�%�k:ٓb���)�J�Q�����N��	֧.h.ˡOC��H^�V6b�R���X:RYI�׈�Z)+�Z���DR�|c{��G.$����ݝ�8��q��
��A��]��_���E�������b�Q"(2�m��Ƈ������C����jjO���JEm�x6�9���q��}��$�S����؆���zv?�Nc��J�+]�]����)�dx�������2Q�J��f�\Z�vU��� W��;�J�8��٘)��>+�n&�/�caTo��Q��J�c��!S�3�G0���ֶ��XtJ:��9����'����w�[[޽�1,|� 3�H��{�x�`��ҾȜm� Sa7��z�i��Kɱ�N�0Q��& � W�����s�g5��L�h��	Q���_��y�`������BbtY��TV�T���N����ۗJ�91��S��q|����Y�"��\s�lcʔ�9a~�ڍ�&Р:W6�j�A�~K\s��g3턽�<�*^bv5�7 �Z�^�=-�I�迴5���9�w;��ne�EB��P�aw�9J�����l����49\�Fq����L �T���?"�;>l+z�B:�Soy�QW}K&lm��Jx���xb#�^�NȚwgsx̱Z���rx:̺GX�&Ѽ�ȩ�WcA���z���"\����Y˞[Ҳ�B?L9sH6�4S������Gc�k��\O2��'���al�O��ߝ�4�e9�5pX�Y�)S��\��(IP�	���Z�v��Z��vCq��x��G��7���U:�ԎlT]��YJ\��y�r��h��4$�lF�1����f���N-��_��
����+�˨�
�i�u���E&�E$��x�kE��jO�Sߍ���qy�vM"��X)���;A1��g��|�w�ϖT���H�,+��`������ޒ&f��*`?z}��41��	|-����⬐Ǳ��b'� �s1s���~w�aR-;��$����}��of�6�E��R��ނ?��� sD���9�]�\W,��<H<>��� .YO3�1KhiY��`� ��i�"�\�:D���tdȷ��S���}{�U�{9Ȑ�q��t{��g$3���s����<����W]E��v `�\�p���a1�?��?���[��j�Σ�r���?Y⤵��E��V�Ӕ��4I�h ���Z��^��<�k�)P9K���~9gߝL�r�| t����2
�9d�E��*�j���Wp�؜���@lݹv�ъ�Y�!U�Z�o���~�"%*hW �]�%�u�#QE-��u/��րzWK�E��$\���0P��XJME�gi��%����v���z�7��"e7�)8�Y�� ���˖u+�3��R��Q��.��r�$3Q|E	mǈ�?\����i��Ӫ�M�|B1M;��W���Xo����y��n�ȑ��%���52�F0"+.�)>�l���$S�{Nw#:�@������p�c��G?���N�{Hb�B�P�~�j`����U
6��Ж�:Q�J �"�Z\��"�'���?��dE����1������BST��	aLӼ����Ӿ��`"����;�|@R��t��`({���Qȝ�~=�@�~�u�ߔ��9��|��wG�}��i���S���!�i19�>d(Z�&�">�ղ:٣5�{Q9~�7 �	�"��T�F4+�E���b�E�&�t���1"�hʴ$�����{eV��}ap�V�u) y4��Z"�h�#�,7���X&�%���2�G����0���{�HU��.'�G�T�	9�#�s��S���><N4q�D)�ZQ�G�MRWB�:�n`�m';����C�}�+"����`���h�W��)%j�v��.�&˒0�z�0��p͇����vP�h�R���	31��
�!�Di%%����6@v.���#�`����S�0vZ���u��:j(��;��X�
�.�Ϊ�ԁbQ�_���k��Y�x+��a��~s�s�(VQ��޿"rJ׷��K�x.�ё��d��}�ͅ%����O[��R��Ш����_D5$r \�,8-��lr`���v�����Ω�dJYZv����ӑ 3��c��d
��g��H+��u9!��:0%�?-��Mo{]���.�#����3���ȋ�dz���j���b��V�P��cY��ꅩ�X�ΏjM�V�A��*5�� �ɧ���u��h�@�	��|�r�c�t���Ґ��W3Z��]���5g�1��9��QQ�>���I��5��������.�� q,�n҅�Κ�(��¡N"Em��i���؈��Vq�������Qk�m|�cܵl+)�)�����n��	��f16O�a���;����Z���a��7�L.�ƍ�y..��Y��`�"�����n��f�H�p���ۋb%7 ,�g��}ԭ ���*#�%��`J���O"�%:WF$��N�V*M�{�l�[�}�p�����@q��i�!~4�
�b�M�(,h��rH�"{��{�OS,� I9�;ǿ�o�j���`6T���`�
c����&�G�G�n��Aw�Zј����v@d@{���B #�W�B��[\F+)=;��x*��$�+0���p,�-E�#D���C_��q����/$Z��UL�@۬{(/����T:=/�vJ].� 6��ф��g�KPy���+̋P+�B>���"R�qц������4������y��2�Ȃ/s.�0<�kP���ƧJ� q�����ň݀���ll>6�}L&Pf���GE�� |�a���T������E.����{�"��]jMˮGX������C��EۿE���y��7��6�e/	۸�T����s'X�7F��{�֏��I2ƕr�j���u:��u~8�g�������{�`J2-�a�Z����ǐf��wg����	�0�HXHH�P���_�I���MK!�������a�����`��~Q��YX�.l�_�>�l�=�*�������ن��,@�<։E~������+�O�����΀e�4�@T�H�Dq�A��!���lܜ+�(�"�z�p�|��%�;� kt��V�!�J`Gf��l�Dx�)�c��lz�B�����Z;��w�%l#Ӂ"ͻj��� ?l��00 �@/J~܅�� [��[8�v!#�#j���'�8V��ZXL�������i����{�M<�F���F�؋r������dnX�N7�I�,?�aB¦�IPp]6呺�O�Q�����S02*�0����M�Q>Xa~���u�o̶�[���G�>�M���A\O�ddW�.�ӵ��߫�z�'>Θ8�&uIP_&L6�_��a��*#j��(Qa+X�R�p�-���R@6Q57bM��Q,� ���F������iV��U��>o0����,�p�5%�®��FEj��t�;.�4���,<��{)�������k�4�{���=������G����-�?b$����F E>iI�T��1�""}=������]R�R�&�^�?_��$6j�cZ&а�J'�T`��^bNӍy�3mc��VӰ����rX~	�2"�1��Fqh�:�$�/��b��?O�� �i<mG!��+5則%*1�[3��ѡ6���ю;9�C�������	8)��<)��{y���L���3���)�����'no$b���I�KV�
ބ�H����^O���2X�mw�>��s{˟�c`�AэIy�B}�܆۶�c���.��p�p��8Zd��G3��R���qHN!{�3�-�����B�� �h��~��4^�����?�5% ��륌�yxk�t�5lȠ��.}(��%\����Pwy��8�4�����F$���Ȟh���S]�E#E��E��P*�&����a	J1��͎s��L2Mǎ) �����*/'�`�
#�:�B��;�~�X	 �}��2�L���/�,�(�*Iď����@t σӦ��?-��M��[ᔂ�*,�\�6�◫�Y�DNo� �������t-�4��P�T��5hm�\��m��hE'�E{��Ys�lE0�,��SHm��S�Q��R5Ph���Q���.7�t����A���E5s�Y�u�Κ}�dN"q����6�;e.��/(���|��l�s� �^�������w=���n�y����j�'^��&6}���A�04I*�����NhRg�g�X�~Lj|��΂1�ڼ.�g��H�(�M��ey�Pd��'������Rp,s�U#
E�ꔧ"���kQ"�.Y.�Εl7[u��ު�ٻu��lp�N�KEs/�g̥1VK�FR�����q�uL�?��,�l<�O ��s��6Ut�$�Q�Xpj����K�/P�)�?#�E�u�"�@B�i?��Bր]I 6ːr���{��g�e�����o��ViL�![��.��}Y�U�^���h�����{���~��,�"�%!�����Y����nt�����C&�/d�KO��O�c���lB�^y��Q���s��7��Y���4��-j�����t��H�&��W,���6��4�2�iɉ9
��ܭ	���}�]Ȧ�^���6w�������h���p�����Nɠr���Rf��0�׮�nЍA^w��SW��v䎉N<EX���_Y{�>�����rlK�9�½5����r՗�%���2�������*���(������	��Ez�N%8t�L�8'��x����"���"�uT=��J�������H��{�T0����9u�C�	�lm�˿|���&a��;�܍�~�nwj�ź%������Eɶ��} ��}�����:�mkl��*�$�݁֡����'=w�6�(47�}W�Y���<�����R���%e��luxO+��
���T?�K�a�/-HSoI�g(i�R�h�A5J/���(z�T`L���ٍ�Y���+P/�ӊ]�Og=����>1�uW�8����.�厡�i�c'f��"����d=�_���1!iqF]puc[��yj���&�R�b=�;k�Ph����d����c�p�[͸(�ln�;$~��#JY�+9j�RM�?ف�9"컹^�K�Y#V.qmD�����r�[�fj�X�dϚ�$V��n��[�y�E�:��.��ݓ��=����i�����R�.YM�B�����؞�:���үi,ng3C�8�Nʗ� q#��":!���l���2�ɗe=�k�Q��;zM���g�ʾH�8�pX���%����>���ށ�]���YF@����Qɂc%;܄Ĭ�t���=�mP5� 8֐�n�� �aȞ�'�W�!@�ߠ%���� -'��ь��DMap�<�=��3����� �������3�~]7Vȃ|F��ab	xj��M����5N����f2pqb�ƪ�F9vE�'�F����}��knr�s���=��H�:����W�&|*E�3ҠRe� ئ��w�X/���ndz�)ISz\' *<��x�A�����o7��Ư�!1ނ+�D��P��ɟ�Y��2�!��-�D�m�B̊TA]�V���8r�A��(��V�h7hl��j�x�QG���.6�V(lR�)�+Ɣl�"B2R�:����}��&ȸ��[�%�c�9]���ׅŦ�Hk�{����î-�(S�g�DNr��3z�F�Ma ��k�6�b�al}4��f[=��d��� �}ܥj�YpL�X	�>M�:��)�s���-�)��cuꄔ�����v�c�+��'�mM�}Z	�A;j��휶(��[���?��Kv�t��\�9��i�A��V��o�W��l��S۸��~qx�s"��! ���9E\�U������j�`aJ���ӮB|�e��_���s�Ǌj�{�h��#��kR@���q ��C�U΁����O'Y���+c�HWسٖ�Ŏ���#b�ϥ1�65J �u�Z+C,��zZ���&�?j�lb��6�_��A���v�U���FT��`�<��V�	Qc�8��T�H6��=Ȫ_�nnB�a�%�Q��47O���9���s���*���bm�����/8��'%q��!��_�W�;��9Is�|O�#����v��4��U8=�#�m����#�2��#�\|�D�����g�1N/�~���޳%� 4瑡��Nј~�G��
(Wc��������'.o`��X�g,�"�BO����P3-�%�꟫����A^T�=V���y<ul��J�$D���h*�����S�Z	q٦bh��B��a&�F��Up�yf˞�ę��ٔyW��"�Ǐo���]�/��!<𔄵��6v�;����[k�,�,O'�v��D	�UƵq��ɚ��jJ.�K& qm�LN���bM=|/�N:�;L�=�|��~� ���&���b�p�V}���6�:4��rí׈��D�s;��T/?��p�L��n��h�����P�vrH6_�y��R�\��.�����G-4cٕ�����,��gL֦�FT��E9����F�;{~�J��hr� ��%x��m�>4���;�-K�=`�o���3�ছ��3}W��y>R�.��WzE g�G�\�*���3��"����������	�Go }�f3|�3���]�z�;�D�C
�
uL��n��t�hoI�Y�z�#��يX� `w|"T��b�c�6�DI*�μ����O�S����vТ��Y�q2�(��٥���Tcz��Z�M�p|8/V���!V�/я�@Bl�g
�*�-^�ٝH��*�=����/�f
�.�}��}���`F��U����p��_�K� K���n��_?��r����� �p�i'�E���Xz;� 
���x���Y&�IC�p�����,�~����+o�
-:�\̶�9�j�� �o,���^�r��ɫ>��\���0Oi����S%��X:�"�5��|��v�7a-/C� �aJ�YчV� ��8��'�lE$�ub��\��3�B�,c ����j���	�ع<�H�iH���C��
ڼ
 ���^P��r,7V��ٖ�[�D\T�0��v�n�ppRM@Gw��$)b(��`�%�a��:E�	��_*�7��֊<�C5W���c��s��(�NB�ĉ�Wq�i�����ٴ6Q�zE�ѓ�l���o���#�PO%�A�\N�_�������4��P/8�q�\��0�CZ���1T�5�zO��a���$$�p{P�t�|J�X�QfYu(����-�Z��_Jb�k-�J6��'ޣ\�����ů�"�E/s��oP����?p'$f�`�_M|P��ij5Y9$���!�/�=��6r=YkH���x�2�t�A��ȹr'�G����l��Y/�G:NGu"�s=_pf�#Z�LTb��b�3@���w��,���z�����i@g��+$�1���YZ�8N����ݭ�e����ѳ�ER�%�{�t��3�.�F����EpjQ�I=`�et�jݏ��/C"b�Ő�WQXx��r�6�@�¸ff<x��D$�W.1R5Vn[�6k�0�f~5��<���+����0�%�0�&qK�9���:}���ԧ�K�����U1�����ѕˍ������?�Hl$4`�&��Ӱ��22̰l�h�T4��`*p.éu���\����� �T�@F
�j�4hG�#\D���9�����z�J�X�gZ1TDy���T_4�P�D ��oX�m��׆K��a|
	�0�N|��V2��V9a�,S�.3 �o�#�.����sΞ.*����|q�3Ls��)q�\�d	ϟ�xy�?l#���C/A&��zt�x|>�>�B쒆�7��q�a����R�KQ��\L,�/)�M���`�&��dJ�c�������ж��Jy��8����;���Y]������ۇ:Y�0q�^&*yYjR�4��M�2��?�a`k!�av�\?����6>^��~���l��o�a��a�ِ9�O�4��߉��SD�ؙ��p]l!`5?��U �R����H��o��IC�k�I�''8*_cY�h��~����5�>��@������_�K硱����bJ �9$��}���K��O�E7YŪ�!�����f���+������ Q3��_BM�q_Bd�D����'��:a�<�s>�@i6�t�$G�kL�fSN
�� �⑕��6>�Z�}|ׁ���3os#�	Eo�Ť)�z�}#��e��Ң��dL{׬�'G7HG�m�yN5��t�=�|Jv�tצrV�F�g3�wS�[��I��G�r�V&GT�iu��M�b�1�Kd8%�'��%��4��8u� ߗ����L|�3�]Mq��dG����5��������mO"���]�l��@�t����LE宮_�[���I+uH*�p�{`uQ�m֠w�YK�b�Hb
�� �L̯�9ʤa�4i�(������k�[(ߙ�Rٴ0�x� H\�֨Mt�j��Y0�8�����!�9p9���u7����{� ����Ό4/.��b�3�/�"ݯ@��T~_� ��m;�n��j/�qс�=[gF�y����Tq�����m� ��T0�פ��cr(?\�˺�t"�	����g!N�ɉN���>E4�O�=�����] k�6s��lwT��uX��i�(�٘5�Ԡ��5�%��L��_ԧ�-��)���Qc��s��,#�Z�[�_�F���錤ޥ��W�s�G1�Dr���)�ߔD�0~�I���<�gXc?
0]Է�����fOn	0�'Ǆ�S�9-�6��]�����&8��b-,	��޷���'1�Za�}��J�<h[I�����}�s1�;�3�Ⳗn���>� �p�tzWwO_���3�+�	ێ���'694$8�+-]8�H#����P �v�\wV�]�sZ3W�e\J�L��y䠷f��|2�P��w��*~gV���"��5�al�m�����^Ӄ�T�`���c^~ձ@��g�ߜ��ic��?�Ǆ(J��Y���n<^�r f��(|nR�*5g�!u�?ԭ�3����o#p�\}�5�P�����I|}�P�R�7���{)�M`�b�v�:/}�8#���
�H��S�7��59������	��O���[�5'D��G�Z�kոk�U�9���BB��B�WI��8���`�-�SD8� >�rp�~�~�J���F8��cطd�X6w*��k�����{��XcH��7>C�<���ADw�6>x���`YW	�>��Ȅ��nu ?a�1�|]�k�}3ӎ�^���g�U�%�;a�ج!�T5"T̉�}{�f��l��AҥP*ʦ=0��6�^�G��9Ύ�*DoD�Y��T�O�S�y�x����z�xM�SBm��9[)~(DA�BE0T���R�P��ANӋ��h3R��\�i��|�r:�p�c[��0�(�$����f,m`�XN �U�<�H-K�I�t�*�O�S�v��s�`�̐�o���w
��(h�|�k��S�:=n�+q �L6**I��6���d�8͍��k�({�f�:9,}�3��L���X[��oh�u�����0��'���j�l��ٸCo�k��j�����vնwl���x��w�O���0��t�Ի�FA�����(���-�9��'��WE#�~=�����B�e�C��Ƃ׼H�{	��ϻ\����K���=�N�ϼ+��,$���f�(��0?i�D���c������gb�.?Aa .�3"BE� �������Bi{u�&,P��L�~NO�U`�,�����ӥ2ʉ&�l.d����qf�!��R�l2-r�a�:�-���a�Ѐ�	&�,%�)��w�X���8N�3P��V�3�5��X�.��@G����� �,�`�0��H+��U�
�~p�쩟���9�8����+�S�i���<�T�c��r�'��ķ=�������� ��cıG`�;!|ц�<9���_")?Ǿ��!n�,�?͛GG>¾����2գ������apS`�n	��3Ow���٩ǖ_aakJO#�\�L%;��������gp睬�I�@���4��*_��+H����q=t�:�PɉD3b��b�ճ��/	Ȝ��:j�rp��	��0���殀�|'�0��OddV��1=�zG��Wg��E�Ehq�.��rRCk�F��C,~oz �lۿa-�	���1z�͓�r�8}	�3&x�4&�H֭�Yh��.	<H�64�!��)���`X��{��N��������u���b]��;9��6 ☻���JJ�p���d�ώ=�N�d�d(^�So��`���g�Ƈ�������Dx�;��1�"����[q�w��+ѱjYG5)6K�~~�5`�>�w4ԛs��π�ydg��d�-��ĸ��%^�I��'(����E�%��S!b�$�����Q�4��we�Hv��j�!�y�`Y�0{=�׷{����_U�תI�hX��W�9�!z��6������O3�����LDHAs#��EG��٫]P�8ˢ1���f��_}�PI�6`�'�/X���MZ^��0GV��;_�\̃�t�����Z)ň��`|��F]�&�]��<_Lw�\ zT���3̎I�PS���W4��d�#��.G��@(S����6I��UG-��O����?H��%Z~���]K��d�w�Z���+����۲Y���(4@>(#�zy���~�\��J�����b�P�RDx*"��)#��^��J�*wl(t���EZ6.v�(
'�c���P5�|�L(p���y5'Ub��5�K|��>0l��q���uX[bv�� �~�9[�e����{2~/ �u&g�!�`��&w�s�W�L,QᾤAK�!Xg~��'�Z��t���-]3Ε%L<{���"Ō�ISJT�`� �Bp�\g�P ���v����Uɻ��T��z��[�[���s�R��'�� /-Tn��ݏ��=�n^�ɖL���Ҟ�(����r���	cѭ���h
E6��Ga$�ؗHyBa��~��}� ՟O
u0!ۺ��`����4�:�]���u��X�Z�%�~�MO��#���m���vr�>7���/�}|웽��ɮ(��;72Q�.�҂ �&S5�vL�?�8�;�Z���#�$55e�_�Gw�܍�M�s�w zR𙼂���o�䧾�<��e�ƾB�E;��F�*y���sD&�ݝ����Tuc櫌�`�~DT�j�zf����\�v)�O���~�M�������C2��|?��K/{����dZ�?>�/ ���ꌸYj��A�p|�3�ڊ�엎�
ޝ��Z�zN���.��KUxUۦP��vK_�T�������fK��GEcC���
�+
��{���8U�)��Q�񚄛�ų�#Q�wf;]�gpB�*q��ҟ�.U_�M�˶6� �1	� s��m�,Z* ��HE��E}В���/��?�́���
`2Q�u֤�je�( m�E����L�*�	̺����ì�8�xb�+�n�LD��_��H1����6���m�Һi2��0��P J*8kw|6?��X�5��+�0�Y�q��I%���q�BƥD�����t��w\�7�!�e�/b��c��/lE��jQ|� E@�i �x�t��J��h��i�5�N|�ֳ�����i�=tL����-M��EςWH��n��)��ĭ���RNOʒ�,'�2h��{��%���Ɔ���)��v��.���QU��7�/��o��&=���h��p|�B��eԐ4I]�]�H��*��+��%���~ ��zy^0T����K��0.:R\
'�&l����ݖ�&�~���fH��M�ޮ�rb�L��qv����.@z��mx.|�$�T�]�yfU�HX3�
�qF��VO�զ<��9�D$d��oN]���ԕi:���n�|�g��|���3���m+N,����N�X�L�>���u<5����������Z��x��H~|v�\4�fqm)���b�Bi	Yt:	�����Gr_�y㓩��:}�"aЄ�A��	�VX�y@�ȫ�� �l��x�r�v��[��{��d=�d$���2�[pbrl��kW�y���j9�'+J�`����1&�� ��V!ڃR�+vT�x��jƕE���Jy���=@o�O1��b�ŶK�S\mHb�r�h�L˥��.�X��¥T�S�)��P�z�qza��#�%�G���A�fO:J���!��
���X%&�76Us/���Ŝ�(�C�5��Ȱ{�j��r���bO9�wD2fS����]df�c'��쓉*��Ø������~�X��l8>Gfc0׀���R���Z��������\G�$~5���WJ�AvZ���ϒ\��R5A:~NRXUO�g^��Þl˛�f�޺s������
[8�_n�3'�+�k@��闒��pz��
oa��Ǐ+��q~��R����F�����g��!�a�s�\����8����{��F�݉���@��^��o�p5 ��""��Z���.[�=9��zC1
� h��W��Ǿ{�
Mi�>(I��vp���M<�sJ���^p�D��_�,�Rs�m�X?�+�"���Z�$�»gw�%��V	Frk�j�v�{�������ˌ�����o�\��v�ʮF�q�㬂L�����۹��O�\o�z���,�㍰�h���wڏWiQ����M<sB���n�G�M�
�j��A�"O��fQ��e�����ƶ�  ?���9_i����mXh�Q�`�B�=��Ók\͎ k�Ô�$>q���	m���:��8ך_�y�\"���@���G�l�%�\�0n�QՌz�n��Z��Y�I��� �Kp�P �����,1���ݞ2�>�|��-�Ώ���la�J���\��\�0]�F�i �t��#!�L�[��ƥ`㩶����j�桼�\��N�d�����,�$�Čq�[���s��(2�Է�MZ���c�p�,���y>�\[=��`d@�7�3�H���Gd_F����
�����
���G�k��Ĥe��Ή!)��[-���O¢�2�̒����^g��ml�U(b��p���5KP�jbK���!��������œ*ķE
�٬r咍;�MQ��	X{8�h���W��Z�{���j������>��W�2@���K������3qq�G�x�>�L���R��@�2�ǔ`+�'��LPP֔�oj�O�4bOMPH��R��@q����\,��v��hy9m��6�b��jߠ����N|b:Ӭ�b����\0��"�x��u5۶�����Zfq�)�^@0�~�#���g�����jX��$�Kn�	6�F�v��L�L�tðNe����z,�����@H`�������"EA.6���/���g0x@��7���}>�ɯ0�nD�R�q%E,�vS`��K�T
��PBb��Y��y$(]�Y�+��+�h�^m��e�����Pp8;���at������SU�+�Jc��-C���zI�ո.�'�O��s�aAZ:�m?�2S�2[��C�h?d:�o1<�旇#��6�؉�E΃V���G, �|�UR��ԝ{�ڀ������K�y�H��"�&��O�C��$�jU�9e���u����t;�O�c��d�V��_gZ��t~P'2�Ɠ:R��q�IU�d/�S���$,��=�W�\��-����9_����3��2E��V�V
�@��"a.	0�$�4���kf�蟩��;�����6�|�۩���ە���r,�}YY�Ʊ`<or�[nH`�9���1M�np�֜:]#*d䜁~�4˦!T[���)8~͑If���^T؆@y=��h؞��z�O�!��CΖu���ŷyتd�X]�n�Gx�TW)��9�#��7��)�� ���G
�:5 <&f��� w,0]�����𡵡��f�R���q�T���2�rTN:���g�@٠�E}D1I���=��yY�j6�!���E��
[V�Å�|�o���&ny���0u��e�0!���� �n�8�-u�R�8�F>�����P,�w>�{��XD��~Z�Cwy���	��^k6�Մ�=�W�d�Ab�����z6���*s�i u|�~�',�_ި����˟Hl�G�m�d�v(���H��'��K�����1(��kۼQ/�-�/+H{d�N#bWC�Ǽ�5���}f�ˌ���Zw���;r���"�)��&�쳣�X���ϡ)�u����>�Yr��a�z�`�G���^���(O�2�8A��^�V3k^m�r��ֲ5��68.H��}9���u莴���,�R+ƻ(�'�+ׅ��Ƴ���x�$)8�H�����/�7|~gTc�����҂���x��ác[B�Ցƨ��B��-V�]��xڿ9�Mz��,�-QUxϱ�m������[��:?s���e�����b=��g����7��5��Fl/�l��BE\�z��{�)�؝�(H�U��y�-T��g�⮞=9���j�i����N�gϧ�M��*
��̚�<$���-(�ȇ��V���3���{��QH�403%�;E_ȇ��$�$�;T���Β�n�@��w	`Y�As�oYw�ݙ!e@3~��<�8�Xr֌jObvE9�a}�WI��,h,[d��"����#9/ϙ�����X���qB\�ؽ�
4.܄:�mϷҶ��-2��4b���S'*��*J��::u������"㷵�?J���>�5�2����	�~)P^�<�5�J=ɿ�e#�!����l�çyG��,l���/� ������f�lЍ%cN��s�5g��7A��ٕ�fX6P҆ނ��2J<)M'P�Y^Dޜ�)�M����pWS����N� ����� ��n�Mrwa�d�.�������5�Y0�1&���$���)n~
W���Q�\��@&j	�ruU�\��w��{���R���X��oD���A�O�����h~(%[�DԷ����lX#Ԋa��ܙ�zt�Se�v]n���4�Ul�)CC������'�4��,v�4 �&�����V~���B����[�<��"<�=Yv�$e�-� <I��2X�X��������)�0�����Qw�!\�wSc�n��'�xwt���Dr,2aL��3@}rC6>��� }}�q���&"%u�'t���ɗ������c�:\�@5����ܓ�4�!�g�}$l��ua�m@.V�}׮�\�ZIj����hH ���!E4��w���a9���jW��vm��͵)Z&�ަRi��,�-�LHy��]�A�Ce�W����� �~ʍl�D3zS��(P�����a<�X4 ��VaN�|h� _��g�a$��n]r���T�����[n5w(�3AZN��ދ:oR���s{�",���"���b7�ɚ��\ӱ��=�'-������GF��%o���-���#	��5��=,�]��Rp��g ��Y���տ�64�����[��g�F�����"q�h��L���әv��?$d9H����S����n��JG� ]O0�c�n�m���3���R�SA�R���[�v�<q�7o��pE�@C���5�L;����g)6ٞ������Ȉ�t<���s�>��Ws��ŗ԰��Jg��cj���Sj��E;��^��I��*�I�ɆBR�^�G��=�5�c]ʢ�\l��Na��'�F��p�o��\�\X�f��Sv�cE j����)���羒�Z�(G�g���Xb�Vu�����0�4�Z~I"(d�u�C�*�B 2}�9�4B۬X��Ē������?���G����르�.�Md��J��0a�}"RW�x+}ZٶL���Ѿ?�n�<HR�<u�c���.�t��5b��;v,������>ӵ�ɍb��ͅ�T&�<��0O�!(�C;
���c �+��;��S~]���-*~)u�=�^+������q��}���S|�����N�0}{�ɓ�&�ZDG��@+�g%<����'�|"R��^��b���ھ�������-1��V�Z�d�~�<m�{�%�(���aY�4����Z�m*Y�/�A.g3�|��*H~lz���q��-���ͱ����l��&-;_�"�-$P5I��H5�N"+E[?y�Ӓ3Q���O��f򩌡7�ɜA9��� S�^�"B:��t�	�r�Wg��nު�O�$�fR�&wHp�3��s'��4�ν���7�0��ARLc���p*x�aWT�F��G�u�#`6/�K���z��3�Т���N�M<�ە�$��[�:[ϫ����,�xYy��B<J��=Ё�� �b�tX��G�1�'�m�_���P��~r��mo�ҧ#�;�i7Ml�9�� ����
{H�ʱ�p���Y{��b�;�p��7>�{4e�Qp�p�|�q�>��N\<�laV��7���]<�8siA�0j�}�
}�&�1�ʙ���ˏfI��fCq���<���|r����fZ�m�x��&���@����2�!QD���:�D�z��ϩ��bE����3�I6��^��$���_�� &s�Uy��B��;f�����^�@*����;��F.6�{l�֎���D���|C��i�c��/z!���a�vq>�M�4&}��!=�x��:z���!C�9�r�q۾�*�P�D]��n|�97���3�&bw������;���f; 4�c)Ӫ@��.s���˷�Y��b�3�ͽ
y��2e�����̺B�6�i�����?��!�Q���I�P $��wˈ��ҶL �H``A�^_�ҡ}����-���&'�S�ZG��O�s���j�,|�O���e1K!]�)��6�(�^�ͫ�ژ�	����'.���%���?�1��Q�\����9��_`�cwC�&��S͡�y�M����pk5�o�0P��*�o�R�|�"�"����f��x���E�c��j���Q3]�
_[���U��q������G:|aG��\k�^�1��g�������/��ezʅMa	�"�������rj��� 	�����L�Lp�n�l���LAl��<���8^eS� �a7�߳��X�Ȟ*|�u�'-�Y*���q.`�)�˒��Lxq��W������2�;{�+�����Z̸dT؇�š�������p��Y0O��Jz�V��J����r��F�&�@oXF�����J�rv������O�G7c����`�-�%����}I��d7��تW.�?Rz)r��ʪ�����#[����ga�U���:�jq~%|W�+�G#�˚K�i���B]�>��,�0ɥ{�j�$Wa����a��/=��[��`�1�Z�Bd�J�z����%$"�ab;�ɪ�u�"���Z���'���߂�R��!nLˎ�a(/A��ݪ�(ulz ND��-�]�b���F��pS��3x��2��Hj�{�d���3O�4id����*1`�{Tz	QH�;��R��Y��[ <�~�k����$���̓X�;ν����W	��GIMa?f��&6�"'�`��)�_N=�[�<�[<��El����o6��^�
�V=40�2|�` �寐WvVP0v� �F�+�QUm����e�4�h%�X)�}}��b���� K֒��(�����ҏ��`�[��5/v���~�x?��#�W�v����x4;�v`$�][�?"}����I��4Lg38n�$� �y���W��9���X��E.��rU�LWͳe��Q�,��͉�)�Q�Tl��%-����|��BY[�R��1��;Yc�ө_����F��s���ô�r�Bu�J�����P	�HE��IAc �<��j[N/�0* ��8�x�̤�jIo��=��!
����HR0O�.qozc4�D�SX��{̴݃y�"#�e���g�t��7�Á��أ�^�/��63�nabP�f8)&��Ǆ��%͉C�T.]��zdV���Lx��\�F��ɷQ=6Ю�`���eՎa���F������+N�^r_ ݭ�!	M8KT�k���vښ�$u��\�\�M�Ѽ�K�U�S�19ؿ�E�_㞾��f�)���S�G�h$���������Z�I/-ut:�{o�i	����\<��J�?��+x��i��
�Zig��O�E�W��X���˟�+f�2���-I:&W5R#d�{F=9yڰY>�����v�g��ϣB�%cx��\[<Hy彎`zh���$Ep�O��XSu�h'�U@�a�Ձ*o�7��i����.@�W.v�Z�La��Rq��d����
$�B�O�M�:+��F���Jsss ��!m��1��hj#��N��lU�{�\�X��S�}p�Xs����W�l���|�܃��1*�:�g�L�"�k
��;�/fF}A�������Vo��)�Ww��z��1$�,�_�(����^��~P��2��j��5����ԮndbB���/�n�K�1��7/wqt�k0�����L\��ܮW6�WY|�5O�6�n�����ϸ���p�@Dt��O@A�˴PQ�p�'h�#�,�Q�Δ����ǭM<�s����/�����%�IGI��y���mNa�0в9	K�s��f]B�(}L3.Y3�$���Ǽ����!��RZ�9����6�9ۆ
��d�P��.=��L��}��Um��\��h�X�*|��紛݊�n+b�S����1�Ʃ�4�����HNrߒ�on�Qb��$uၲp�\�0�}����䞀C3�)-����n��xo�7H�1Kp�'Y�O'��m��ٞ�S���-�q�J�G7��!(Ō*��/LK�ݡ����f�
�a���(��z�q#kꈂ����l���}<����nF_�r"�9�͠YAƛ�hDבq��tˎf��7	��*������E:����8�bqk�%��D^�D�����{y�ֺ��o�DJ
���G�Mw2(����Tj�;�:��O�]=����<�H3ӭ?��N͐`�d��JVI~t&����g�ʢ/�h';��c���_����m]�H�|��m(�,�.��^8�gq�1]���s�x��P�XZG�� ����-��(�d�VP|�y�F-��Z���G��2�z�ߪZ���jE��{�:5Y�XA�L<j!�GC���"w�b�@g��=�KE!XR vK�$����� v�&�^O��v��������Xjy>]5e������K�Gҕ�w���a���
>�OP�ik1��!-�b��p�&��Cˈ�Ɉ�aa� ���Z�#*�Å�r��8��6ά�5b��܆�~&��'��J��1�$b�%Y^�n�;v;M{�v(��<��Л&��\�B��0���ǆ �'(�%N�2o��i�K;�����B���`[��j��{��+E\�O�a���S0��W��p�ҏ��l���;�-���v��̔����b��ц��Q�j�M�|�7Ja"_X��|6Y��T!@=���mo�c�X��:\1m6Y�;��0�rb\f�Q�=x�n"�L?Ne~MՐ���� �kC�r��r<'TS�"=~�UΉE�����n�3ܗ۞G[tp��jÀ�x��GZ���c���|�}�`[�@ح���1�u镁U]2�69�v�'��E���!�f���lؔt�	�oN��=�1詀�� (=�S`�H���[b��↺�R*x�q�Ʋ�Ύ���A�E�R;T6�����&-��Em`$�Y��~��6�[��6R�8�N#��`ef�5�R���%�Xc��rfb��q����ƴ���4��)E����$~�o��]q�|��w�fU�D�φ}~��Tν'�'�?}�zb�	C]wi]j=����F�N��
�A?@쐲Cy�yK�k�09�y0ǳ-ۼ2�xK����1;{�J|r�=�� #`5炯�'�[�%X���qI
��ʁ/�r���XA��?}�ᒣ�&>:
�ޛ�d�֨�_���I��)�a�Ne� �IL��z��I,�m�'�,�g�`�K-�ܿv@��素"������k'41�lz.�G͢0V�7�����l��$�$PN�\�w�XS�����)��e���囹�2�����D��<��Lj��$ k����lnY�4�l�]�,V��{��+�	�3�'�١2:�N~Lp��г��%;7�h��g���R*S��,EZ|Ul/=�D|/��m4�����]�|�h���pV3�UQ�n���{܎���^�r���5������<E���&��m�e�(6�A�(K�ł��ãM���/��&�w��_�]�3���~�G��ۻW��x�)NՇZ��Xa���VR��a5��N,\�@
:� �oR���"��%6���CA궰!
�� �c����i�V̔:ib��UY��u@���w`��x%��l�]]WN,}�M����[���G����߇S��^����|���J�^���J��m�׼/��S`��:V�y�����������~�	��ç!�(.A��c�͵:�;�1bWOIj:y�O���t��+�)A"�]4d(���~D.
�������9~���L��������mݜ"����v�R��*P�ܷ��x%�����㖞�-���z�r�1����Y]�zb!�5���*z���h����G�#=�Pn���s
a�'�6�9�,{0����A�o������B��	mI-I������ڬ8>�i2���՗ �p��{�W�cq��g�g��
8~���q��1���*�aV��i���
 w��q����׍"��i87A��#���Q�)��������q)�dy���藞.}
�Yl�]ԭ��H�e9�v�cL��1)�9��)c=���w���a�ح�uP`�[�#�C���s�w*,Ǫ�v�����o�u�^��%�[B"3�L=�a�e�[M����P]jJNYپ�/.ae�x��6*`���C��y<D�f��*U��e�!b�	$"��]�ȕ����$�	��s�94
�{����E��P�A�|�eu�l�@���u��4P�{������x��޽r_�\Q�0��dg�6�ڟ8�Ӡ^��-$���P�^s�aU&�g�@�;_5�wo���'.|M숣X����+�B�UV��Nh��Q��R*إ�d�Y�;��	�w%��>6���P���t�r.t���`���w��@-�A;�?)4��KR���}�W�⪉2z���77 �@E��x٫���\�F�NX�O>P�urI�@7G��P��z~倦��:+��(�bz:~��-�b�a�:�7��R���yz����\n/��ʸV�9$z1���D���$��K��纶�Z%����n�(F�L��sx��`��0�DԱ?saٿ�8�؋�"n�",.��]I��~Apn�bR��YV�<F+�<s���sM�C��֣#�Lhf2Jc��<)��k���4�LC]W��+�c����d�g��Ph��?�Ѫ���d����%��L�����>j
�(���0�4���^UrnPڅ*6�M�։㷝K8�,� M�<�3���E�o�z���b����dx:AG�G�����E�H��q�
]����m�?Ϩ��H�,�ς��sp8�U�*��܎P[v�|��r)��HU�x�T�3��l"��';���@k��9�,�O���3�<�O�	#����U'�[�2�o��V��u ��z�A��!�b�8^���1Qo��HJ�~�i�a�ß��*Q��D����>-�?c� `uk�۩��/��VW�Q<>/�e�0��~�j�C���4�*��B"*z�W-�,b�u�0�$ /h#�I�/z}Ma