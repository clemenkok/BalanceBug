��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�!��
��%Y l�׾�Ē{�1+>o�^�\{6CT�����h#/Y�a#�:R�m�n�W��wf~@�ʒ~��w�H����S���Q��;?<�m^�Xy�6,��\g���DJ�+�y��3��&u@.�Ҽ��?F
r�2��#�s?�|6Bʃt!7�0��^h�O���%��-dޟ�hB]8���֛���GD�?�6U�$�?�A����{h�Q������D��X�آ�	�T�H���C��K�H�a�=slE�Qp����Ѷh�쉌>�w]�
�8���-�o��$`W�d8�
W-�\�x��[>��j�i���I��c�#��UT<Im"�/��L�`'n̅�)��$�S��.ǎE��Q=�ź���D��+�z��P�9h��
�Pw������VX���z�Hg+���H|�'�8���=m��ë{��]C��O]%Cn��|�9e��7�Y���j�0oo�봳t�N�o��$�P��'�l�M{(����}W���[^ik{�` i�0F�z�M
�x�����S�����s5�SeLvn7�_{Я��EdiksEٌ�Y�P0����I�7##b�ܪ�<~��Y��w����2#A�>��*�ӷ�
����� �,f�����WZ��Tבv�6"ǶȖn+`��Z0����,��)�=-S��y ������W�Ar�ܸ�B
	M7B.)6?�O�]q�o�ޅ�*�HI��VŖ\����goM=�{I�n��C�q�⛯�W8��R0���:$�6�s��8��zJgB5j_��=�fg�_gI_)����i,l���^Hcs��E2�W��/ʒI�.�X4���\c�>�?��$(_-S��L>Sj��7^�W.�.Vo�=�w�M+x��i�0É�3O�y���� S�ln0Ua��)L�v��J��V��Wx��S�}�>�	#���9�;�'+g��i=G���w�]oY�QK�MV�^�La�}W<�%��1r/��8<���7^�E�Q��ꗛE.	���J:6��9�A"�o��1{�Ɣ�?w��h���T��Q8-�q�� �;)��˯��	k��� ��eU�f����.9Y渼�����J��Ƣ�z3ǅ��sÇUpd�D�AVm^t����x��9����?#������d����3{��9��4j:�����r��!�f�/	5�6
:wE� ���}���ID2�s�܍uu�!��J�g��	ft�GxE�h��a.�-�qVe.��[��%nBrfi:���+�˟3/��e�}i���7� x���^�Op���>H�I���u��]��Ҽ�r�8"j=���u��C��j�:*U��BF�]��@���Kr����c�æ�ת�K[)�:��E��d$���Ie�T�����lݱxR̠���-�U��-`�k��;$��|��$�<g���������}n1�q[�:�5��F8mY������ں�[vv80Z�r\M�\��;�^5�/��;�l�S'�vwF�h�<���Ȗ^��m��-c�Vu.$��!ݤZn.8|w��П�c6Y�����{��OFk_���A�\H*v\���U���޾ⵡK�m�S&M�df4k<��b�Y�XaPW�����}aG5<c)���˦P��}	��量�G��7B5��C٘��~`��Sd|�[`��FG�
SZ�i!�{�Idd�?���[�'�"�H���+9��w��-/7���X����)QBR�T�y<d�dZŜ�r����O�O˵zC��74�=�|�M�:�8�$�f�-�Z����!�Z0��n������P\��su{*���ᷫg6�e�o��,d��9ןV{c�4�ΐ��+������6�;�?c��á�4�ܺ=���x|�~�-lN����K w޵pPB1K�XH��v�-?d�Va5Y9US©��˞�.�z$�{�)Bl���lj��+-J'�g�|K�[V����րd�b�;��C�%[>�!�����mbW�U4׏6����?��<�@2kI/]8M= �<cR�Hĸ@��g>r�f�o�80�D��g���ֿ��j�S��;�����H��&����Hc��&�2������.Hė��CoդL��y��}\��L,�OG}�*#�`�[�k_f(�y^�K�<$�)k��>������{s��Կ��mn���8�l��I�	_B���R:Il|(&!��o�>�Y����)�Xtoo�X:���3��gãL��Pn�Kܒb�����Q����/���wK,��E����#4vǌ�D?���y=��qΤkN����kڨ�R��I@y��~ \�u�P�!���@���]��sw��O�߁�?�*���w.\}��aL�Ûc�����^}��<|G�V��Mq-�U�m]3��( �����5/��=!B� 'mjS��e�]ŀD��s���T�Ll������^|�o4��
��M��,;ÐCF����.�)�x҆s3���$ ����z/��O���Q�?��d�!'"���	��R�OT�j`�وg�xu2�x8Em:j�~�K���t�+�C��{��9xI�t���$;,�P���j�&����yD`���J��Iuge���Ҵ]t��_�r}F��!5����b���ũ�+=��*�ױ�_�%t��"^jӦ�j4�%���2X�'���隭Ӕ��u��tǬ��7�8�,L�'�vin���wlS�=�f���3��*y����paPr\k�{SV�A��"Q��V���t��Ƞ��b$RM��5�m���+t���{@���@Ct���*ʤ�@���������h� L�v�C�z����������̂F~�m�Y�H�5��s-�	`�1iAA5t����u¹s��7�`V��m��"��Jy.���o�9�4t�c��ʴ窫bW[�Ԁwc�x$�I��āS��,�w#���-�a<�f-�u"� ��D�eDdD�_ƺ^L�`,x�:A����o���d�˷�e!W��ބߨ��0���ɟ�_I�0�Px
�pm�UU�B�-����`x�z�o<z�w����a��� �>�֩���XY��&�ȅ%_��\�E�9�P�n����7�����������{cЊ���V �I J��̞=���Mz����sEU���з�V�%��͠���k�XFx�X��M,�f�f�.� �&��o���$��y��?��ogp+O�v�5����Y�R�M�~�:��[)ҵv�H�e$Hi��6���HZ5rX�]s^)�a6sҦp�j�S�����l�Ҝ�GY;e=5)N>���|C���+>I�6gR-t�<n��N�%�X�n��߀H��e+J��LO�gF�D��˪�A�3^b&q�j�Zm���dN+���Ǉ�����"4C�
���숪�6�W	�u{F���bs$���1���X�~�>��-ȧ�����Tq�9�
��)#�Tq~�}ǯ����H?Pr�����6��b���K\v���4�E�a��k�\��h3ʓqG�A��(��-��$rYyj�%�Ab����JǪ��GA ��e��8M���&{8Iů��Ox4[YP�ֶy"�'� ��k�&��\z��q��Gk����>��[L�R�HK���\��s�ҟ?��^��V+������:Yɔ��h^�ɍ˫ΰEΡ�Lb�6��w�2I�sϭ*��� �]���Z��MR%�hV|]��M�߆L�=��,T ��� �/���s�7�@U��#���;�Q7Uعm�}ч}��2��A�3�:/�2 s���ݙ�
�kb�����7v�nF��r�p|d^}�;��
�D�g�l���LT�.,���S��AQ�d�en�N������N�O���xs_QE/�淥	�Qk�}V���n�砉a�ņ�ƅ�`�V���'����E�Nkf�T����do�bcE|f��=��e���~��t�g�c���
;��.C�0Wꁸ/ո�1JI�l����Q$���y*��]2}%uT+�H@=�/�lPW�˦��K-�g��.�������	�<�M�D���������Q�ɟ�؃J���W°&�;���� �;R�P�rS��TA�d�=P�Ls���%={����-��ܕk+zF)�/3+�V=�KJL�i�Q3��?�h.�*Nu5*c�݌GU�6.���������Os���oQ7�]j�S$����{u2�c�(0�8vW��7��f��U�g"-��*�0~e"g��lY�j��[��t��kJ�V�Ϊ����%�D�=5��� p�����S�j���B���|d+�3EP�C$$�y\�QBS�&����0�'�vW���"`�8P��p�X>�:�9��pZ[�Ǭ@k4D�\�z���;����5\q��܆x����c*��r�!��ۥ�f'��5�^��7ိ�9[�sV�zAqc�~ ��DĶ���㽦�4�~����*��o�tA夁���&�uI�W��z�����ӿW	2DQ�'-�8�)��M���V�����IE��	��e(�)���4�jvmI��V�,��ke�x_��E�cc��Ԃw����VS��}�I��FC��;Uw��]c�C� ��s.P�Fj�#�� ���*�*Z@�G�%Yq�Y���<�M�����e�V�yy��rSZ s���2��ܸ�kǙ�D�e�)�*�/�.��ՎM#ک��$�]���|,��/��>��/���G�Z4�����C\>��Mޗ�O�a�w�G8cP���b86��2C�U�;2_����{����Q)����I(�2���8lQaK��ߩ�8����0!��D%���dg���'ǌ�ٱmܤ@#������kk�h�ݺ�p�@إK���S5R��Q-!��h��c�`_��
����\������&:��-�Ϫ2�g�jQ<�L�R��|V��9DԖtP�u4�9�!�-�Qw��Z�i�ܽ��$ʥ�*���[���T`�I�*�;��̽ Q�Qo�x�Z��2��V �]���h���D;�����+r��0�P���)��;�q��M~v���Q��H��[���?��yjj�!02~�-=n�S�<�@�� *�H�2�#�b��/����A�E�e�.Q8�N��`��^zSO#�Z$萍&�Fܴ���6C��,��Ǒj�x"�$M�m�l�J��_CX[���v�r2����1cC�>���mĪ�����`x��2W����uFߑDá��~j��B�"b�\���P.H���i.H���� >��B�oAŕ��uh�w6'R�f��`��w��b���� �f)5�)�|�.,� ���㒦��bD��V��Z:���@B��@��t����F�Amu���U'd]@�J�_�Sd�� �U9;�Qxo'm��޳!X[���#J'�����������J��d���+�����pF�^e�2 R��E)c�[3��n�#�	��a����^�wjQ�^��Z����j(��.�/��6ٵ��+����t��I�8����A�yfs5��._�xIK#�ebg��A��
��T"�T�������|����sXm�S�{ؕ4�ј��N�f��i�և+m����~�����k�!H�4�k�(T�}w|@!v}z��Yd�Z∌N#�uS��{�,#B ]u�P�]U� �[�Y�Y{�c��9W����X����,9o�T+9��z�w��b����ɦD�P�/�;���tNQ�fjk�r��$�߻@��鼬�}�<uz��H?2�L胡�>"Tsx/���T�V-
���Y3e8K=B��+G��8Lh���i�T^;�uV1�>a�w�Uil�\|�O �$��{t"�ڼ��P}���%<�G��cVD���r��/��]�g�r� �P�|W"��P���b�*oi��-�ٝ���{������
�s��e巷�F^F���N-�!1l��n��U\�b%�2�a�@��2��U�ߛ��8�j��G�[Z�ܕ�d�P����TuР��Wd�r*�<���X���z�����iHKǑ�GC���"���d����������ȋ,�ݼ��<9lW@�	���g�B�P�}�!�T�<ڂٷ�۫�RuW"eM��\�k����̴NeP@�Պ�M�ˤ��ƅ���#K����;����LF/AS5$@�.�0�.jq��8nQ��ʖ�E����Q:�m��z�P�}�1���z��`'��N��0pt�(FI>���S���t���	�9j^��N��*C��+��d��b' ��sN[S 朐���_g���0V}�`U�����+���W�bE'���$��(X=00��K<�܃F�$�WKk�8����ޏ�7LP%4�����T���O@���H����c��KE����I��A���.ɭ��;LٜU׋��M���Q��8�O�~��������rk�N�P�g4�Ei�)RZ1p7a�Ҕ��ĉ+�n=@;s5�_)�Oa��=�D&�a��M;_q���8��	:��a�aD�3���1|����_��r�"��BeǏj����A�p6_I�Uz����n�U9>�8^���{�����[�Z�v� d۔���YQP�+�U3`Du3>�뫠c�q��304��(�9�z�5[>և�J��סq*�����#D�+�Q�'Xu�a�]Uy-��ж4_*��uڗ�wX{�ڮ�ERW5�2�[SzZ�,J�Jbq?�R^��}���et=�*S�xWn�Y���
��Ƴ��e�zJ�`"�������rC�)��G�����1�/�����ǧ�T)�7a ����Yԝ&��(l�R�Q�.t��:vre����>*[5�f�v5�;��T�sM�zT�2Y cK �t�և�2z��ĂM���B��1Ŕ9�e�����8��l*h��!�;R����lC���GV�j$`�KR��v�]�+�gFe��A������,����#}�d����ͱo���"�t��n�F�F��D3`*��w���tĲ��Hg�U���Ն�\֫���#���`�o�p�j�A__����(_�3�� )�y��K��GG���
}�p|@��Im�Y# Z.sTs%`��oK��Ԣ5�fD�����Ux3W�4�ko�}���B�<��[p��|�OJ=m����X�TK���?��tß��'?o��$0{͘H����a���X���;K�ς<f���E�#S*'x����s�1���H��J��ۦ�ڛ��D����wӃY~��{2 q�m ��
��Lk���X�	SGEw�����։-��C�("A����2�
{J��m>	����0�� o��� ~�襼�wC�n�".��J�5f������:����i�rXgԖi�蓒Ƙ�"n��e�DU�&��+!h�@�+:��{^@(�i)��a�O�z��_�W�䧋-wW�Vg�.��ۭ���y�[K����J�U����P(�(ʽ6E���C�}'&/U����*o=m��)��ˊ~O��B]�Wz�p��?єك���v��m����I�֪�g�2y�4I��&��e�l��a4�I���.��LgH��X�^�z~��2��~�r� �]ݠ/U��^�fn�0t��W:�c�v�� 	Z�e����C�,ܶu��F�`k$�9Զ�h�Z��@�:��d����Z�U\�lp�X�M�2����_��g�O6E����ʠ�es�Wk�L%�	u�GT/���lsr�Bb��1�l:�`�
F��a�p��V��M= ��#3�V�`���[.���8�>���|�|S�J�N�ҷqO�Y�o#��ȇ���(z�+i��|�+@U�kFH��K�%���L�ߒ����I�$Gᜧ��r�S檦�!�NjUo�1e���0;<�Y��;�3H1���ylޙ�="��L��yY��U-(!�c��x��@U��09���+~OW��љ���1^�3^�c�v����:���6�e�ܯ���#�fe);B����~x�p�(�e����!��y�f`�����8"���>��0N�,0N���|���:PОp�	�l�m���͆]�h��N��F�X/�� �UK#�>)m�@�b����r�1��\� u$�ڸ�nj��hʵc��m�a���D��ǣv��ȏ{E���igҦz��W�q�>�gtL{�R��5\2�S��Ƴ��M�V�	�V{��	#������r��*6�n�و٥4��Ap2��E�$��5w2���a���0���d����y��_6�������
߶jr��͊X��2Y������� {�������2yxc�W��֝�����&+��n���l�Z���jT�{h�^27uލ$ѳ�X��ifp�\k�5/�U��ǧ�*�i�є�8h�F^����8�����v��$�ƴ��(`B�ǹE�7To����ۏg?A:����������%PC�`���������`�c5>T$�tǫ�n��ji)��(��wl4'��s��x������Ь-y��E���b�#���B_3Jo=���֭)~|	k]����c�-tq?�F�	���q
��ZJ�����Ȯ���y{�eЅ&�|j�J���[M�d����Z�~7�v��	n����G���J��G��h���FS���?c!P���҉NG�Pjd��xn먷RS t�
T��w��,ǘk�5*]��o���b�+9��6o���{:C���-��Ӱ�O�Z���+Q��b��ư&M���jo��������J�h��$�ڶ�Rº�Z����1�~I#v��?��~���;�Mm�y�U���x.#�*x�B<�wHG�ԝ���R��b����H����@�d������g4'��4f=�˞p�a����0�dbFT��1|�<�C�&�yR��Y!� `�$��4�= �,�g�s`f�@]�r�����φxb�뢹S39`4���h�-j:���`���1��K�(LsC��MQ굨f�Vb��ʣ�s�~l�X���U���V��Ҧ�X����I/����Y7I��Ӏϥ�ڡ�O�`��j/V,s�!�t��Sd�Y�G�f�Y�l�شb~�j�{ю�u(]�~B��#�۠;��Cp�Y���P�-�{u ��J�S�&;��Wϓ�A����
8�D����0fd���Oj���E�#
GzafF��/�k�%�2��"��ɥ�-�X8�i1�2}�{��3�&��.:����ʟ2��x��:��܀:��b��FҫWZ�=�����Bz���NR#Y��Òؒ<s�3+>.w1�qÕXE��Ѹ�}[:�z"w'.�JÜ0үR�+�!l�o�rx 
���}��fiS����!���j��:�1�GO��l� [��J��zA �0yF�^C�*�/اK˂=���ze��쑿������-�!���-���r�v������l��ي6�	�ǓW )�dPp���zq�M��G2Y����/�1Y�d��2aF"�7߄�3t!l�ƛ#k���~�Z��Z��	��a�*n���֖x�J���ã��$��NS硸L<���<p�79��]xӗ/[+O��br����"�n�5��"�* }��j7E��N}ê�1r��(	��C�z�+Ҭ���?ouy=hV�;;���c���P��}�l�Z�����l�+�P(6�Ν!U�-���ᖌr��[���TA*�xA2��5�4:���\agIu��l��=���ߑO>���J�%FK/�)��D�X^��1�ڀ�1{5U��ZA���^����N@���Bd��d%��rf3p�8�:(��Rګ�//?����(�x+|��Ղb�ygn�BO<�i���L��4^�f���߯�[�BN�z |x��4��8�jW�ㅇ
����u��&���P�������[�,��� �i"��҉��34�����o�L�F���(G�O�h�v$�rO`�E&�v؎j����HC�Źވm�W�>(����.'�6x��}���(���b�;�����s;�f{��I^�I�<Y��E�UA�1Lʳ�Yr��WĢ1���y�g8�ņ��-���H�����W����Xt EI�tMBƅ���f JvF��Sm#�r���G2�Z�i`�C6���4tb�B[�$wN5�'B�n~mX�,�:��"��\�s;kz�NB��N�g�[��Q��6����.F���9�j[��^)+���õN��Kq-�=���:*�+�}�i����V�~���h>���y�0�VN:.���D�H�	�7��|>�=� �-��b��`�f���9��*��Q\�����h�� �d�^�RT�JiM*�$�H��	 �T�y�-��f`�Ѯ��
Wf|P��?�����&|&v.HL�)6/Y�Z��q/Ӊ|\셇�.�Ep	�y��u����4���x,���� �K�siA�O�g�WmdFf(�;M����G}��URI�-�㋪��$I����j�ebn	�3�8���gM��pK�dF���>C�a����ÁE�$�y �]��8�\z��yu�<o�ĤG�a�T��)��JtM%S���X8���$#98�V?!�>�ȷzIn�����|Ա��tm$&�kY�X�E�R�C~iU~m��Nibc71¼@��^\h���҇(Yc�)�ck��e�����MĢ�q����9G���֯�u�z0Ӭ�G���l�;�ԑ�	��$8iP)a�;��1�m�(����*Ei�z�|+LI��>�A_�Z���:��X籎��Kx	.t��u���}]�q�IB��N�.;�������D��<=�(�v��[��1��ۍ�cwgG}~�wo�����\U[W⹃x(��z�Ȃd��"*��ʖ-&[�{��l_�`n)��C��
�GU��)1I� ���ǵ3����{-�1�?%K�n<8@*���t�y|�{�AH쳷�7�>�P��T��_�=.r���M������}c�n�d�8�/�M���e�Q�4����yŚ%��FO���-����]��� �wq92�i!��Ti�ʣ(A��S|�7��۬w��M��nV���4P�2b˛aҧ��������F��+|m=w�,.��S*���:�#"k��Α_�9TaI�{F���7���ڗ͛� fZ���g����r��q8��d-j֏��u$��oXzU��%�P������i�k�T�u��/yR�)�+���m�ң���.�f�H[�GJ��؀v�}���Q�h��FU�9U������Vr������^�3�ࠈ��P�̛��o(�PSy\sU� |�/��!����h~aDY��n�D_5� �7����q�y�N�M)	e|�q�j$Z��u���^Mu�X=Hb���<�`Ϳ'K��������a�]ʥ��T=�q����P8�,YS�M?��B�=��S��d6��mM�nIS-��nw��ӡ�����i��24L�
6WR��M��� &6�ɪ�+��e$���)�$��СzUؾ/��8��>�(^W�-g����'��q�g0��l�FV���^b�φ`�/?;ם�X(h�t�ZN5	��8��%{�;^�Z-�� ������_-'t ��U'��F��~�!��[�-��ʟ�*�����k�勡��eM|�B���i��`Õ\	������S{�l�<P|��"����̥E��B
5U���;����b��9����㉮8U�aqC�k��3�-vqI����n�z�A�-��M�G�Q_V�kV�u~���2�����iȕqn3��a��\��N*@F�G��%�-I��#'>DW�ލ���t
έ:�=�t��a���J%�3\(��M�@�`&~#Ů�,͌���ъa��
*�s�e����Ћ�
a�uu�M��D��o9پ�.���X�T�-�c�1�ӞI��K�/�G�)AO�x�T����w(<*��>��ͩ�*#߆�ui�}D�im8m�0h��	�) ��wa�;�-����KT3�eW[2���R#B������p�c̮v���+�X0A�gZ&H�o�
ƻ����_#?GȖA�'rX�n���Ip�$�?���������Wn�kKd-��tQ8�`�R�����ѫr�pL���o	L^I�K��`OnE�_��)-�d�׾�z���T~NN����}�"����r4,y�j1q/�6x;�)�C� u��"[1��fHc�C g��=�Š>�3�s�	ʭD]��~��o�{��Xy�&�oԾ*�|>�U���ڸ˓C�6}xM�A�8�Jp��b�[.-/ې+4�8��[��H�k�����LeՠS���$Ӿ�g���/3i����W�4Q�ڭ �:w�'ED(NB�%2v�R����fR HJ�� v?���i�y�cI��d�
%�7-]����@��v��y"��Me�Xz���e1�*W��'�L�g���@-I��崏����~y�F�5��E����1э 0��:P���m.ur�q�du�K� ;�,�����^�P������
�m�_�NR�]K���"��N�0Y�@����%���*�7��gX8��vF_U�x��D(G�lM��`䩒�W�9+�k����BUÞ�"�1��wm�3Թ���&���6�E��0
$N	��vQf:������$��Y�蒂��O�N/0>8j�CO'E��ꯒ�u��+��$�io��4�"	���W*�k�O�h4IR�P����M)�1��B��s��w��o׫�g�l���wo��(L��O��l�R>n)��\cpW�{ �=�e�P�����B�OP��:j��h<�xT�����h=�� {��(J%*�V킹/qp�Ω����#�0�dЈ��K�
U~\�G�S�>Ň�D_f݈[ s�x�����D���:�������+�72�g�  M��⛴�xd[|O"Ɩ=b��|cA��?(�j�%u���f����AT�ϪlZPp!~y�12
8^�O�01�e�9�Ywv�f�����Ȯ��!)`:XOG���G��DG�&ݧw��K��b��p��>P��2ɂb�3���61*4�a��ܭ�k����Q��<M��`�|�j�C���!�o�c��+����r��✅��r��	2��~�\1��� ��"�$��t��LV���9��7;�ʌ97S/��w�ڿ�+S�yٹ��9eޖ^�?\Whʄ"U
z.�;c֜��u@I�����کh��Ѭ�����|��9 �R%�o�0��A�P,��r-`^M�P��U����jpe�P/Y�k�l�vm�������4�-/uJ�3-3��l���B�r�po� �-PY�-^dݘV�D3��\j�V>W �$��;�����f��q{Q.���g��ޢ�S�����n��������_8���{�l֤��2��=�з�����j��u.g�cAx}�������	���h B0���I;�|�dJ�U��A�D�$f+-�}�_�
�^���[�rY�֕��m^��<&�'o!�y-����>�z�>�g����a�CL�9y�X̷��NO~�K�X!�Vc�w���YG��ݚ� � �����i4Y�r̓O�j{��&�ʴ0r��� ��HDA-�a�L��sm�����y��e�J��`Ü������2I{�ʬHdF�m���{5�j�2M��3�	�`��8Q��?l����[�ق旤 �h�-�$A~1�qD+(�]��ҙ�s�)D�z�� �ː��k�ӣ��fU�*a��{;h�wX$į�.w��_,Gdx߱�+� �JP�q���dۉmr��0{x��K`��Z�"����4]/bj2nI�}��4����K��E�ϩ ���M��`[�8�����C���Ap3�y�1�R�H�U����Z}�ޭ��T��SL&E�����
q'�)g��1��"K��)e�'_x@Fz*�1��� �Y��FڌI5�)�m�]�|b2����@��}@��&ݿ�e��^&T��孊x��* O�~f�^gE���v-� �j��̷�
���(O��~�Q�Âp���i�fm,6g
�� 1����O�!2 D72���p��|����1y��Ωez��b�x������,	SQ�U�X��[��ѓ;�tT���I[3y9�� 0BX���W���Ƙ���v/��,p]�S�Ɏ�y�i���rtܢ�n�K�h"�����9�8��Vu�l�7}
�O��f4w�/�P�z�ы>�H���	���G ^ق��Y��6�.\j
��Lڸ��?�=���;�9�ؘ|4�m�Gm��U8Q��.lP1�tֺ�%!hF/�h���n�>��]��T'���f=�)��"�	2{�`{؀3�J43fV=����*d���e�߼B�$O&��z�N���������H&����@3V��J��O���JQn�0(X�4�:��� �Q,>�����i��F(�����踼�C�u?��dAVλ;����ߊ��M�R̒��%�����ܘYO��[��E�^��9A�=�IwA�\�5�>a<�^`��z/Poj��}#���(QX��	�gQ1�7ۣ D����}W���v�?zI���[M.�		5Ъ 6G/%g���  ŕ'm��lq�K��Z�@-�(����M���1$��B�d�)$�¥��rB��JhK�ȧ�t���T��	�-�k�hF'>��H#\�>R�,�'LR��#�x�A��UAl��pK����Q�6��P�4��h��[�kJ\[��k<��mG��J��k�(�LsӢo|���M��t���&��+�k�H�1���!X}�����P�n��r��R~��
Q��CQ�/�&���C~^�	��6��pB�M]|�+6�/p��ϭ��$��e$��U�P�P=(�V�L⢭/!�w�SǼ'�XPpCs$��K��t�ʴg��
&����~u6'dI`�!&��x}��6��z8�.�_Qe�'�D׎=�Bm��K����$��a�6�r�kV�ٓ紊 �YG��o1@�m�xmW`<vK��[�=,~�=?���>�&�<�w�<�	4���gZq<�m�F��u�e�Q�:�O��u�*�"�@�~F�,�IO�� ��	�E��f�P_ �ƥ9�"�F�����n+m4��֏9`b����������B��-	�g�ÀH�~�x����.��o@�0��0�]Y�L��`7a	m�6��b��C�+�~��9����!gs�*\&�8,��i�6���>2z���k��c#㻽�R6vfss����_�vH�$�q.��K�Q�����=�퀋�ݔ����L��J�;h����Ӷk�̘��P�@;����2���2�2LL�q��%�#�B�����@y�Q���@��a�!D#���N����ܚ�kϔ¼��u!��s�"��k�'\Yc[lx�<�v��	u}g��#l#��#y��bOJAϨw���xH"N8�]������s�����?��5��!|pf��@�5���P���H0;)Aj��� .� �����ڱ� �tv�9"�X� "k��MB9������[�5��o�(����������*-=�V"��=Uv`*؉[*
�j�+����~�_���HC?a��>%05r�d�=9L���m�J%�ӥ5�g]�"�/G;y#x5�#����:!���=�=��]�>t�j���tH;=|�V+Ɂ���'*����;��J���5?���T�K�<�^�i�9�g8�v{.=]�6�v����v5���㤞�O�1ՃO�uB���݇��3�&~<U�X����bi�i�l���$��ў�1��+'��7�מY?�3<���!ee��T���(����a�j����ZEW� �ZX�lj'�v\c�(�s�CZd !�+�
��[���K�©�̡��זoo��O�#�"Å�s��Yu����ܺU=~���-���9��o�7��IK��*�-���^�R�a2�ٻi*�K��>�� �.٫�\#�M����r=�}�r��?�l�U�9ɝ�c^��%\���v<K6��,%����Sq���|*E�_�_'Z����cRb��0�p�������+��c�����d=����qV=�����D�Z��qq_+r�L�۳���>�u\�Lj�Y@[���e�0��J�;H��.�L��Cΐّ	��_s�ӭ\����	E�[W$����!�B�;%��r���^
�����_�GOX�Ŀ�75��4���:����D#��qi��U��CH����ڠ�]�]��q,�ѕ���v���h�D�mo��x*�R���s����^#�Qְz>#
������eL�|H�*�v�9ƖE�F'd��X�5vlR.�n�O����b�������ap�) l��r�	�C�E�p�V#�Ƅ<1ҵU�n�A������19���JUnp��x�*�@����#�Z{:���D��<M��R<�Բ�8�� ��W��{ /������-����7w9��H!�,⍻��ZOS=�h�ɘ
��H.���4� �DJ��Q�����L~5C�ּQ��k�\y�����~r|,���z�3�i$��3y#o����)��u���L�r����w	蔬W�DgpQu�%�x<�(Ȅ���n雒wq������{d3ҋ��	H��~;�T� ��e��Z��С<�����DD�n�N����z|{�&�E�Z=8X�V��5�����خ�;:.=qy8��aj�oY�kwm�W��ϧ�;��@l�Į����p�[<��Ed����������T'w��^=�c"Y��vLv�@�S�m��s�s|���t���"���.����OX��ٹsǣp<����&��k����w:����\S�)t��ǣo �ZK �t��92�vɟe_Oap]�c�+��(T&ۚ����
2�Mm���J8�cS����4��O��(r�{�o4a�3��f(�� ��/�JI��F��.}ˉ�����Ʀ�CFnJ��XJ�4R��g��Ȗ�p���T.q2�|܄�!ҋ`�j�R.y��=[_`��ve�3��sy�jXSH����;�:�8�<;Z�b%N ^>i,!j�XI�^,�9���N���9�YVuR�U�����g�
����<@ ށ�+WO��t�,�	틥/��}�B�L�ȕ ����0�D`�R�$���(�(UHy�e=M�훼��A���i��>|�v"_PF��p��-k��	�+E�љ�'�;P�@�������P�|d$S���BF��v?����h��x�h2��HҀ�������_�d"�6��6-�����>5_I,,���*~�j�\<�-�_�&i��-E�N�^�Ȃ��Iq)���R�۴��xmILus��ʂ�Mv���Ջ6c8p�.�p�6Qb>O1w���8���z di�8b�S��<X:�3��ZlC��0�:���U&��Tj��R�;Ɓ������Y�Ky��E1O�h��H�C!��];m?�����W����h��dT���Z����p�o�]|�vNs���Xe���������w��Tې�m�m������0�s`�Qk�֒yr��pwS��:ޚ�$R��l�kN�(Ot�H��N�*wf���X�b�ŉfe{˨�����Fa���OM;n^Tfi��@�(�ۆc��\�&���UF��ڷ���f�����jf�A=΅/�[+
E��&n>{Ok�u2c�z�mޥ�!P�ގ8��6�E�������O��:/�wĿ������^�X�C���U`R�5z�E�`,�`�:�'VX�rؿ�\�;����s�P�0�K9��U��oQ�8���_�<�t��^'4�r�#�����d�#��Owa��4^̮\�	\�_�����,��7%-���}rFM֗��'�Y:�7�ѩ]���&�7�]��� �}K��l�;%$�H~�g����Q�@�4/l!�i�'�����ܛT��w��IxG���w8�Қ4[a�X�t�xPa�<�(�d�QK�w�X5��p��>DZ���6D����Y"8���y�y>P��DVCx�tQ|S��a��ȕ�&L�1�����Ĥ�v�8=|;��ݞ�r*f��4�D����4��${&�����s�f[Qd^��q��[�K��whZ=U�6�b�\�ܩo�ݐyU�\Ƹ��5����S�^�ٛ`�0>�@��|����Ύ��� k~
���F׶O�$�Z�Z��]?�/�����T!�h�-������7�q�OO�:lu~���~�S
���J�����VY(��=�x�c���n\Ū��A<��ؽ�͝.f���,�P_Lb��7@�m�5�
�L���\oN<mMJe,�@Y)���1�.���D�����*�q��x��o��a��y��"�����@�66ˍ5h&��y"��S�~p��ϟ�
�]�T��A�$Jܪt�L��YQI Da��fvE�&G/p������
��N1S����ȼKv�%���%ƁO��XJfa�k�`mzd���
/���X~5��j $�3�D�QQ�*�7i_���S_��ڄV�ͼs�ϱg;ԨKN�G�}�;Z��LZ����ÃS�p��=RA���lO�k�!��Qy��H(|�NEn���oG͓zL͛9>�_@eH�虚�#\;�B�U�����`"�WJ�e�����'A�=W�\�6K�&C�"1IN ֻsNuJ9�R���g�Ō���x��}1�R�����]>����~�������d�d��4^�Q.z�3ީ=�1�5�e�w��b��a����b>RgJQ�!�0�8���o�L�{Oa:��(��q��ne
ݘdɹA˙�@輱���{8G�td!�k��>y��qۭj���.Z���#x�V����������vh�t�k�A3��B@���� ͹�UD�P��a��4HE����������'�U{�Y�@�qs�\c���(Z[���[���Bz����g��Y�W��F���"�k�-�)r_�;+��x}m��~��H�.�F{��O���,��dVڢ#R�5ו�6�n�h)�%*����]ӴO�6���M|l�r��IQp^�W�q����b�p/�M�p�|^���(!G��:k���b���P���)0�{��z܍���~h�BЋf�R�����P^�N#rhˊ�`�ڮ�h���ce#BӚ���vd�z� �r��4��\��}�������4�/y\�/nۦ�LJ�^g|<}���_U�{����ƽ&�k�y�og]��_T�$6Lǹݜ"!���dD9�Ǉ\��|�����þ��N�K�&�z��E�ݞt�=3s��T�,A��^�Z�Ѵ�i/WOR�ڽ� ���Ep&a�W$��7��qj��⩫���I��@\&2�U�'m�ו��]crU/xE��,�&l=$+?"������	�Qš���H�䄯lm�D��d5x�J�xV�=����3�u�#����&��Ot�rƟ/�(5e�JϤ�u7?�LJÚv%C�SmC���V&���E����XuN���� u��6V���L�Dj;��o���Uu�oq���yF���(Z�$'4E���#�b��	e�BC�7i�ɉ��]����l�x㍸�ؕhx���Ƨ���%4 .�5Ww��.h�]#1=������+����G��o�t�v�����v2�f r��NiVx�=b���a2( �4���y$������M���a�j~��^h���g��Ű�X�n�ltS���3�zVFA��	�_�ez��y2ɹ�CI����"v/5w�/�qm�����n1����6�r�V���2��q��f�����`���Z�g�Uߩ>��)��^
ZXF�y�rJ���T����U�눗�#�. v�m0��1���3P��lG~$Wu�F�i�e��F��e�X�Y4��ͭƶ��,�u;ZX��]C�2�ȟ'j�*c>g�w���t5�*�c�QX,*��k��f�~}<���?4�ʪ�
i%?m�Z�W��s��В�قˀ�sR�������|�R�]m�~��Ec*B��Sp\!c��I��4����`������+�E��J��!%w����z�1 T1D�\,Kl[a���T���BG}�X�̷�o��8�%	u�79��
�2<g`��%��7��&�����S '�B��D�F��/�,04��֫��m<eɢ����R�VC���fa�Q/�Jǳ�κ�X�=~`�˯���Q��ftS�&�� >B���7X�!��H:�}�K5��}\ZW3�
	�>l�Xꉴ#!�.X=+�7M�)��@�[W����K+��(���V;�{��%~����16�Jݤ�QJG*��;��uI)d	��Jl�?���[y �
�_�hr���<���iGe��/G-�&�9��ɋl� �B;���0,�s�|ű�����;���n-9X��ؼ\J��ZQ�k��{!A!��'��)TAu�.uG��z���\��ڹ��Ѡ�V@�.��z��H��]�����W��j���xҥ��LTŹ<e���#�M�{��A~�Kz�Tb�İ?@�O�۶��'�Djצ#����Fpq��+��a�!rt��.�|�V.���!d�N��b�^�ص&��w�?� �k��n`����!�do�;�8k/�� 0Hlƚ���`'u��{ݝ���.��Z ���=�4$ ���E��Q�߶(-+kxr�+�?�Cu.��J����)�g�?X+=v�F�@��	�G<�IH�m��C�>
��88�T�"�:m<�g��♚4��#��J!޶p�N���;��乆. 2fz:��c>�21�|�_
%�g=�Q���aV�;	^��i�G�]9IhV�����r`�j�М�2	Lv�'t~�T�[��doQz�2���J)���#^�<XB�I�ˍ0��|*�ڎK����4�j��kj����6ᕿ����$$`:�18�����������9��Ve킀{�:"��E?�:��j����Ps��Z+C�	
��2�GÏ������8�(�*�̕ �%J"52 v�b����xH�4�r��8�a����zi�f�çpW��
�B;ć^��PP��/�Lu�!mu��-�q\����c��1�&��m�t��R+?d��/�:o)��)��_�p�k�������l1� ���3Y{]i*or�q����A�L��p�J����hT��Jk�͏�b�Zi�c�WD��V`ST%s��!6c\��!ԇ����!�C;��؜�Վ�J;��1 w�ߑ���f�y��Y3'>� �P�0ꈗ�a�`�ð�6�\��!q�դJ�\�����>�p�v�-��I����g���F�yE�吏w�Jy�Q�l�>����'�Ӄ�N�,�&j�+�>��گ=Ăo�b)%�I���J�����h/�@Ɋf�)�E~���t׶��ͤ{��� �m��~�@��i���s�ZE�o��ߠ=?)���E0��Y�_5�k��@=-:�^�l�Z�-��������.����2���J)dY]K�њ�u�]5��N��c����S�.t	��_�����S���� k�`���:�Jlez*`�z�QΓ�/�u~'v�Qq��ﱙ��WG��9�YI���]];��ߣmM#�8Jw�;$�A_��E����%�8�U'`�/����F�6coh�'�����AB��:�EF�~,x��	��h�n�������A�6Ϻ6��{�>�|��b��{��O�+��6�6�	2?���ͅ��B�?�̅ybgm���U D���3Y�3$�} ̅�
J� q���`�u�M���	%e�F�~�yOxíAr*���E%l=2��0Ʃ��ƻ���ֈ�^0�叉�C9�F����"�;��5)��|�\ m*.�-`��`�
�S��鈩4��;
�[� w���%�~���љc�m���U(Z�[�L��6�|j}�B�pٓ/ghTڐ�)s�E�K������6~չ;nI�HLh�` �tG�:��i�Z�,զ�U��pc,��!���|(j�s��3m�<ݒ�sҎ�K~ln�=��0��2^}�:�Ɉ�B�ʙ�!�����|{4�K�����PMx�}&X�v]kb�c���v�k��l����u)�[�O�@������&��I�DYA�^!���A0i�.8�U��c�(9�^������ܠ���t$g�ê��}@0�d�k����FuFfŴ�D�I6��9���Y�^���8"*m�]Jn]���s���{7�P	(?9��f�ѯ@F�>��A�ԛ�g.b���!�2�����D#����8���d��zA��,?���gV���s���ʩ�yԴ
俁�Z8f�>k-2�-ug��X��f���]/S�/�M�_~E�Vt|��*��'�[X�&�:�Օ���~���tW���[�0�����{<����,�ՆjE��~�WJ�X�݊�\R`S��{*�v+���6N�
�w�@!���_v��+�.���F8�.s��:w1I�Y]���5��'7�%fT7L�y�N"-��bXE2k�~5B���ӝ{��B^��#�?Q�-�F�deH@�2��i��7X�������F].�hj1��+�Ri�����q�S�a<XUЗ�2����V��?�Vf� �)�\��WC��ޭy�Vh&� �Z�	�9%�P1J[%�!2���R����T��.J92ȩM�����҂�RñWǖ�̸�H.�KY�~�jC��s�N��U[�{��`�����R5��9�-�)��W��܉�/00
����Jq��8��bGF-c�O;���D�}%]��ya�nvlՎ�/�}EIg��+d(�m����C �ѵ(�"(f��h[��2y��PKz��(���Bm�����8ٯ\�,���"�j�":|��2�>_���ү[��A>���)�$L��EBj��
��%{J7�:X/4��U<A�K����D�Kr�4M�=���2�]4а����\��0}�͗:�Թ���*����N�oƯ��F�^�i�Mg����#_��)�9*�&�Տ�Ƭ����e3�����
����[�a������Kb��4���~���=n�=�D2��0�C_(+a�5O�Y�|#HR7d,�h�Jn� ��2}�ȝd��a H�f��ɳ¶9�G��@-C�0BBb�c�
�X*@Y,�N�����R0�!=F;_w�x]*߼�>�dY����h�.�'�1�2�@���*������Ii�V�	��FY
,%K��Є=��Ĵ ۲��=�A�!�?��8���)ԍIo�n&�{��.Z�$�2�{�a4��1�f���Q�u�v#�S�a�Q��2C�P#��d�x9b?G���a�(C�q�|~A�hSR��H��!�<�R��kD
��`�A��3&y?�ٳ�*)��c��������D�y�^�E2���n��)=�t����8�4atG�'�'�G�탶�$>��������d�V��ܐp��~�g�!b��(m�GvH����3t;�}�s
I��ӽ���n�����w�C�	��F���:�>�KekʑZ!_����;�B�_>�"��NgN���x�����])��w���y�;Idr7����7�v�?XP��a�[)=�b�
�{;�l7�'���o��`��Kd�`��%7���8�����V�VBF�>Ecc�ڢ:�x�#Z��q����"����ti��d���ȴ���B����%8c�p����=�s�@�'��1̽���sK}�2��'�SLT ��{�j	zW�D��5��7G���k�)�.D�:������T�>*���?�qX(�/��k멿ºZVUg�n����K�D�&�j�ܩ�#��_u:QR�%X��$+:��b?�����1��a6�'Q��{.��@��\'�<�KK������|���bd!����eA�@0�W|D" s������|�.�v��f�2�[�Ꝑ��w��0/2���!�b�Qn����kK����*�E>=	�-��o��d%B�QIC(���λ�B~_XZ������u�R��u����;���C������4e!�3]b�;F0����Vf1_�ڮV-���<{�8�z�fD�+G'l ?k�L+(�	� }�}��"& ��x�!L�h�{i�#�K3���J*eh�y^'��b1[��
���;��(_ H\�mmex�L~�$��T3g��'��j~P�v0�M%J|$fie�Î��,>����m����]��k�9�w��==��d�<I���|ZS)3� �b#�j˟��x;�G.L����晠��kpA�
BT�����X4L�ޏCe�����r� � �X����\�'�w�E���f4���Ou����"�wĩ^,z�3��l��`�e�.��!	��/�y�]~��⹕��v�Z���Ϟ~5�a}��:��J'�����h{��d��)􀅂�f��=t*���`+��#��ϯJ�p�@��u�����;\L2<�X���Ŀ�J�m^�w�;2�g���c��FbJ�X�����P����i�� �mIG[
����m#y�Ī�_�0�K�v�o�R%!����k���wo3�=1�$|/ש�C}Z!!NK���,j�N� =\8�vArn�\��y��+p���ݶHFXoS��o�Q-OJF�@��I��K�l<�X_R�g�-��q%ُ_7�x�=N8�+K ��_8�:�&֩=3��#��FX��<���r=}�*;�5���P��tOR>��m���W���\r{�a�Y���|�|E�����߶�AH�Y�<���w��]�&�-X=�V��|��v��;0e�Pl�!�u�Hͪ��L��@hy��x@��W�Fg37u��]x��vH�2foj �]��	�W�]}.���ab"����&�9�a����^��`འ�DM�ڕ��*ՀA�?��^�R