��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��s������\�Ἡl-�y�f�����f� �ѕ:�nA�kb-q��_���ѹ(4�dê*���7��N2�ɐ��+ٞ�4Y6Mx�ejǴ�y9�����=���D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�!��
��%Y l�׾�U�����l���M\�;˝�v�HV)�uE���l�>p�R�o�C�pT���
�:H���ʱ��y_&f�n�U&��j!߳��k;����(���Y��e�S ���',�cf�ҙCsW�ʊ�`��g'b�w�QH#i��'�?��N�ϒ%Q�4��d�3��SI'T�:N�cǢ-���7UH���Z�UI���k�h�	ɺC�6� U%�F[ߥ��չa�j|V3�!�M��[.�_I/���_੷}<\�b��[{�� x��4+d?<��U�-�$hڠ/��(ѐ��	^��Ze��C�&���˪Ui�n��HT?T���U�R�Rj��x�63��R �O<��s���w��]R��$2R�Y���E�zݲ׺\ޱFp�_?�=U�;Z���p�8��J���PeݶRLo��s�F�x,tJ�-`��m�tG�W�`�sP+EH���[i�T3�3S��[泑כ��,@����K����у���y�X;�z�`��2Y�Q%�:j��hi"�\�@�=XR�<Qt����;���|�-�L�Z���&)�<�F<)���9-©=����ld@l�v�QB�T�p �R�S�|�m���� f�Q��漃o� � �Z��物�2�=��O���zC%��,�}��=�X(A��z��i�;B΀h��<�s����]���Rw�hT8��:�`FO.���5{L�P�c��{]��\"�W�K�<��#\�K�n�M~�dJA<a ˾�4	�%w�|`�?�2 ��Box��^K
�l�9�)8a�)=Ӳ�U���U�3�E*��%���bӪCh�7n�t"�$R��e� R��s�	��"�����l�� Y���,��=��ᚪoW�+�.�����& :�Z������ۧ-�yWu���k!2'�z��,�Ly2��q�����{��
(n`�g/���S[W��Ɨ"���3t[�d����;�}�	q`�/���^��7�y�" ?�C���o!W�´�=�ANl��r�k�����1�8�s����k'���h0� ?��IOP��	:�,���Y�x{H�\�����A��e���S�*��}!R!X�j} �l�eؑl�I{���p������ a�'����o椤�lV�N�["i�>A��'x�~n-*�ʧkJ��Q�U����͜��Y����ʎ��-�	���"�@���֝����F�C�[]?�]�"yXp�j�GJ���*�a�S� '���a���E�!cw$Ń��q�q"6���?����vm&�1%�?p�T��B���WX>� X"V�>�iW.�w�^��$�9���J���Bs#ѽ�w��e�Н�md}�J|-��xU�i"�b��1֛���:�=>٥=�z 	sh�_+���=������"��.��V_v����/2�/'�8��P�O�W#I���O�>y�>h�	�� ��|���γ$I�]=��$gD��1�����!й5Ĝ���ϽJ�����n覆�U�9;~J�Y4�ld9;
�+���&��D�O�N.��.��X�9)6�.�pU�Z /zM2�m�)��U�!c�]���dn��͍�)}z:���J�]bj?6͹����  P��x�#a7��� tV��N�CL�F�,.��#T���[�r�$�K�
2���s��i}�X�/�W��I(}X���w����:5�E�[�z�j3Ee�6^D���t])#S����b��%À(M��g$)��h�g�ȥ���iW��O�s
1a���F&t�����{>�O����A��
�攔���U$h��1��ޚ�N}�z�[N!$��C�r��K�-S�$;��4���:Ν!q�=�|�N�%��9��&N b!v>d�jif��Zy'�7�J������Aj B�Q�s�t�63�.t�*Y����VL�N�,��q��P�"�yI��5<�����>��T�S*g�Qn���h�J�|��<�(%8D�!�V䛿(�`k��k�+U��t���>�� ���4��kT���S;��l
���(��x�ن`(+�%]r2����(%��;�*�m�ܚX		��̰�r{ٓ����B� ��������=6Y-?T#I98�A�ӄ.L�ٛB��-(�ư�4�����c�b=ʂ��smNx�DL�ui�>���&�|}�pj)�wS�� ��$��� �U��($8�=`X�H�ef,��K�rz��(������t�ӷe����2�`
�����1>�򢒻�3S����kݸg��y������9v=+�<�Ɖ�W�Hvx��7�x��C
��%�>�D/�C����Y��߫����������Poq��WdT�����K�;I�0��$�Ce�=ޖ��L��p�4{� �~���]	Y�|,˔lG!v{����}�l�
�ᮖ5zc���ѓ��D�������`�&�����M��5�O��h4��W[(-��4�L���R�?ec�����Β�3n��N:�Y'@�+L簛o���@>ٷ԰Ȩ�Hn��@�H�JEB�NuJ㱎�X
�aN�U���&'������%e<l)��C��0��{�M뤆J����=�i���X�C����qЁM�xqZ��:u��v`��-��%T��� Xm����c���}G(d�DŁ(riY|�W!���6/�z���r�t>��c�����11%���;�|�+�G"u��>؟h|¨|礡�
<qr�w�2(s<Q*z���9�??�h/���$����u�	I��ς���AH��c	(�qh�i���$U����Rq3|��>��\���_� <�zC��{蒕F/�%�u��#��&�1�׋�?ԯM�n�E��-[�
��s��K�@�6�D���l�W�%�?L�5�s�a[��eS��<(��>��@�!~�8���I5��xzF�i�yt$xא��Ӕ�`�t�/G���O����c��x��
Y�s2׶h����+x�h��6p�o��!�<P>���Қ��A��E�S@�**�\�A^�ENf+���Ϗ���Pu����]���q� �Te��8��c��;
_7�O����]�VD��nS�����_I�)D�x�y�ͶR�R\a��n����;z���]��Q&o�K�%	\�q�������D�µ�.'��|��@�-��-W9=I@����<�gg�|K�}쇎#�\+�8:X�(�>{rI�l���|jϦ8�j��l�{+�*�����!>�����3��4U����ͣ��$�˕�}']+r�������@Et6P�m�ZAD��8���b\�˂���)}��nl2�׬	Nk�S��F�t�IY�=�뤋pZ`��0�v�e��lLك�&���ύ�+�C��C��T�)yV�-��R��'yy�P����Y���)JYI5��R�H�^������,����ms�;��H�}�FhDG��z�]y��6o�BOh�v0�\vߣ�dJ�8�cMm�q(�<Eo�cP�$�DQ�_h2�!p� E?�!3��^]gS���|瀎�k%���i~rDqKw�x��ӧ�qM%�6x	�"F�5�Wmc�sLc(ۡ�R<65�;����Q��?�Қ���������]y����5�Up P�A.�^W���`0���N�]��F���z��x��;a{L_-n���s��/A���p�`�v ���1y��9���nRf���9M���ţ�����k�9(��{�r����{�]e�Ì/�0���8Bw�1�\Ǹ3�3��T��]�����A �P,��m0=��#�p/u�'�����P?��,�֕0�
Rh��k����ZXz�ۍ^��8~2a�MG��ލ���}T`:VPjLMOƸ��e�x�pI*��kt�i��Q��Y�0@�?�y��x �v��H����lz�7)����w5��U�|n��z/�T�o��:}�f{��>G�Sx���'
6�"Ζ���x�w 62��������Ig�X3 �Q��B�/�����W9�"�mf�.��7I� ��8�(�UL;����i����J��tchp�2C{OeX�l1S�ep�
Y��CΠ�Z�fϸ���'�xN��)��7PlP?�Ti"ة�ֹs2m�w\�yvuh��Xr_��HB�����L��I~�H�=�����З��D������в��B\�լnnO�Dz��jJzPQ�b�*%��V���E�M�]�[�k&�(n�*Mi�^� V�����E��su�'�4bS(]��0�2�����;��,'�v����e�|����ൈ$\���"���W���D�n�Z;V�wa�J�̊cmAf�Z_�Cvsf����m�Ӕ�LJ�@ᵿ$}�i���սC���ƬT)�2�+C-q_�|�A�-Ӑ_��N��l��� Ƈ���a�4BD_�׭>D��#�9iO��Trt��_u��13��:'�e�|��x��ne&��6.{�ăTm�_9e��Y  D����)<�d;�A��uE���$�͹p���{�螐�V��7�FIRf�&ڴg��^k��2Y��l4z�_w��g����4c㣯�t �F�˫��"N4��@<���QƉ�L[�����<��;e��j9��u�:C��k-5�&�(���avתz:�x?9����"h�k��+��ˊ�q~]+�OT;��r�u��?sioI����������]O��7�
�j���i������~�- C��L-�ed.9�g�!vCq�Zз�1ʅ-^� ��c��GW(T�+#|ZeƦ ͈�$�� �)�E "�MV!"�K�/�,)���N�R��@`�����a(SԑJ�J���@=\�I�B*�S(.���S�n��_>�n���t<�ޘ���Ǳ�6$�;��t	{��59Aז���v_G�&�e�Ƅ�Ff���K�2���]�S�W#���Q5H�5��Fl��	���P��B�-l:*�A����+��{���������'N�f�{$��|h�yj�;����s3$���/o�S���⏎�a��o9t��Յ�_���r�(^\M˴�& cJFf?�{����M�l����'+C53e�L��q%[�7	�	t���ͦ;�D������:9a3X`��Qۮ�d��H�1y�é�iZ�I	@�n��4wU����`���cg�iz�f�-rT��I�t�mx"�}
q��E�#��b�ǆ�8�Z�z�L]�r��v/2k|��-ў���kA�yA�:�8���/Aֺ��tAcVmM�7La�ڹuNT��w@�:]s����w�"^Swj̮_L�ZX.\ݢ�2�(��3��3�G������䭏x��c�C�b����mD`t}�(���~Qw�j���y1!�zǼ�e�}T�ĵ� [+Bm
3Ŭ,m�(�5�BF�5b�獇NDRl�x�M��dEu"�L��ej�GQ�+C�e����;<�n#t�����#����3}�c})n�}>%��㻷��0�ʾb*��`FA;f�zz�.I��}b/�LD�g�tX��J7l�)FC�芞Q#	5!�]����ʙ-�����k/�UÂ�'~F�?p�����	�C9��P��_�~;qc56�ƥ���3z����9ܻ�s�~��nH����{�gu�2���r�
�	�}_^�n"e�m�"y���EÅE^k��
�4��mn�H$�oO 5�]�gD��)zU*NĘ~�\��o�+�E���ـ�z��ܒB
T�Z 9�Jۍ��ۙ���<�Q0���R��4󲏗Z��|{�DjvsȅZ��/x �=����$�6�o�e+�[�O�DӎH�u=
F1wn��n�?�`[>Ņ�9��@�c�@M���)C䰩���v?4��	尋$���OO������y�e�S�)j��D�<C��O,I�+˼U�d�i?�[� ��)�-\Q���%\���t�ҥ���nͪa�z.]��9i��)�����F�Ⱥ�+w�dr����kOD�����a�m�k�4<�F��݁"�;N��˪-��5���N���{qba	|e�Gfz\�ֳ�ʢ��nڑS�n�Y�qz���N�O4�:1��c�����,ZU���Q[�E���r)���{�>[��j#�O�aAt��T����-�0/���v�����^x%%=�\���VX�,���H���%��p���_�P�'����]��NOZ�V���$�W�m<|a��;��Ŭ�l/t�Y�z��Mb����'��_�(�6�R${���̩K�a��H3�x��e�0��5�:�r�<��jiw�Fk���_����6eG�|]�n�@�7"��+�{I)��ez��wy%�K�N�C�0�奘lCYzOX� L��@��0�|9?�K�
[�9�1�힘dxci/�<̒�6�����.��� �Zy����˞�d�l�f�ȼ �f����Kˣ�,B ʃ�V)~i����6\%�ȶ����G�ٱ9�F��W�R���c�zL�����cY��e�Ȳ�|�)���8�|��u�B�:����@�:k{��1F�6��{�CD�R�d�b)�Wf�,���`V��ޓ���B~;	�����Ò�&r�b�3c����.ZV,��^3|�#�1� �D@������v1�!��(]DYѹQ1��g[�����ꐆ�V���6L�5���&"W�NTDD���K6��:_!uF�FdY&� ��:��"q�Y!Oݺk^4���~�����w�d؊�E@ܠ3Û;{c�a:�jQ�:-�Ϣ����!B��P=���W���o�1�NC+�?��0p��fJ���XZ4N��I</t?�T�#5Q��x�@��#7ZPRR3Z{�I���+�����5���e���_�\�Ry68��5�D7���*�����-meh�����>_�{.q�8��퉈���-�/�jj3�B�˽ُ����[L� ��ݨ5T��T�}(�G�{�\+��K��=��;,3�@�c�� ~j�},�bqf!�W�yNc�ǁ�O@Б��F�d�X��'�l��\O8��SS��-�$��8Se3Ήfǿ�)1xu����Z�:�G��!r�_�s�>]>j�3���rs�K���3�|[Й�2���?5	l__>R~ˁރ�z�}p�_jw`#�hs���$&\8i	�bK( IO{(NP|����f�1E�'�nC
������D��g�Ɋ�lD�5j�:�9�S�FBm�ģ+�dj�L��.!@�v������_�n|O_�x��p>�jF\�`�p���}��K,˦K�e�K�"$���le5����\���o7@/k3�������,�\����iZ��`�ʟ$N�*�����9�	uU�.�Z)%x��ˑʃ͈�	Y��"\�u������	�睁Xj t�s��XR=W���4l����*4O�>�5��z�U�t��(�v?�-8���g�dmR1���z,X��ds�E�.�&�a{%O]��>��)KӺ��#�*L���n����-M�b2	PA�gI҄:O�V>��X��5���0������&B�8ӯ������B�����{Gɬ-ܔIv�\T��o����;��,2�CR;)c�Hm�v��{�⩯�j3�B���� ����0H�P���>�%�J�_�E�^P��N�w�l�I��2�Z��&
�W�&��o�����������@���D��\� �V�W�g#�f��j(�㝓�����>���
f�M�a]ݓu-ߌ>/�eΌu��!�h8c��i�>��(���c5m$��!��#���Wޑ��s�亄F,� Z���j����V��)��v��A��\�����C�,x��M�qrX�Y���C"/�R=��Ւb��)!�32mZ�zK}���y�ɗ�_9!?�w�{p�dz��q^r8 x�[�!�<�jl*H����Z8S�L��z��ߕt�:+�h�n)fb���$�2#�+��;�p�A��R��<Pǳ�xo�1Es(�Э�+b%���-V�'����l����hW��材
ΥDm�������u��ε�-E9w��:��.�$q��+��0��2�ڄ+�}�T��A��3���h'V�st>�7<��W�Wm�/$F�V�p3��0̈́�1 �'cI�8͌�53��}H*�D>��Uj���O�Me��|\��� L�FO8B�G���������	1*�n$�1�~c�:>:X��8�a���
�/�h�fa�� ֟I~�;��g3�V�{3~��? ��K<\��H�+�tԀ��͟]��jP�̿�?� ����%�w:��z���,��͕7��,Z��mj$<���f�^���;n�T�tq?�JL��Mש;D׵�,����$Zﱌ�����U`�N=�0��
t�o���z�Y��C�\`�^bϢ�����1��9�,0�^�gy������ҡ�X���R�za��â^��9���h��o�� ��`X�U |��ۏ	)<oQ̟O{���h�)R�\�Z���J�17<@:_`00��܆�k; vO�&���B�:�Rx���ن7+g���K.��{}�C&�v���ߍ��~��f���iA�RA�f����-��%�AiKً�k-�CF�EF ҙ�/��Զ������:�}vg1��ĸ3V�|A���(�%���F�+�u3�I�`;[R�I����X�9@�)3�$��@Ҁ�u/�x�����,�iT���<��GÑ�7��]52IM�u{a�o;F�t9�UB(?v�u���8��1,�Mʧ�es4P���s�|��U��8��]�m�T���SW�0�bg'�B���q'�/Ͳ�G�#�$��Jt�ě�e��s Q��Ufֈ�&�dS�H-�Z,��4�@�
'���݆D��W��-���M�K��������a:;U�ģ(p�e̊_�N��+?�E���K����M�0n:�y�^��0�t�o�*�jj� �ϒ�@9:B�D�NO�a%�/�a�B��@�%��������}.MC�;�)�TVo�+�b�X�:	�ӷ؍����ujۤ����g��,�fS��+�"q`6F6�~��֪�g��>eQ��9j9n������xŇ��j�5�h�>F�h �"��^���em&/`2�<�h��g��%��d�\� �q��It�V�G���-�t�.���W��4x�MC�8$��U.Z|���{4�a��y��2�U"u�`RhnY���NBi໌9��UC��jL=�ٟ�rmZ[[.NÓk��m�Z�fWp�<L��������zٺ�@��p��$���m�%g�,oi�A(iK�~��q�w��U�+}0�h�`�-󆏠�~����q��%v���w0�ο'� \��t��<IP@��1�+����
�Kt�0�i"*�/4���U�&� ��dI]n��)��(��+,O6�={���s	o�~���Ai��&e�XE�)�#���p�r���T�T�:ru�ʎf������4d)��{�u�)G�)�B�$���yo�m�4O�uֈ��X���=��_���w��5.� �$cf7�aP>�/qfh�5T<-�g�Q�7�\�Ϲ�"[l�`��d�W��ڸSXl�K1	GE�Ӭ1�����F�iU�7#:k�6<�� ��)A&y~Ȇ'#ֵe�������^���f�����Pڃenք��@S��v���,E:�ڱ_���;yPvG�V5Lmr���e���7C�U�oD��N�5\1�V��ktt�۰@�zz00�\cf�P��Ue{�)XV.~�#NZ��]Gg^��B����.��'A����
Q�F�(+�?��18X�`Z�f%�falϔ�����]R��Ί�d�r��d�8Vr��\σ�H �a]���um���))8̛�}�^����o���Y���Y�L�O8���[��]G�,���w���{=y�#!��+�����CeϘ�o[�_|����4t/O��	���X|�]�O��@=�0�P��l4�	�x�7�r�5����������a��D�-6aX�h��s\n��H^�Ud�Y�Ц@9�˦�k�����-��	I1S��~:Ա��[�ӡ�$~:D��Y@BD�	��'B���j���ȝ����KG�@�_��(+P�̫u�!A�!�z����Y K�X�4r~+bj)Z��j���[�=� ����{�6P���J1�BUp�!���ܭ\2ق�I�p@��%hG�%25���p������iQ1��1�Z�ž�>�-��*8K榷�#Hl�-�f`vv�)ΰP�f7Ә~���z�_�י�@�,�Fug�R��eU���B,���ᘎ6}k�|�#��x*K�HG=m�S�\��O�+;c�� �5I�0�U6W2ӧ��/L6�h~�ݫ��⭆�A��e ��Z�t��Ky?,��sm�N��L��V���st��Y_.ᎊ�dm���3i�A�l�[��3\t�Y����?j넿�q�D��P����P�K%����:H�dl����H�� ��y�z1<"�5���,_��]�-�d���zIE��z��+�<���y�Ivc�F�-3(�gS�����ҍg�T���X9��w���r<�Pk>�C���!�!P���K+�����ڲ\'0@	�Ú��<����3ԑ�FO����R$��ͺ��0h���͹��JLe����;�k�̿�\��|5_��r��+�ZN��`2'r
��u(��`ʽp�Z}���1	��x�8���:H_p^�'RmHT�
U�=��tG�T�k� ��V&�ɑ���do���΍�&�Jh>ة���3ee�i�w5u
dqPZw����(ie���ߠ�7SXw!${D��{�	(�7��mO�ɮ�U��<�m�bU����z�~>-D���l�00����U��)�P?��a���~l�Z0>ě,��yP���X��S0�nԾ�������r!���6Ģ��ܑ���Μ0�GF��D� �7��V0�{��<z��&��ؕ�~[�Z#��t�F�񬂓A�ِ�S\Y�7��ˡN9c�4U#�5¾C�3%$��%�Qҩ�p���Ĵ.�m�+���~�di4���"ge����s�CH�9!����h1��E��\8��������i+��M���7�<�{}����5�awr�6�XO>T�i����B�5�r�{J��@=�SXD��C����l��#>�"��<�aގw��Jʛ�-���0�"U�u�}7��mb��4�JN�hs���H�Vm�6�٨G(�ŵd�U�
��>Q�?K�|M�YZ�P������L�>pFM����ɲ�c��>�S��?�|��V�=%'\��zοW��}Y�}�#��ދ�ޥ��$.H�c%��j�q���@�#���W*―�9U�d��u8���[��?L�C�Y7�Đ����p.������N����$���`#�v�6�����0��f}g�|�q��A�=l������x�c�P 'N�S��ī<�����֮!h����� D��6JPQ��lܙ���__�VQ�3�"�,i��KD�w�k�n_�e���E��O]����7&���ZrT��j>M
�h�i��8���P� ���ʴ�L�j�[ZaQѝG~�w-��MhC���x�� �)څ{Ѣ��Mҵt+G�q�eMp��Q��}���"�x}�-��+;$$�Tq�"��ۜ�εhoj~��
�gz����2��NǱm3��R��'\���S��,����	����\2�_�BwM+��-5�>��`P�]S������[%i�I��f�q�[�����ݡ�/�JHׯ�P�F�ܼ{�9���J"ӓl�7�W�z���y��SB�`?*�ɂrk�}'D�(�a��7���7�dt$d##J�Ň���K�jx�P�u1��=����D	9���pp���N��J9�c_C��O��;���8E��P�)o΀ʄhMjśUTǅ#��>��!����=㦬����8�~	O�_'Ao�@�C�ʉux»����i�ԣ}�'��`�kP�R��!�"�i9��$\p�[�Ϝ��s�%V[�h3�ek�ڀk{ېhAf��./�D����3�.8�	��>h�{��>���T�eVF��� h�AH{��	���������g�4ͭ7�}%x���s ԧ�VĊ:p,$^�+������<���f�P�v^#��H���d�Z�46�E/ј%P9���*����&�?}�Ռ⍟\V; �+eŶ\b.�N �l��'��$G�=�dFU]��NRN���]��z��:Ϩ\�L�Hۇ�v3녻���:/�;�T'�����:2Y0��S�DK��6��՜49B#B���!�6ߗ(�W�kM$�)t��8x]�/d�!�D)��.�����;~c���'Pbo��&��:�@q��^&֎�v�8�轅@u�Vŷ'�E3{��T���O�D�zc�&�P�M��߮���\��6#� �AZ�m�[6̆����Ȳg}S<�� "���|����}e ��q��'�e��!
]F+q��@�<I�n��n��#E?Ra��uʭ�LH�̥�����.J�FZ���Ui�j�u����N�����K~Q�(�P�ЇV0�W�Y�W�9�O��
@+[�T��<1�44��c��X�����~����� 0,�B�C�c�
CVM�Wß&i��`?)���Cu��\֝M��:
��c+94M&��иy�}u_9�ay`Bz<�e�[Vv �0٨;Ƣ��E��9�{?��t��B�Ȣ���p���h%���Xv0$յ��fԵP���%�4Av��Q��Ax֐w	�8�e�cu�D�Vgî�_P/�rB/�j��t0�r�BA_�6e���b��d��L�<��M;�D����<�Y�`HBC��ȎY�j�����di��t�ۙ�Y��G����g�3a���k`�VE縩��#q�i�L�P�Z���`��\��21"Ů*�B�O�{x〃�Q9�{TI�%��T���˼2_�A�i<O>�<Qw��q��n��vL.s��N5�Ƈ01�j����&8p��)Z+UQ��=ۂ�~�v(�avBZ�^��ZA���1Ɉ����l�w����\��X��'^���$��Q�����ƥ��k�G?���b̖��$y,	��(� �g7�q�zLYʕO��>�,Hp�I.��G�����<��&j2	=���K>�{�TS�u�����bR���_|�� H��Up�X�sa���g��KK�*Ri���}���<5�4e��{��J�ߏ���?Ee��d��q��$���V�h���YF�5K,�p�f����_r�p�p��	I�S჻��4SB�T�������H���Պ�Y���"��"mM�S�� $&���S/o��
��1�-����(���M5�RL�j{�
�me+��4��E�m�#q�IZ�)���.�"0���H���R,��]�ej�Vk���٦1u'U$|>��wԍ��u�4�	H��YxU��bR�ܟޚ�A�^㥂�y.Sa@�)��J	�����Tԡ�Bգ�^��B����=U�Ru��:w/��^�:{35w�Q<�b�M�a�@��r��̀#Fշ�j��'�9���~�L�'��- ��s��O�'z��-�G�	jU�%��ejZ�i%t�ZK�R�oܰ���9rYK}����b�J30�^)�o���~"kC��y��Ud�-�M쉑�a�@�Cb��,aNe܆:�3�nz��J:|I����E�ʹ��$3�������;&��lɈ��0-N燺H�n�I2[��d���V&��y-�(�X��$� ��3p(�C��zT#*��:�����w�����̟-�UI�4wx��E��vĈ0Y��X��0�됕iC_��F{�nF7�(��e��&g^��H�G$��5H|��b�D���֌�p9gm6J�Ě5L���˿hU�kTh�԰1^��t��T����%�@܇������;��cf_��l�&�#�[���zC����7BÚ��A��B���&�<!�}������	����vr�ܟ�ʑOi��鋆"%|ǈ�Bը��������׋e�Sp����oѶ��:��&8�Y����R5J�r��%H� @�b���]�銚�E1ųh�;#<�+�n��p��bX~@ɒ�+��O����A�=߰)��p��(�cD�k�{�}��c��taW��:�"�Q[>>���^�f��{z���[�S���)64�JQ�;Ux�H��5� 	w��Wk��'����/�>k�FjHfZ���+.��o�ԸVK�a����w�G�L4ב<�G�ȩ�dA=!2j�$�'�cjN�zw���`���<B����3m�	�>_k|y�M�Ch�`O�,"=��TK� \~�7���+Ѩ��NQ�y��Rx�1uT���+t%�_B���Z{2���&�HO�u���>r��i�����;��%�]��l_Sx��'������S�]�[��O����9�ԉ�=�$���6ɤ#koՙ����OT����; XY���Tv�Ig!��_ q��d���&	��q/\�:jj*�8��c��;w�t^��xu_�G�4w�b�d����\4B�=U�*�{v�-�{!��X9&W�ԕԐ/v�{�����x�� ���Z�k�I����TGf�Y��(k��@I��FtAw�h`�7��;xU�0E�V�\�����k��K��U:eP�u)����݁ZMy��;j����M�?i=�Q~a��{40Q�#���y�~�zkۈ]e��be�l���g���v/��=���A��P⸖�}cHC9�c-mC�D9&æ����!�b�})�=���Tw�?a	{�=k#6T�U��p���m4l���cq9+��N�w�`Z�V��2�%��x�i�O�B�g$WqΉo}�F��K��=,/��0�06XN�����ǧ�'G��*��=r�f���ѵ�Ty�
�Ub�#F�{)�vT3j
V���֯�/?2��C)��D��k��J8��C�C�c}TǗ�e]� z�v�3���gv�O�DI�0��������Vm*3�	��|<��q���-J��i˴�0�� 1v��Ut�bJ�n*{�'�3|�ݖ3:����,uO�Y�k$,d]�>|�����I�dȄ�&+B�m�
�&2[ٷ}^t���U)�#�����|E$���΃N^r�Ĉ��@R/%��\Ѯ#|[ǀ���e�!�]�W��$�U�H�XȚ� ��
����\$w=ؾ���Ը��y�<a��BmIǘc��C���0BK�֭�
^�:�t�w��I~�au�oT���.Cp3?鱫)�����$ާ�{�o����QT�s�#�W������r�Fm��!ti�D�#ܣ�o���I̽���LQ�0��� Hq5+�1O/`o�;>�;bt�_��y�%͇���� ��P�ǳM�Ԛ�Y��U�%���C��+A��0��1����v���<�]��:V�A~�����)�d`���7˲^�����h�t[�	��/��V�Km��?x�~'�e?hCùL�4�<r�fq�F��a��!E�C�b��o�7�Hὰ�L�=aڕ1k��հ��
�6�0�YGǢ��~�p��,)�)q�`��پ��{c�C|�	*��ߨoH������9ĸ#1���r�ކvC��*�K�`����n8/�zP5$p×fhs�Rj0���fm�k:�|��\��ۋX���S��L㔀�	�R נ���HF�&�>�{N|F�ڄ|����߾e ߗ�5xH>����+.�,x�e�$'�[������9�/�_�];�-�U�K�r�<�Zv�/$P}�y����`��B-®s���#z��7���]v%�V&[ ���/1*����	喽��i0�w0�K��E
��N�C�,��~�횀�����b���҂�&��r���q�D��_0�D�J���BOu6[�3tD�mإ��^W����nR�~S`2�s*,(��l4�����d�~,m�����&ER�|E,j��J�����U%z�N�{�Xշ��s?H~��>dr/��vβ��tͣ^Lʀ��� ��Zz��=ܴ6$V�z_��˾؊ʗ���#\�z9.����I�����6\��5>8{�O���0��S����H�ϵߣ���e�t��׮˽�"�\��6��	�[�ԣ1E������m����Oepx�Xk���M��A6��zM�ś�`�^[:�®����(*��.�<�E��(;��Ju�kw�۲���$zᢡD,��)|��;@=��p���	؋_b��2(<Ǝ�A��rL=�����)�56���UÍ�I��p%�z`�yI%�������womF:�+{� ��-�����\���%�vUao�Le�;�F�##�%���཈;mr���,�9�l��
�ru��}WKA2�Dg����cJ�d�۸��ȇ�Ԁu�^��.x�����Ð�~�����d�,v��c6⇫O���n��,x�i*3�ÿo>�ǔ�l�����\�
���aq�ۂWg�ד��Y5�S�4 s-��b8܄{S'h����W/�NhƎS��8�a.*������r�dSP�����y8ڇ� �M>p�lXh�g�S�0ں��B�tz��RL��73llak D {-Ejأ��#:Tn��'��G;e)��'��{u7�C�ꅐsX\f�mP�d��.��_;���R> :�%˺r����k����a�ډO��b�׆=Z��U�*�$\4/�(��hɖ�D�L�+�/���y���&�%to?�O�C��%��/��0��2#���p��&K��t�3*b*9������ˮI�.ˮ�g7�1�]�J=���$���Y�@{��]��T�>�!��I�6z�6E�p�k$��R���	����d��6��.!����?c~p�ܩp�����v��̏�H��9���:��EG�К%�B��g	6PW�$w�7������ ��p��b�w�Z7�J�e���M����W�y�����y��:�×��w���2�J<�&I�d����Z�#��+g�%�����qQ��2i�j�����W`��(2���ژ�u�l~��/u,h�`�1���8�_��ɨ`��{��W9���/�=v����l�S�i�����Y���zBl� ylջ��q��]G#a��E�h<߿癆N��l��j��0��/����XU�7r���Y�u�u�"��Gsn����b�6�V1ԈN�U��ԇ���YnA_�,�������H�u2�Y�gS��^����O�&զbI�����K"�4��NhA_���i����1�L�|���L��9#r�\�r��jZ>�W0�1��_n�����Ƙc-�M6�+�$�h���+9f����"��������x��@�wXy��!՘;h���3��ss��/��@C����ӵT<p�YStܬ�� ���mN�3��������41���x��U���Ds�>�JR����Fd�@*��6�}���D�@׿���$�Q�ҨՖ!ӕV�E�)��˫<^?[����e�K���c��@��v���W~1�ʭ�󗯑�&߆x��g��y<L�(1�'	�� �͖,G�9®����%�(t�;�>���Ǫ�I�U���v_ǜ޴��h��kٍb��ZW�m#��&������F�썹ۀ����!����M�#� �#�t{q_��x���I)�X�rAG�-G��A���f�s����N%q�2a�Kp���*2�"��Ey��~]?�)��3$�
C�EE5I(��Fu�O�o®8��)�E*��ɯȖ-�H%�ވi�����^|��/���5{�^�#8Ixיu�N�r���s>�J��E���WN7rPԗ��it���ɤ��W�B%0�e�P����� ȜY��ɠ�a�#�UV�/A��j&12-�-�⳦pk_�+]��s"[���`���%�'�7+c��%e��*��V;[E�s�w��]�`J�U��f�^�`U�	�76	Bm�X⌃�`���&��� �$Z�ٜ�N.�e�T��JE؞�-����S��2��c�<��A+�9���j�?�5�'��1<?&}� �����|��"��au���mroR~�jx0􊬛�c<�C�c���X�:�6���;{��n>�d	|f��O}��7#&_5�w]wQ���QL�y�-+���+���/���bUtT��V&/�_�OSᆁ�a��5�eߊQ\�h�_4+�,Oxȼ <�(u�E�kx <�T��"����{h@�F�D�S��u����=׿Ζ��cz�քg�[*��.�Ǵg�GD��3����e���޾��]�~x�쌚�R�e%I���Kd�!����_�]0#�H';���Ld���&M�_�,�X�z�1==[lp�T_�G�Fh�M��C��G�s�F��i܅J	r�m\�.�W��'�ξZ�͵�_|��R��l)��Ƣ_� ����Ȱ^���;6�׶��׊5Z+��׬<������Tl4Q�a��ܟ���**fF�aT�D���c�u�_f�:�B�?8m{[������T�#�6��@��E -�m	���s�d���T�1V��{vބ�6nxbؿE�L8��s��jAF.A��
 ܑvw��r�M#6h*bL���pm`��mm��Yw��w�u�]���#!�D�B�����	��p�Q��m�?r��k �`icݬt#�.�/��͎�z�}�`���J�/�.�#/s}\�gN��:��<Hq�9
���ؿ��}'�]�@f�i��������&�R��;�؞�Ța�	�і��cpE��s��S�,�^�����׮����cx����.tu���s7�<�G[Fe#�?���W�jE���T�%���'�E5�BVmS��y k��u#
F�}��j���'��DJ�[ʶ:\H���WV�d����[�@�3�z�G�In(���"��$/M�f�V6��jt�O� 	�G>Xe���YfP�L���ߋ�ݧoI�	�����l$��XH�GR��э}�u|P���>v�TZ��B{�'[8���S��I��X1���w`+�6�@h�H5��	1�d��[W`l6���{N��u��#�A ��Y���ԋ4Fs�I�V��[\�	�] ���3��[��.<�R����Ȱ�#>�'��d튢E��m&i�;�� �߾�M���;
�!��وr�4qy�^W��l_v0C�Lt����Қj� l�B��07[�����z��>$C���|C�P_ξ�b�~�A�S��I,���dB��ӳ��b�]6K�/�"���_��j���n�f�F<��=�-�r"����sն���?P���	��{��D�C.��:X���x��N4u����H4I9p�A�ҿ�S����ҧ-��?L9Q��o��"�ޖ�f�[����]��s�c��1M�O��b#���a��{�_���lD��O&H���=&\B�o�eT<e^dId1��QN\�3����b|�ՎOC\��m�M�*ےx�F��F�S5*i�ː�Wd�~�AV�Ɓ`��",��y�0Ŭ�G�� ��t�y~�D�R�<����}��܃�:�"����Ж�Z�~�1�
����j��CV*z��M+'Ҩ�M��<1�����/�>��?�3Ҿ_\Jtf�^�:��]�O%V]1N�U)�ܰ9�:��	�v��L����BP���<q�����MZ�Alኧ�/��RGa�כq�����/C�[�n��'����NV�.�=�E�To"{ �o�D8``l��� Ym�9�����ܒ�cf��m��n�-�0��Di�Ϡ�{���uhl�ɪs�-�9���� Sq�VD�8A���X�'�b1�W+��p�v�z0�u�x����97-�T�X�[ >f,hf��*өrJ��JVBVAYU�cr�S��>'UQ�*�_��P��f�㢙����*m;.ZM
&�Vx�L�*S.T���g�3�GeS�%��2>��z�P_�r�Q�5Y�����_��4��K�]t�/��_��鈱�%�8��}�0��.\y>���gQK���F�m謌�W1��^�S|%JK�������P�􀛭|�1������;�J���Oofy���!������I��?2��if3P�8��b;���h_��>5�2�{$�]�׿�J!������~���ՉÜ,S0=17|�:�5����B-p�2��_$0j����"w}�cǪJ�H��x��H}#m�Ǻ��b����6U�={�T���� ʒ�8�OsA�x��˯���~dbc���p]����'�S�̷�C�m�9������{9�;2���بߧ�ԱHp�8�[�)T��R
�ɟ��`��q ̠��Y��,�0�n�C7�ٮ)�D7�I���¡��Vq�4��E��~�-����/�٪�H"HG�[��dԚո�w�3S)�;N�CkSV�	ϼS�ʀ��!Ո�'D��ι
Cօ�e�G:�O'|�5l��D�����p��\;����Ǒ- ���ڑ�]T-�g	��y��n��]v�N��S��)����ѕ�:Њ ��~���U�����զ��Zo�c��z��<ئt�2X����F1b�Qj���6��6n:y���j��n�n���]Ň�oϋ�l1�C��ӷ��0�(��oJX��Me,�#�Q�cʝ�e��@��i�~WGՕ8p�6ϷZ��b�$�h�_y�	|����6m�&�r�lt�o���I��g��Z@�7��|�%�oQ�C���ٮ�8����r´�1��O�G��&X�Q��y��u:w#�Y��J���MQ�Љ?�u�u r~�8�`z�އ�e�gF�H5>�hk�հ��H�8��>�_ώ};;�w3����9�Q�`�䤎���<n�+����F���=P�5�LǨJ��e����2R������_i�j���������v���5��TO����������n�h6��R
�BB��-G��@.D�wa����Z"~�:�*+�_j"$"���J��%�z4Y��:$_�jDa)���\k�� u�!���p��jał����w��>:H�_�A
�c�ΜF=���W
�t�ʇ����vB�r�|$����ԁI���P��� �s�PQCſy����kT�X4#�{&�7��(�'Q֜_CK���#�!lS�Z�e+򸡔�L��1$���.E�G�7�F�x�
g�Z;c��	JFu`ݴ��ÖvcN�%�F�)42�ծ�#��#���i���\���S���|�G��M��$gVң3]�5�W���0� �D����C��Hk����I'�h1K �d�?]ȇ���}�����^�7�3�\W��c��*�Dڨ6�tA/٧K��TW�Ӱ۷Kcw'�xG�˚ivJ��Ȁsx��>!D^G����
�{:B�ٝCب�2Vd�]Fv��l�t�Wn��v�T]Z��\L�*	������o�=�qF��U�!�)�pZC�B/Q��śP�?�ӡU���;��P�{CC'_�����h��v
� n7�]6��'�6��k/�Tc�z#��w�=��Fa/�w��2T���f��{�2�m�q��><G���V�)#~�jrȮ7�]sE.����Lq|^�3:��Uʢ���}��+��hT�LP	=4t��{�Ry@i�9QP�� #��_��Fc��۫��8���ҩFt��֥g��P��>h�֧|�ld�Z����Jc�F�[��Z��WA�e�n�GsJ�/b�]$RD�@���CJPu���f����F��#����0������P��L���Xb�&5ԯ�
��u�s�1X��91rN�Rf����q��A�ٞCQ+1p2�&�W��ECq(�"z7�@Z>]>�+4��.��p��s�W�����	II �%FT�x�:��8�Ui����F�� @B��������Gaa��X��`�	�O��Ќ�&�Mr�+[. �7�G����}�\`Xp'��"-�H
,|���,�K^W�`�&�G�U@�.6`�	�-��hT@`�ݝ�m �,\+�Zz�g��u��g��>�>3�}������ꊈ��y�%��3%�c���7�w�@�r�xde�U�̫O��'��*'������݀ꣃW�KN�)'`n�
ͨ'6K�J~� ����>P��RU{E�O�2�s�v��5�a�F$�KΩ��i����0�5����|`���<�E�=���sw�uYE����E�g�;f�K�d�U`�Ƕ{�9v�u�j��Í�5pͧ�1:�ˢ��>P��-zq*�*eЅ㌪"�~޺�S$����{�"���3�fV��$��m��4Tm톮��8N�{'s�6P͓F>{p�/.���ف�ν�5��=���/F7?ޡ1��`�l�ƻ�AZ�y1��d�\*ů_�0S, �P1"EG��>eb�;b���)z�|K�2��H�N8�[{�_cb�E)�c����8=[ ��(�XԲ�x	�ްR�0ǚ���Ȉ��)��R�ܗ�>>��G�N�P,�ai.�I�u�=�����4\���e�u�zB���23I6��cq���elBY���ea��:����)G�-]�W���)��gcͧFSy4ez�z�=Lk��+�y����mɫ�}�>5Uc�I��#��nSO�����5+��]wU�@��ZɆ����x7�馓��Q����2%�3)È�CոRj��.A�?���0���X��0/�Wfd<I�c,�棑�oA�~9�md���|-.���(��\o��b�����tWQ(Fs2p���Z�&���Qr�d,p>h.E�T.he־8U��`Voq�"��6�X��= �F�G�i�,�>��|���W�눶;��x��y�<#���c����K*�5�+QP�?�X��*T�
���7o ���Z�_;#��T��v>�x=��CRv�t�]?~�e]��Xg�h�E����n.d��;b���'�jO<���i�A�{�o�7�*2�a��ٞ�����!�����~wJ�jN��!'�;����G�1��O2�� ��DM$�Dq��n���`��m&��Ǒ���c�$�`|taXz9�$p�B��1����/�؉ +{�k��$$�L� �����eRD��Q�$��g��2��:
�`��T>�B���=�tD���`K����Y@����iN�vp�� �qf�"��

!Az�EɊ�'��&�.+�z�7��n�$�̛u#6���%|#���A5MMT��ȰB5�>�Л�I���.J��Q&�F��x�(# ���]���H�%���hg��~�����V���]��L��Q�{X[��$�&��$�ζ�vV	�*|*Y���γP�B~ϟ����&)U~2
ͪ�ogt0�"#�WL$.νGy,by���|7��o�-K�Cޝ ��bc�V��l��߄��"����[�:�pFXm�c�0�.N�.i)���� ��R���YMC_�N���B1"����V�P����`� �k�F�����"
`�31�=�g���C]7�Mw��N��� �bb��*�6zY� ���C�U�������7��_�H!c�,
qˑ�w�G�6A���88��N�ܕ  ����ՖX��w<%S�B���[d�JN�}�;�G����� �Ĵmo�szυټ��a�@�]8K�|��b��\��6ܝO�q9Flk$z��s�v�zꑥ��KrOQ����=l�T~��Cꡰ��d��&n��_��G]�K)[�uS�l�)� 0�|D�
����\+���ۜq�#���ЮQ#J
��L�r���[:�t�+ZZ�6r��^ZK�ֻ�?�I���*�6�
:ǃY;)�^�y� ���bE��ٔ�>��8i����66��8�B���El��Z��6�E��A��d���������'�@�v���(��`����~�A�f��>�)_>����ڴ2Q�VH�����>�SvT��\���g�Z-!'K�z%٢�dڬe򔵌"v�o</�!T�Dz��ϭT��Jq��PIr��k�M��W8��E0{U�f�	�5�	u�����X���W�Z��
X?*�����vs��i���GB �,|$4J�J\o���e}��`	��w5��rT��PDв��2K��K��(Ҙ�`��<K��ŝ)Wf��r��fR z.m��ި�s�
f�Xl�I��&L�*3��u~Ie4ﵗ9�f��\Y��r�qÏ�*�D	��c�SS���n�W�ѵ��o���dUv��^Mi��y�΄;��1�(G0Wr�y��p�P��g0u�۸䑶;��=y��a,ѧT�� ӯ5�6��@S��c]��ά�Gq���y�աhE�$��_��/x�*�-ڌv����I�Z}f�x����,��3�������"��oA]����t��k9ܯöx�J�SͮH�VZJ��d�?7������Z����C����.�4���d�;q��p_*2�b��<��nku��B8ڀ_W6�lǟ� ڡU��A}�Й.U$VW��HY�Q��x��$��x�ܵ��#��"�g�jKYg"bN����S��ꅷWt����ǝ��"����&��g�ͱ��(A�#ƿ��1.k@D�d�&l(y/ ]:�w+�_-��r ���j�g�ƶ�e�e�a�!��'
k�'���d�CCC�6�厥�;�)��t�������$m��oY���#�2/�� 1L�[�^�VDn~����]F���b�a6�$��L`n��t`؞gaY�:C(���1*Y���P�X�r�v�c`������A;������C��۽V��43���	u���T��r驁�����#IgHԼW'H�O��Z�*S�����ս�`�6�O�d��JH�4�n'ΰ���f��Ҽ�i���лSW&�2�L�?�����ҝ/<���C�<c��K�c�����R3}��Ӽ>�ZB��gS���s�+�)�/:n{d�=j	�3��zԚ��ኻ����8���A�f�J���L^)��
zL�o� �k�t���̎��pdP��w�����w�M��:���`�JC��/-Z�@-�-6��/L�f�n�VW�e����@���v'�y�N2o[7	�MaX꽐߲�37���u��d�u����T�(vtӷ�B�j3��s�=�"8ѐ�o��2\�C>>\��N�~踦�&�h�E��(H˲\p]ڞ�&�r�5�ĵͤw-w�:�'%���K�A!��ƽ���$�p�e)�iw��C��8���tH_�!��N������.'@eQs�#1�o�Z�vw��/�������1��3�a&Y����ܶ�%0��������*56����\�_>}wA
�M�u����|�)$��M���i�j�Ն)��P|�E����n�޹@Y�×`@�#�1�A0'���J��*�k� ������{	}0�0�O$�I��t�g�`LV�|�y)��
7�l��[i8�m�B�uYi�n�P疧����ں�MY�0K���ҭ�=�s!����
�ȓ	�Pңs>u��`��kN���̾rX���˺~b������#�[���|o��l�����%%��������9����dt�:�P�/�f�@\e	��*Ɖg�#�ŉ����Ø�M/J�on��m|�������,��j��a�#���i�`:0���I�)t��8wr�xmi1�&��	�b��a�#8����@�xy�@�9h���,���\��eK�!�*_�\(!������� �]2�d2
��y�����UE��ծ�;����A|�3*ݗ�Qqd5���"C���Z8�&�����IX)�=���`hb�T������釶�~�p0��"���P�W9ǝ!� ML9jN'����`D�._�6����1o�������ʉ�����$���\���7M���~V��X��A�{C9� �?B'��F:�Ѳĥ�lǵ���c&F?�*]�Ԟ��p=F�71���i���\�ʥ1B���$(���UǺR㷐"��3�Tr���Ux?�Te8��uE���öQ@`S�{�oSRG�����Z� i�?G/\�|��F��˴�"��b����d�/��:�[���+���gX��Ӱ7L�0���^i�2������	�k��\~;�wvNv�����2���������}��qP����U��#-�q����d�]Qͣ�N6�'Aka�i<X�����h�Lou�%�`��
N�"'��O�s}E>eS �oV2L���キ�d�x� JU�E�U��$�`┡(���	V��࿿���m�;�����$��n�Q�ځfsP^h�T�;�*I 6!�/���p^�r�JԾ��
�(d}��'s[���Hķ�=
СN�s���d�"���s��#�J;Q�R��j<B���iu!}?��׷����:+D����9��I؛���ÆB�(���*���mR�je"9��χ�9!�$<V����a	A�.�C(^-g�4<�d-z�j'�A:Bg��E�W�����u|�z��`�lG+��4�t���k9�����y�yL�e#�x)���
�ϩ���;6>՗ �	^�P��z (���]h�?�Lܑ5QGQ�ζІb�X!״�3�3C�5��-�T��h��^��II����fZ*�/��2ч����I]bXq�z�7�5/� ~�Ma�sv����t%y��3u��2���;#�K�*�Yt1앭��9�� M�@���c���s1����<���m���Tj$�����9��'�q
j����P�W����T��"�&k�K�1�ʌ��'k�Xa�˔z��ż�ɨ+c��: R0hl�LȦg�_�JO���q8�1����G��h��+����_"_���k͹���ò�ISX�3��3$:&V<��
C'��z��^K��S�e���<M���E�����B�N⩊������ȿ�_�j"ˌv�%6 K���#bS��;��k�~6:�w(��XO��~�u6�d(��`7W�á��U=\�;�.$W�0�M�I�а=JfB��iR�-�A4�(�'�o,�9mov�/�c�2��+��l��s�(�e~$��N��dum$i�fd�*W�������#�^	���Hi,WL��!m~kN�i��|xRj�~�/:IN往�*QVӑA�"eӨ)��$��Z���ri�N�GJ�a�A�Tẁ\o�g��d�D���92A�sX�+���A��P�����R.&?�/p��B������lL=Zʷ�{.a3�C���Q�tai�G������ �RB��#pqu��H�F��nk�ub�6� �����^�X=��K�9XжFE���	2�TǽH�W�pպL�p�uer�ڰe�$�$*�G/�-0�4F��s���KGG�w��p��W�,Gt�.
~ۉ���D�ٍ�z�p�%��HYن���R�R,���� sС���g"�8�]�r�h�K�����񟣆�4���Ԋ\#��+��cJuA[K�DH�9+6Y��.BH�_�z�ڥ4�
��?97�J	���D5P����~���Ur�p�ȝ�������qy�hb)�I��H�F`g��7�_�9eg-
T�1�=�;-�-z�c��%��y���E�׉R�^������:R{��n�!�sV^uS�l�%�M�ś�lf���Hw�]���yQ�
gΥ
9�Py� ��9����G.DvEh���ҳ̈�d�+%�I��AHP|Y��sm�6�P�UG4ǌ��8�Y]��Y3��l�{�kItő�ja(��"f�݃iK��Dg�����޺�	�}�t�5u�Mѕ��7	�� �!��ű�N����{\�Mn���ލ���wMs�^כ�dw@%/�`�̅��p��X,� %h�[�����:*�f�-��rb���y)&MTNggL>�XQu?�Ee����jD�笪�]Mt"����/kSc��&Վ�#s��0QIO�δ4q/���a �,����:'E3`�dx��f���)�Д�hj�z�_��WhO�2�����Q&� y%�RI��˚E��ڴ�jBC�S+4����^s�ȃvk�>C�,"��ʊ0j�xE��7�y��M_�ro+���{��M�������1HvoB�G�m-5�=�Q8�
����mQ!��I�SX�l�W� j���"͍�68+�Hq�w��ih�A	��"���s$���G�.ӣl0d1�r�g�L�j��l��9��uߥ���_4j�m�E�j��|�
�!Z|�z3�Bf	�V��u�n��vP��s^�N �տkX����"q)?xfKK�,����,�p���G�g�������.P�	���(	�e7���`�I���Q�0$`�%5�����B䧚տ�m�{m��)��0��t�𙟼+j��	M�/�'9R�?I>j�`_+E
��qL{?ϥKW�vA�p��ژN� t��8%e[�-��+���}/!��;]�;�m����^���2���z�mK&�P�c�UFYƵXt�͵Q l�|%Й��-�{���T�O<wsV<���@i�Ņ����%�Ѥ7��k�
{�u�5UҚ�0T�l������¦쯾�P	_����\�E��[��g̚���z{���m�����h�g�?�7�����Ga�x�w�n�C��Bt\��^ml�������}���\,`�e��R��8�βZ��]��ǣ�\&�P"�SR�Z<� �:�>Ej��pˤ0xw�љ8d@��o�?����ײ�$PP6�X���[�w��u�
��e��e�҅�'.�0��z`�R����	�U�lR.��B��`g��X7��fU��E)�( ��:�[�8�Q���p�Z�6�3+L.�j!:��J�6��I�����t��>D��q�Pvqo
j ={�.4��l�J.i#|z���!���w����r�D�����$���qF^ �=;��[��E%�h�X.0}��?��ä��^J:��2rǗ���X��
���e��<Mp]G��6�/��T�E�V������S`NpC	-d��֎G= {��������T@��2�Khw��
���$�v��Id3+���������0�_ik�2���1ɮ�!(�)��cθ����ў��*?˪ 1�#����q�W���;JF����L��Ҵ��AOt��0*u��양\��ZvgR�MA��JQ $�����f���u  �
f��v&��	Y &@����5ن����r�m�&�!'�y6t��
q|��o"��d�%=T��҂��|�^��mm�Z˃�R�=#��N�����-�T®!K�:m�z�!{�8Ȗْ���-�G�Q"a�+��R��\����GR9.gy��"a�3�[����UW$`Hjʳ/D[�/�s�ɿ��c������:dg��8P�m=)�F�e���WLo��m��E`��8 U�hƼ�t�"@T4��{n}!�TT�=�̪Q3��aO��&}>����:�a��ϬT{�c�1<�;G����F�nyg��=� �Q�}���Fa�W���d��g8=7g�JV�[�9��9��ۊ2^*o؝�a>����G0�M:Ti[�'��'U%���ޥ�b"w K��(���.�̓.��^��X�сR��{�ki��-S�<%̜����Lq����U����~@H�g�� ��p�;��@�}��z[j�y���[�q]wyT��Ls���a�r�و��t a����`�dw~d��:��.d�j[w �C,�է��9�����hI˓Qơm����
߸y4�R�A���D�f�YB{��Y:T��rT�ҽ%@�������	9��O��Ad���m����ƑW��@����!�`��{���?Q��ޮ`�%n��~���f�����5�CzsI�#�^�G��a��:B� ������nYݔ���.��fu�U���=����]�ч���|�;�+���ZIm�+�Le��4̀:���;�-�3��A�(��7��8�zN)Oȯ5@���%)$'���k�81�'4]0��	)T֢<93�_�ۄ�J8pBcgJ0���ܧ @��
BamN���7ny�H�����E�non���bj��@&A&Q7hV=m�iȪM�|��:����;�_٢nكe3z�V�<��a�~i�<T6��K�:w ,����鮽�2I[�����I��=�Gh��l��-F$���,����e&7B��Xn7�m@����6u0��_��jŏo�d�g�w��V�A�.�v'fF����(pY_�C�xi��xr��U��
���B�r�GM��z`��i)�FJ�4(ވ�"&�~��"�x����ܟr�N���)�.	�?f[��o��F�MyZ�ۃb���t=.���_���� MyV�N.�%�MZ<��g|����'?d��Q��6P����o��2"���|���!�.���h��\I߸WJ�U]r�j��g��䧔j�=��2�������!a��t�o��l�l�k�dp-<e���J;pp�P�R{rIC_�q�e2�@��>�6,�M'ξ}��j�yP�Rߵ��I"�0Q,f�d_tD���<g��1:7W �u퓤���h��`�?@��=UK�����E�`ʫ	m����6�ǟ�ĭܲ�ў�!)z����0�p�ꈕBB\�s0K����d��㠑��}�̽�Y��Ŵ�r�T�x�T4�XX.Œ.�z��x��S}�%(�BPN��om��I�e�S���@���oŋ�}���cBZ@a8M�l젙l��5��,o���������ĩ|�L�!�j���GV��������8)w�
T�a*何�i��<�<��j��';2�����	mXꟿ;ŗ
�j�@8ip� ��7e	�����$���<Խ�����(��'�=lo�Tu��Ջы�����	8�GTkk�o��o�&�cSb����4����u�"d�4��+��bϠU��8}����f0��b�����������f��Q��.6�`���xhc$[x��V�'
�,�yDw��h��i{�K(г�;6�^�@�/��yq��*[z9ǦY,\�{��>��z�u�0\6H��]6?L˩��Y��ư�I_�L�B�	h�/x�V����Y�t��Ҡ��$M&�^F-Y�X�����en	�^$K�2�)é���~�mh�<�Z��}���y|�U�s��!��R������QUO*���ƭ�`q�>7��t4�g�U#�9}��2�,��pFV+��2KW
*��
�-�����1��t,�	,����wq�@IE�ds8mg��9(�+���(����
e?r�����"<�̎re���a+�������½;<�����G(>E���G��3����[_9K�e���r�[(��I*ܭ%i�K�d�q�/=L��E�u'xqy$���c�`�x�"3Fnx�I��{UE6RA�'��$��|�.$�z�x�b ��9��x�)��9����	�3{���:%���O�u�Sƥ��pb�9��l�0i���x�8�ջW`�_�=��+Q��P���x�%��c�/<���gIO���vL��<�E���]�����F����6��͙4��*I���A��|���Ed����}�*B���o�?��!�M+Q7(0�e{z��O��c�`��E5��)�;�� �C(���m~�9���g�Y�,����.ˍɳ!E������x�y����$\˰�>��Bw��Ǔ�&�{�#��N(�0�c�`�՝WdU<Y�p,�K2��#x��\;Q��f���TV�ZN]߻l�Ԭ&~%�[{"}~�����>�B�k�oq}���D	А���ŋ�(l{���?�a6��HHy/XpTHX"��8gP/�і��U�����Z�.�x�~����uL ���E���.��������'<&Zvl�b�R*ȁv��;(��}���O�u�������r8T��~��I�>s�IJw�����!�[�P���պ	�u�[���M���	F����DE��7�&Q7D�������y��$��_��B�ٖ�Bl�s��6�8�|P,�72�B@����n��H�f��ɮ�$f�*#��p�*�- �?��.~�����z���e�:!E��%�A�$�̐��4c�6w���������iX6u��3�]�o�i�8c[xk��Fi���g8y�^���A:<3�^�ԭ��2�hG~�HlŚ�r����Ñ��T�4���wH���&�	����PŘ�Z���7�๾��><akhu����9�@.>�Bz�%j0��ѕ�?�xP�i8�~5��\;���}A��ߵ�,�Ch�_Cx67>E�6(��eb�D����C~��
]G��Ko�
�g���5���2��\��7���O�xs�ce��G�GZ+�}	H<�r �ޡ�~|h�#W�~��V4�-׬�gZ����|.<���t�d��\��|:5b��H�='�g�T���|̻����Q$$���'U�*��F�Ub*ؤIqKE&<̎�	� ����6�#�ҵ緌ݪ&��=�X\l;H��r��hmƹ|�)��6󙁾ܱ����$!����#�Bn��l��t'���@Zx�=���M���䦲�l6"0~w����BNy&�L��?�kǲÅ%�y�m?���\�"R'����֒\��Tɸ����H*Q?x�=���3y��C&W�k��~���g��h�����&�7����[�-���s��|��׫��ɋQ1r��h �D�nҨO��CF}UiSJ�Q�o�Y���L���\�����!���B	O�O����ůu6,M~�F�P�ϥ���w�P<��9�&}�����Ҍ4��x�����}�ނn�� ���݈M��d9�9��П�Ilb�$�ҵ��9DG+R�y��T��^���u=��S-/��\ж�"5�����uf����a�"�1 ��&ܭ}�TŋLAE32��-wp�G�4��aWq7Y�K%�?���c�ǅ����i�09�����y�,���a|��O�b��}Τ 5�R��+����{F�h�� �drw����ӫ0�E�L7�::*�R[�FT�aM��x>6��)y/�5<";YL���<�X��ք�
(Y�<��^׾T.e�p9/��R�9e��ܱ]]�l�tZU#�v����uvt%`�|%"��Ac��Jc�B��޼_�O-i���ݜ���Հ���̊ߠ+���������4Þ�[�w�H�S��֧g\�y��Z���m� ���Vd��ɰu�;)'�)���Z��jlˊ i�W�tB�}�ɤ~SvZp�CF�N]��z�/	���؎�\gm]7��I��2���#� O:� `��іk���v�k)x�ǅ���<9�Jڥs���'̽BƢ#B��q����Qu�2(|l���+�߿m�A�,W��MX_���C�n����L�ߟ�>�DȺ,0&�2HO:��3�7�<jl
$�wK�^]8=���8Y.�1��܂RظK�r�762N�r�)�[���x�)��k���]��/��}E	��V�ƿ�Z�6!�y
G�a�|��#�]�'Ǹ	�cͱ�|t��v���D�®Y;��r�V_�ړ��Vt�X��	��+���,`x(S�*Ζ�\Hg����H��Zo��b,[=}���S��a�����:��A_�:����wM/bMy��h��޾c�����C'P�?AIxA��Y㕶���n�0��+�<epo��'
�!]H�VO.���h�7�p�6��^|�F��*%l�ў�	�RF�������X���ip�����:j��>2�<mh�cS�t9��A�y�3R�~���fϻ��"�H/P��x�4���b,d�~�+V�O�j5�t1�ve:�u���s1˄�EXĢ�SQ��a�}PSۢ�'��Y ��N��Ƀ�]n~^5����`����CB?�t�񃕔�<P��<ЬɌ�ڠK A�����3�!�9�����K��7�	+�WQpA�ks�!06~Tθ�9�aֺ����c_��?�+�1O�@�o����^:�Ge�
��Di��i��MW_��[ c����LL8�	������:/�D��;��Z d-鱓��*��frcRv�;PȫY���HmUqg#��\E�膏ɔ7��uF6�G�yCطqxҹn���d�l�u�V��I�f��ߥ%�G�+�x<�[KS�}��S�����U= �� Pv�7���m~܀��r���)���^krj������U[�Ru�����UT��s"��_�ur-�w�@�����=ҙ9���	�m��4'7ƐK���d����V����?"A���;nl�Ɏ��
]:[
���tw��f�}�D\V�@�q��1�Ƀ���ʵE>�ЄIӲŸ���W]�,7�RC������X3-��,|���ڣ�(w#n���r �=є���, �]��ɀ�#����>� p3��O~�9�csY�u`(��B�,wI�\f�	�fJ�~?@����H4WH�2���@V^Aq �@���~��t�������,�$!�O�������\�t>�Q�m��� ��Ά������K�	Z����Y�e�Z).���ʚ��M��._8����g�b�M�]�WS��`M�[�
Ud&�����`������[a)��fh�g�!<�:�1�Y�-����(@ ����tp2���:V`��;@�k�*��W�p��BW5���3_�Q��#�kf�t�mäV�}���q#	��\�ښG��1�H�v��VW��I*���Q%���"���0TRy�3i<��"Ǉ�K���=\�|���y���$tꠕ�nx��&���R�Dg�.��k
˶ �ڍ�\.p���oY&�KڰU��gl�] -�]�\RV�)�PC�����8�J���]/�|�;b��+��1�꧈�x9�\P �hn�T�)\&"|��r�'�1S��p�l�l�+�%b�e�/�ES�d���^�4J� |(���?S�`�,L�}E�*Z��V�u�?��4=�ڭ�y��p�/�;T��x_j��|`��L�Zn��W������	ĵ&�2�,�-%�Ksڶ��zpB�CN������GF� $�p�0�}��[zEN.�����׃��������Lk����
���zȇ�	��E�,�}�	��д"6k��"ׂ:}^'%	�4w����V�R�l�p��Ӣ�������_�������#
��}�aSfU���.'�d�b� ��D���!o�mB��~i/ 
�&p�
V��Z�bV�E�?�I�'j��K�w����J;	1���N_�ʨHnY�Zv��!ZD���h��P�1�Sh>&՘��v)��	���������UMvÞ ��G�d�z�{����1�e�����+7{j@\șS&����b� �1E*�2dҌľ���c쌼�b<�=@�jP{�)>��@
�I��3�23p��=4<�	E�S�EG^1��a�Qǆ���{<4�)���\*��G�@_B�7�=1w2�3܁m��rJ�`^�y:޸�r`�s���s��1ه�kk���BtɅ��f�F��8ǃ�S��e0ڋ����CԬ!�ցH!�\[�of����)t��I:�w6�8�.,�j��Nߟ$��0��4�K��f���cpQ�bD��.��=|'~x02�����]���T���2��g������P&��yz׿e�j>��ĩ?�y�C����e#��*����t������mP�/7�2���Y��M��a@-/�d!��e�Ǒer¹N[�Hѡʢ��d#�ܦ�Y&���R��ɎI�e��=�t���H���D�����	4�k�J�[������X���〶��y�^}E�W���f��\�	�ET����Y)arU�A7��*7��
��S�MkX�X��� ���p)KOHB]�|�ch��|DV�Ҭ�D��	~L�EZ�r�X�Cz_x�{�h-���$oxԜ�c�Q�J���m�_�!+�"ǲ�׿0~7�'`�A��!�Գ��;G�Z��9γ�0U�� %�&H.z
gU��5��x�d�VÃ�0w���ᘶ�7v0�)�H<R��3���q�4�+��w�GIC�C�[J�[����[��q6ώ�	04�A��:��ޫ�M�kNw�����&ǫ:���v�o0���rY�:>`�]��+�1�,�</��&���\���̍���-��;�E	;�.��o\�|6��4i1E�-1k �m��7�?%����_#��.��J��(Z>�E�guZPtLA`�/��L�+_�\߱\�͆��@e^9�4����V�1�(�`a=O�h�iq�?�
{�s� :��y]�J�a���X�&�%���=��4���W@j��۩��|���C�t"�����*��
�Eeȁ���B
{(�6��	�M:c*:O�iY�]=�yw���F �f��,(R���dF�@�oo-�"����j�S�_���Rf�U�%�� �H��
��# ���S|�<��Y�w^%c�V��ӰċRj�Kˣ%�R����L-�7��݆����.�U�@tk���RkTI��4W�'�4���֊32�߸-���M$ajK�p-|��G2
��t�+�+��mY^R���Q���*�Q��_>����1�ٓ~�Bŉe�$�t�bV��mQN�7���,��êwfM@�w�N!���!&���,��I�i�s�
4ӖU�Ț��3��m�F��*ߚA'�^�I�&8�ջ�[�x5yg��x;W���YjA��B���g�?w�{@�M�!X 쳐б��19�_c�>�.�ܗ��i~���wD��d�)xc�v~�C�������J�6��������q��.�)��X��I������@` ���/� F:�9� �3K����d�/�\�|�nY:@Ҙ%b�Ӗ�7�_E
�1p�����5b��.�Q*N���7���"�Κv��Ð�R�>g�����B6���#vpׅ?�/�Y�������o��K�^E��W��S��M�ʵ�9�,���6ىǰ*���"�L�3�Vװ���g����j�>MJ���</� ��]]Zz�+Di�>�f��C'{��Z��j�4L��ȶ�Z�rP_�G����K���K�h��G!�г��t�"8\(�(V�h���-��K�f&mǖ��\�ﱠ�ED`N��'�[�M#1d�C��܄sȍyO���)�����o���$��Q.�B�5��U��럪,���^R�RfD�"$�Y�%��K��H�'��I%(ĵ"<�wu��{���o=��zT���������6��
(+��6l�D>~+�����"��uXe��^q"�([u�J��e^��8����Fx�[��P�JL��*�8�8����v�LU�vY�#��{��ǵv4�yW��}<���N}ӓ�/f+�/L�����D�9"ǁ�����Џ2Ԅ��WK���L��|�}�&�4*�t�>nv~uu$#��Q���P:<���(�"�p�2��Y��PQ	k�'�+8����������*��|��
g�w��y���k~�X�U)l"�� t��lޒ0$�3M�o����f}{Y�Dl
0M�Pf8�Ia�
�Og%+��Ct�ӛ�[i��lݗ�r��5b�g6���Y��U��zq����%����A��U:��E*m��P�����}}a��j�g��l�Zh��e8
������^e��_���~=.Il��ɴ��	a�W5�L�S�'R�}���c�"�r�}<�$�ۢ�SϹf�8��E�k����HVW5-%��r�� ��T�߁�ƛ�9��2�4��_�žR�X�[��s�jw��$���H/�6C���
U	H���W8{&�gkn���W�|�J�w�}�/�� � �G���O(���8�����n?
�O?����.CT�y8����8�M�E��Y�@@�m��\�P;������;2;��)+@�0+�{��I*$W�������;���߄��ސ �8����d�|�PuE��D1%��H|^:�8ډ���}SFe	��a��փ��?.{σ8��뵓�S�4����[�?�y�:T}���	r�:2�N�*Jl���k�i���PYr�Ϭ���R������!s��V~`Ϸ��`�@�8!ac|�5��8t�� ��E^�d��@g��܁9σ?��n��1,�,��m�w(6޹�7Κk���^,9����-e vxȐ�� 
�
>���"�zl�1���?��"��"+y���#�l4�0�y��gi�|�xH)��z# H�/�3�m�7~������km�<���|��k�K	|z�X���-S��)2&s���#��C��������[V�K�ϳ�.'�\��"�3�H�ǃ��S���#�2��sc	QG���vW_�Gf��@Iê����� �~WB�-���Y�VA��Xc5��5���n��t%kV�p��#�͉���$���Î��0��O��af�k$�r,�J#����É��D�4�oflp�T R3K��(��b}��q��P��eB9E�fX��n8��'sL�.��)���0w$Z�yA׺�x�!��%_"�����dM�<D�쇕��j�.T<ߤ��c�T���㩆/����V�&��8N��t��g�X8���z#4�	|�p��^�_"�p�QVW�a�	.A�^!� #E��9���%�����.Z��|/��&�CBP���(��/��s��Ay:�z�Auz�UB(<�����4�(ɥ<���y�e��� UW�(����I5��R��yO��i?}?W/e��������GUD˽��{�Mܣ�l�<-��W&�r&hr���}�y����%�>G�>}@_�\J6�:��^��+��L~-3�����6N�+9��]�5Sk��>Ism^*T>�^��*9
o���4ZL%��{6jka�7��m�%%Q�y��V{S0`m�$�����T�^8�x(]�K�������t�Aܶ>�E q6�ᘏ���t4p������'	nF�s�����m���^:,�e�W�[C"���fs ��oጛ�#��.��<D�i���i��m�����!m���$��0�n1
�&�uBg~OW���d��N�m�w���re�=�k@��˗��u22�_
OڟJ���6%8�6,>�l1뜹-�?s</������T�ӑ�ya�e/	�ҕ!�:��]�p1;x���ІOX�y��e+kH_���ޟ�}��Կ�T .\�S��"�Hd��z6�J�����L�Q��&v2䐎���쌩��u��cˮ����-xQ��7S����d�����2�ϲ�=��C�;�����u"��(9��(ȟ�hhhO�.�Ze�z�M�M]��&#�;�Omeo�ɘK����♪�&בy[���	J�>�+'8܋��nc�]\��a'�h�R� $�%oBJRÖ�x�<x���rj����r;�%���c0�=����)��T��t��<�L�a1q�1E�ڇ�M=�y;�b:�0�;k	|��-c�VV���^�Ps1*ö�t�G�$���ѹ��\oe)Zj_�z�o���P`s�#�,�[ȡ����I�o��-n��{;�6��(��|CN�ē��νj;�+�U��h T�]�£s��-	ۼ9�J��K=��PYer��[Ɩ͇�n�]��K�IW��dlckc� L��f����:S��_�B-�[?-'v���}�`0I]��I�d�/�*��Sn.�BtJ(�n��yRX)����`��3sྤ���YV��/c�P����5��3���j;��9 ���
�m'��i�?�,���,���i��v�vR��[J���q���S�[��K���'�0�;
�!�z�J�u��a�*Eec�p�����Ⱞl �=Y��E�p�U�X[�m�� L���Sù��m��Bdӧ���%h h2���^u3�=�^�yw��v�U%7)�K��ZPMM*
���Τr~�*R��^fٞt#�S�@Q4%�DX� �?}��V�̙{��EW����o5�H6�+�SJ��@�q��և��Dfb��{3ΰ���哘���]��Y�P[�۸;	����*���K��Z<�캺��S��5M}�%�S�������_��$x;$6$j�T�T���k �GP*hv�&�(�(�`
��ܞ=�|��|��,���-V�-�_��=mۀ�^���͙�O/��� ��ۑ�mtPz}�.�3.�4%q}0�&�,�3���O4S�n�<���xN���#���#C�"��~���Ś8>Ӕ��]�삹�vr�C��U�T���E�κ�Q�/��}�К.#	����r.��H� Iem\]c����]��X�������^��?�qL����>y�h�+�Zoh>X��`�Z��-���_���Yv�ZfS�����-����y�Y��mU7��id�Q��Qf_;uY���m���M\&\��}��yU�Ҏ5{�����/T^���E22˜i�Q]Q܆�ž�
�����,�F�A �^��w�y�q���*`�/0o����b��ƥH��i&�����8�>IQ���ɲ9'��Y�v��h�(8X�����2�N�u�6�D��.�� ����cb;b8u���"f�j�^��Ĝj�XQ,��\�����s��*"���yV
%&�	=��9Y���ձ�W�����cغ��g���i��r���L�t萅�� �JQ
�Ț�g�z�z-%�G�j¢!�X�e�&�7��0�!�0+u9����(��m";���Յ����d��T��������#����Β�:����_��o`'�c��#*�ͫ=v�"x���6�צ�e�c��Ї��S��e�ֳ=���.����>��pv1�o6�63P|���6�Ӊ��ʱ��t��*	�X�dH�>țQQM����(�y#
�I4t�CG�������+���Y/�YC�,#�jB��<����	?�6��M�~E�8t�O��b���\����.=(5�L;3/YVv�+T̵��
"�<n�^C �#�;�<����o�*��2�O�#�7_��e������
,^��f�(�G��f�����s��h��*
��\E�s>����jWgM��ի��)PV�j-�uh�ݾ���.��{�B�M��!�mx��$�o�����Y@P���N띃��/$eܰ4��K�o�*�6�
v-:9ṙ�4ۈ�r�����[�Q�x��G�q�K�Q��T��2l�k���}DS0�Ŧ�h�ݎ;{K)���7�<V#~��{�q�a, ]���&��#�{��i�<!$ ��V� h�D��QRScI�M��%Uk��@�W��� ����6�N�o��!a�Tb��]8�V�� �����/a~F`C��![���}2W���[�������:����Y�ӧ�YHy'��x$�\N�giU�Yb[���^d��]a���'�,�q�]��W�nZ�ͤ�����h��U�5�>.P�(�"��v�y3��+T�BAys 4n�sY5i�S�o�чD[���ǖ�Eɤj�C��Ee���OQhT���Id�g��7�/������"r��(�ಕ�;�$��&��˘Y���fL�oG�L�B���H��ɢ�&�ܷ��5��05RPc�[����sĹ~7�ZgD[���B @�_� �za�����$��e?��Rݕ$��Ѓ2 �%(� uf__=S��Kqq�=\���<�ӾĜ_UV&ޤH���spY� D���L/�X	3/���U����(N�r��)�,/qQ���%(�j���,"8����Zc5=,G!��\��`ޢ=!!!�1FB����"�
�l`��a9�5H�܀��9��k^KX��Z�ar�Ysd��ʇ)���3��tV�{�l:� G˧4-K�|��AktA?�n75MSo��"A��$��?'��Y9M\�2��O��4�8��P����h�kXū9��e� ����%�6�⇢H�Խ���)� ������<�I�j���$�2���+�چ�Qg�N 08�/�'l[�5�O�-
��P�,\ �.���h�C^����3Z2�?������#����Z&P:?�^�d
����3\�,]��c,!S�fa�\��v�|J|3��V��'c���[i������H>����)^�a'[cƵ��3�e��>�-#�OC�u�%;������_6��ť�pR�����ɣs��{��-��c�y+�Z<�98U-}�]��X���\+������9���دOӯ�,��FT�w杗�<��N�	+��fйsSG"v�D���c�_t޲<�ɀ TL[��
�v���_��A�vX�VѓNJ_��>m��u��IK�F��p8�1C�g�ڡw�R~6'xY��O7ZA�:���j0���U��KKJ���_�����l��j�8�o8��n�mE�XL�"~��|�h/'5S�i��}���W�AR�E����'Ӄ{/�{X_U#�[\ݛ^�'���ױ��K�em���E݊f����~e��B��HznGɡ���O*ֵŨ%�Igbp<��P��VG�O~�}��p�Bk�)��Ҕ� ^�V5 ӝ(�?���z%�p���#߼���*�A7ǯSA�L{����|��$�V�Rk�q*�;�V�Լ�)�8��$�>K�����n��M<�*p���5alZ?����j�ӴX�U��w�g^h�[�D��ڋ}�o'@;u�����\��ES|`<�P|�� �-G����익���I�Bm)&��+�rk�d>�6�h�KE��V�y���&_�b5�k�!�Ǉ%��q!�!&UU���Qe�iJ_ƪR��5<6 1C<��o��h�:��R.�4+��b�c�nt5��[�o�,$�������S�h�`qD��5�7�d�j4��R&ok���	�yQF?��0+�e;J&#"R�a��,�V�Td(��38mZ2�O&������]�%�ޒ��+��FR��^�+�n���1z�6_���2y�g��lE��A�Q���K�!^*$�6��n��Z*I��<o]�Fi��W�#��6(��sE�	�]���\V�`GN�h���ӏL����m_*c���Q��ʿG%'�,Ϸ�>9nƨo+���:Ɖ;e�Z���U0[���xgq�
&���^?���Q4s��Q�:�ҚoO�� ��?ɍ��y�|U��$p��F������N�����x-c��o_  �"�2�x��1WƮ\�-�����@-�"�6�[ѯrV(!��ƽ^L�{�UmT��u���	��^��1�0v#F}�<)���v������tą�(AY_*����S1�����h!VSH�`��K���v�8ɠ\[����Hl�[��^~R��1- ����vI�ys��Il+QXp�;������	Pm���)Fxoӕ�fwV������w�\]��ڇ��_D�r��t�j'�#("�	ՠ{�.��b�}m�f{��v|1���w�֖���k�㬷%�r�t���/6��Z�mӉ�����t���5�B5wV�]���ԼbF�-	�<�¹.F?�a] �Cqw�D�j�'� $�E#
Fy�OR�݉5���O�����d��~�b=t�$kꈁ��~�0�X���~&
T��	���)�5L��=qƯ��M+	�.��oܯ=s��y�]�o�KTdԮ+<�\�Wd��/�8Ƨ$�v^���t�bӤ�t�rh�N�_K���r��ha��r�+��ɗ�a���cA�����I�2y�~�0�������d�Y���`Pͬ���j�e�5vV�x)`{=VZ�&]�q@�=�a`�Ж��J�NaM����:l�K�>mh�By����˒�G�� *�E��7��蜛���0joiV��<����9��^A��%B�p�8߽n�\����]w#��u}�+����_�p`���%ʺ�A�׉"�ZU��Ĥd�`C�sU�I'?)P�n��G��0�$����A��:���c��㫬�t�?�&�|m�_I�����:`a��:���_PN�
���9�BeJ.Ρ�d28Eč�.K�\��!���U~��Β��BvWՓiZ�W�ȳ���ĸ��FC4Z�38Qs=����z�����������)фp#���$U^�1��evv���Q��\�!�YV�|-S�-��ͥ�(�6W������;|�\�/N��V@0m g�����ϜH�x{���0�>Ճ���*�b�A,Ad�".ȆHD���� t��)�f�������4�b��ֶm�*�_}�uK_�EK$!`��ޫv�C,�������8��"�+i�1�m"JD`�>b�Cd�Bʪ�}+�� ~/����-/	Qg'r�[���4���j�4�6r}2A��6� �<$c.J�`"��Ф�0q�zT��֛��>d��+��!�K�^��O�e�S�YMM�'��Bq�r=�u�ݰXRQV�h�E:�턾�� r�ױh����\ʵR�!�l5`�Y������g0�Ky*L��`3�!u��Z혲Й�w"svƬF�)���oZ�4
�g�i"�ӵ���y�$����*?J�Q'4�̄��x�	M��7SW��YX��C�p�̍���9��#�V��Z��F5�N9'(��yH}Ҋ�\��Z۩�b6���K��2C�ӋD�C�k-�:�+�O��K[�)t��Ϳc不���N�x�R�PY�v�,��[
�9�"�Ґ������܂"n��Λ
�'�-����ƽ�^�8��z��z'��6=](������ڥa����!Db�KBI�L�G(;������2�5z�j4<��И�P�y�rr�'�`�*J���yh.������H�]�"A?p��Ʃ�j��:$�7��Z�{[�D�~I�LhZZ�;�ʼZn�!R>�8>���,-<Q2�C�z8�q_���%�0*�#b�W7�WdT��Mvs��7��wF��D/�O��@�~�IP���G�r����r*.Ҭe�w����=�_��lT�\����P�Ԓs8�O�A-�c�����+s2���sM����9�TL�Ӆ`�Rb��s�L�ϙ��	�x�HY�ud���H��c�&B�]R����J��J8��D�3a������t���G:
��ev� �e��쬁���`O�n)��Qn��~k�Y��;�oT-Q�sW탴b�-�����b��,C	�Ϸa?�<07�3Mۃv��Ҷ���[�㎅QA
bҬ`s9�l����+��� �����П��$o9Ե���,���mwJL9J3Tn�5�^���Tɟ��B���:B����h�Rs���3}��NT]=��=A8G�fu8|j�V��ˉ,C�	�x����TB�d=�@�������H�O�k�s\��h�1X^1�LQ�"�u�� ��'����;4��3���J��K�2�U�9e���t��|v��w���"�M�h���fh�R� ?D�Q̕GJ�=�%qh�|8��}���E���^�����Jxu���?�����d<r�Ц��k����.�Sp6/V��̪�v58�reQ��W.Wh�A�T�߱-}l��U�G^��J94�9� Pz ��7ì��w@lk��E��|�N�������*T�7C��
����Oa� 	����E�ua�E��zY�b7x�߾8�a����&װ@��1�=�Hk�����o�ϩ����u:��9U�7��o��b�p�>Wq��+!:xi�T!�ʆq �Qwk�+}]24&� r:wn��rj3#�O[{���BU�w�� ��˵�8�/P����且q�ۉi5�(0�C��t|G��(F�/�tUy0�\�f��$/��3�9<�ѦG�-Z9����Kj]���nq�b�������Ri�Q�$�ĻK�RH���}˅\��Oƨ\�#�)���g/�XF�>����zE�����R�tg(�H����"pfƻ��7KJ�KK�p,fe���U��Չw58��!"��P@.�{�H�#�NO�H�DI�j��F�k��'�Y�ĹZ)�NoqVu�u\r����b����-��]w=��N+L���rGP��wU��1�9����AI��=�aB7p����)u	�
���]8�@*��6�W|Q�Bn^�����A�	J�G~�I8���/�4�=J|%iEÐʺE� ;��-Q]��UV�b�H��+~&���l+��])\�C_7�2�VD��[|��q�tP~%��`���hn�F~�̓�z�n���I��1�	�#wЖj�gY3��Ȃ�42j.�̣l���:z�IOmc1胂��o��Ԟ��𱯬E�"T@��>6VLmp���t�UE�HM_�ko
�\����\�7�2�h��P����g"K&�P)�T��k��*���2���jl'$bJLCus�w�6���uS�$�x�(سYh�Zg]��ܐ��}��-���Z��|R_���i���dٷ
ԭ��h(��Mwr ��q�X��c4^ ]U�R
�Z���La��>��-�PA9�̕'����J}nG蝷���%G�������ܘW�^(�â+����:�d!����2I���L֙�#|\�G��YyU~?82��YSIP�%�;�{���k����_$*��V�{�X2�*|@��R]<�'1�����ݕ�cs�5�s�LF�)K8��LZ���4�IJ�f!_z�ƣ��ri�`�<(-i.x"j4{Ś n���PwO��=�"�����	�4�y���ܥd]҂5�$�}Rc�I��[t��f
�gg3�O1'����?>/��, �9z�:*�� Q��Ȉ�O� I��[�N$mJȝ�k��N��V�r�ٝH"�&$Z{w�E���I�,�=_<�`[Pa��]UZ�v�g}:T�\�xDV،s}��|�:/�we�x�^ga�a?�[q	�����FB	�#IXv�M5]b�~|<#5mxx(����!T��������M}������G1�l��(xG������.c�s�������%�A+��3���Ɣ��@������f�"��&��ց��k�D5���Y�Ĕ5ՍH�]�U3�k��&�;+6=�o�w��H ���{P��d&~4p#h�|��I<��X��ht�'�5��T����[�q��Ϻ�����N_tD��i�[K�*;p�:�*(����=U.�p
��h�I�w�Dba�j�+?Y(�^1��}��mS���1�@���j�RU{HǓLe���L��E�r]��ā�
?Im���$􄥭������l�G=`1��0�#<���)A�̰�pqW�>@�Xd�+��?P�J�z(���s�&���Q0��>p�n���r�)���p���&\g4� ���R-U��\
+�Zg�n�.IZ��9����p�<��B�%�
��ZX�jGO0��ʭ�? �� m�����y��1���χ�'�W�h�C�����n4������7��;I�@��cC�$n-���Y�O��uyp�K��
�3KJD��|���ĪA�T95��Iw�>�$v��������6����JV��*w�PЎ �T�'���
=����)лԓ�]��Y�%�E�6�y�,�ͯz4�pӋrƺS��#
���0�b&�樾^����S_�����Ew�A�췝�ioP�j�=� �,�y:��Y��
bc�A�w��6�;�P��ɣH.Au��7Zp	�ݒ3�$����2<b�uo�B�(�,�u���|�����v(��*�L\�𑸿J:=(��T�oʥ�l�J�.����ȧ�?Q)�����E�0,)LM9T??�ޕ��c��0�j���D-�NE�2���g������� r��Sr��!M"�Oi/��𐯌�^@�0^�C���h�8''����O���$�����-��}kRzا�����rY9�K���ˆE��g�c��<�b��9��RЙf�W�����NOJ��=�ܣV�i^=l^5�P�X�~y*�c�sa��9
Շzژ�h5��
�H����c���Ъ����Q����a���Η{�8&upj�������_���	ٖ6Y��y�Qh�ȫ	ZY2��|�R�Jv����y	�Ͳ�U�ؾ,�1��WX���HP�{�;O�;�gY��v���-��4&kT�����0�6�4����WH�i�QKi�T��5��k�m�젣�1X)ɠ��b ��Y�2���SR?gK,������w�(��A��}Ұ+xau�fJb�ͮ�*�7>-z�Qbg<�V����=�dvFb4EZ��>�C��">�G<�+���z��)-�`EdT�:{�.kx^�^x[$*�;�(�9�?w���!#��-���499N�l|�DS�G��n�C�ԡ�{׆\l�B}���U	�i�DU9�G���K1V���Qm䑋ʫ^��	'R��1�c�V��E���s��43S�m����5h�Fmag �-�M�_�֛O(�%��z9��a' CZ�L�f��ʑ,����Q��ܥF����QR�V&�d�!	���4-��q���N�R�eh��B�=(9�OG3Ҕv�d/h�S
�"ï�kJ����L����M�\�F��|�E��K :��<��%A������^& ��a
��)F-H�=Cd
%gwl�
H�,���{Z� �%��N�O�!��O&���J���[�,����_�jW9V�'�5��V{���������0yqA��z������̓DL��+���A��7�s�U�y��,u���N�_�_�>�k��v>�G��'���A��f��5�W0�r�����#���r�Y$pIs���s�ڄcƚ�LN<��{-����$!aB�.���*���K	@�;�ϕ��y��ar��>$�>�݀|����cLHm�{6����-WysFy0��٫�_�n��eF.��>
YÖp��J��<P�,#`��PL�~w�2KY�~c�=��Y�&�GK[�utli*��u|U��0�e{-�s�{��v���A�����L�C>�- JH�)���3@I��9��MsX�%mǄ�
Wc�#bF䕝�qxEv�����-!2�Tr�&q�:(�a���Rm(!����[�����>���|�Hg}(�^�Q�t+�5�R��Sr�!��*�}�H"K��Wt�3͕e_U���_��'5��%�:������՞���HO���a�l�ؤ�b[�	��?�;9��_���Pʖ���D���G}w�E�a|��Ox�VLX��)b
��jj�w2FĞK������^�6�=�-x���n��wf�?�>m�UK:��a�,��=�}��D*X�J�ur�jW�5���Y�(.$�����ڎq�T�.� ���7�"���*����\�d���y�.�v#��&����Aa�5|d�@�(K�h~�.�{���m�E��$fE�_x�ϐ�K�7�]���{!���=�[��q�8�ȇ�����>=�}%��K����Jd����	�
2*y�>J���j�)aӽ�3ۭ}������`kS���K�{�5�T�-S��T�M]�e/9v���l���b�}�t	/�&�(�)[e�^�pvp�?��'�cy�*�����f�u'��0�YO�����B�a9���2#�oAU�{��ɩ�uZ>��$�em�J���^��z4|[�����Օ�C�M�i�fpX��:h��苍q-6�����U�U��N���9H�X<�73eŸ ���`���Zl��4����rO<E����w{�� �u8�޾x�Y#mk�֧�X�1S܌���5#�I��P��ȸ{d�_�ؼ�� �o�nzM	>�ߌ�,���%�|�&M�#Ƕ���:�|����ꠔ��y�1�U.?O��o[�3�ү漁$ӻ�*��kR�"���a
�f9![���媸��';�֠���� �k^��' 4h��ߥ�I{ȁw����_���m<'_@�]�}�N�����	p`1���C	ţ�)J�K��#�0��X���ʷ.�����Z3����]�d�H|B"�NJ�X׺f��-�߼�f6"{�ss����E�A��𠧘�g�BP�D=>
Z�{�`�0v#&�ߙ��z���Qiq��B�/�=c�Z�Y��gQz�'T\wfJ��^����`�,VZ:
��b�ʛ���-�L�V��0{
t��oR*f?�Sjţ#�tPG��êG������tydMBu���l��*&��-3(<┎,q��M���T�`Ӛ�|�*fu����/��v!�