��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�!��
��%Y l�׾����|R�bD�E���y"�0~E�@���FW�{�;��d���m���/��G�k>�t��_�����#v$e�[UЛ�բq�aT�m?K4�#��.,�0A��(+�+���+/L7�J%�`$�{� ���w��tĶ@%��:�b� X8�cZ�ҶuK�c%����=��(�LO������(��90�_�5J����zð`U=�2���ǋ *���[R59}.��o�K1����%���|ş�&=���~��Ye�`�f��mF�;4!�_�f&�\ݗ�Ir�2.�n�\J���:�H� ��t�n��Z3
�A�Y���gب[��c���X�Τ�#��
Jv�N0�9�+�#S��. �V��1Gv?�1�跜#��]����o��$Q��7�+	E+}�,�j��+��Y�Sas+�~;��?��_9Q�l�T��Lٚ��k�w��=Z������{� *��(�]O�;�ȣ�C�-6n! ���X�qC�B���7�|�2�1F�ߚ�]�U�HqpbK`�����k�������K U�܇��vw�J
�q��+Ȓ@+��,ƕ�H��x-��R�sH,���(SD�5rⵚ80�N�B9�at�F0b1�,�<-���{��$J;��; �?v_�5�&m�Wf��h�S唺,�������`p�"_�d"$����LA2��{��<m��<�1@8I,|,g�qo<Az�9u�ح"G��Z_?	3��[��ǲ����v3,!��np�l�)��)�~	�l��_�@w��L^�w3p����&�f�<�꣧v�L܃�xx�n��8����&^���?X�C��.oK�R�V|K��V�A��HM���j[��(C��xBG��!D�Ԫ(5�xm2�D8>�d>kT��sz�\�#�RH^��� ����12 ��|�2YK#Y���ݢz@Z�^d�S8�Ͽ����n��2a\{����^$B^'h�u��Wv�v�{i݀�-�Q�/�t����!��>���g��]C�&�#��B����0�F���$e��6x�?�$��cvD��_lK�З2g��]���B�����EvF7�Ua��C�/��S�P�5��F+=��WW�_�7���f�Ɛ�4���N��u�ނ��h����CW,�9�"���)�@�ww��Tr�\��'��e�Nj��ْ�'Е[���}�H�mHAt����Jrl�7~�3&��S����w�����FL!� &[�-¯=P���K躃r\��SL���$L'�NK��@��[�Q�P<��@ ?#�m��
J\+��u*c��H��Q�Q�#"�֠>�G���Y[� �=8��v�#�ٻ�!'�|~�`qٸ�Vˬ����9q�H5���u�B(�3��f����%a��3*\�5����:U8pfN̯��g�ΐj4�RO��&��H$�
��K�U���ISkLj)�������LE.5�0j���EH�5�����E��h�Ǧ�X�(����	��M6�l�s�.�+�O�O�>w��B/7��L�1.���AF(D�[�s;H�C���{�8m�O���Y�>����Y�+������|u�n6mLK(BE�ًK{��#q�����z� �|����aWY<[�y�ji�q��'����O�"��Lv>��.u�/��vH1c�]�#��2����\���kč[0Fˍ^���ݞ��j���_h!Kڜ�T��P,���#�7��e�#���FvX�ߕ��{�r���03�����`ź��!x�#�{�i%����<`��X���/dލ�2+dХ�����r��Ml�Z+����K6Ӕ���宷 5*A!�x0uAS�|���I��fO5�0�!�X�񺑑�''-�1=��ϻ�7�r��2��}�fh����i�CY�<�����Y	H݃5��l�m��������4 <�	(���1��ɰ��l�҃�@�
��`��`���8��>����ߏ����x�8i�w.Ύ�>�R-Ȑ�Z��a�qk|�q���.��i���<���I=��ާT���Y �B�%9�ANr�!k`1:<�~+�)g7��A�����08�f��h;�C�w�F��E/�V�Ah�N�Ѕ����!VN}�ƈ,L��(����0�uOd�X�k=��H~��\�$�%H�%�yi60�A]t��,�T�"$��GyK�-��Bj}-�n�]S��sO� ,��B��Ư����v���[�ڃ�bR�� �4��Oՠ.��TĀ����~�^�Y�Ne�ԗ�UA��a�#&^�)h�����r���k0vI�ݢQ0���?���u���٫��'���[{�R*k	`5��@�������NǬ��ʳGf�ާ�QpiIS��3�{�j~�z&~|i�τ�W�	��T�)1uE�j�~�Q�8{���ʦ �d̳����$�w�ֹ�>GDmæ|�R+
��p�V^4�X���4f��c�n.�
|�Ģ�rh�k��|bOS����fYkA��8�-;h���?��繸����ͽG�U�㏳�g�Jn+ͷU� �|2���&�����W�G�Q$��:�aC�h�~�h��_��Y;S^2g������;ݴj�����j�6f�d$j�����؉^�D[.2P����B��wƁ���3�n��Rт�~���f�yFAz�<�����i^�[$t����J��Ybh+�9�t�Lߜ�0S^�\��qK�6L0)��L�y�1��X�Ůô���uEp��ic���ȉ4�0��u�3�%>�HH������\��Z�u=��{н)�t����x��|�n\�kvO�
�$ۓ]�@0Ҡ�jU�J�c�?�7�{@�Ⱥ92%�𱛖:��-�Be��?�ť�Y�<�c^D��l�s}�J��+����Ǽ]�J��	M9�fg����rG;���,�ڒ֖��|\P�����5׼�T*YtK[M�!1+봈��p�K���#w� �i�`�^���N(��3��Ϛ���}�+�7{>tp��C��
LJBxf��pxO��1�3�+b�1q�}��[3=�o�$ j�D��K"1�O�X5M��V�� �w~��sү'���=L�hs^h�`޲W��gJdM�� {΂�ťO�����V=rj��f�%�<�7�<)����D��(�}��h����;���UQE�h ��i"�p����M��	a��\���.j�v����	���e�Ĕ-�4�`��E�Z��&��؀��x�!�u%/����~.7���ߝF`�܈:y;5�)s���C����a��a��~���I�"��̓�@����D|I��-� �,T�-M��c��Yu�5�E/.�����<��V��AQ5$ȑT6Q�*��#m܈�pT���e�Q3Rt���H�ے�Em�y�+�(Qb����rk��M�>Gj)�IP�ij�������(��i;�M� ���	wJ��-�f���ǲ�C4��R��`�Y��6�}��.'۰k#u�.sQ��O����j�>���'�����HKF��O�L�·���r� HJ�y
��Y��QϦ.^�Q���f����/�Ν��M!�ޏ��ɀ�t��U��~<��5~;��$cɳDR���+"�1�f{j3��
�D߸�:�-no�3�
 _�����˝�m1�0��囩��'����A���>���x&BWC�d*�炔?���2K�d�X7d������U��TS���A�T z+�۞�	@-iM>=���ǻ0SqH>�@{�����9>h�[��?Z#w��"S{��nڈI����
	�TN�O�)/�2�����8�Js�N��o�H�_Oh E	Ae������W浮�AT��f%>�wb��&�[G@�0�W�ڿm�|/�#@3v�����Y�q��dW�v��J��@4�����~P|�T�,Փu��!ƣ��.*]�Y�z�en0�	n��D���ယ���J�{`�4�S���=��h	D�$�Y���D*�)=�E��Y����6ך]w`bҶ��9���Ym|j���=��	�������i��j�}}Y@�cD�jvqWx�E T�A��>�N�K�E~�̬^�*���x��vm�6�E�Ǐ"8Z�b�;/�y[F^X�L��~����^��y��.G���_��s�N�;��f�sI�5>�c�٫�	��~����u֍�X�����S6>�Vf��7����E ,��FM�A�`'�l/Q(�#9�B�'9�qGUz�yRjFp�X�1�&��C:�s���0�gȗ�s2��R�|{��P4#J�y-�tP�i|�J.C�i��>���H��Q�;�qc���Җ�����jk8�W����B���+���Gb�:�amƁ9r�sa��?,*9���Hzf�E0G" o�T���(cӵ�U��z���56yl�c�0�����)�T���T'|��p���/�^nm^�f!CX��~z�#�P�[��cH�Hn�׬�sK}�'��\%6�jB����X�b��[��SȖ�b��7���ʀ�>P�B��a������=d,�m��q���R�b7a��#������
� 5]�:��A�L����s��U5���;)1�_FL2�-�B��cᇑ0k���e�N���})�p�i�B��R���J� ����Ҽ7���0B��tt��H��{����? 0n<`2c;�1)��oG�6�6��X������Q@Ü�"�,�����}1�G�~t@���O"�ɧ��'�����e�?��ŏ�����(�Α[�P#b�K	l�^~9���pB �0��d�R���MZi�+c.�n4�]�F,Yh_��\�~R���h^b�P��������x�� w�ױ�5WlO>�#os\]՜!�u�%=�����֧��༩JJ��ޗ�Y��2��n��~^���X��[��/�.d6k�X�8�ͯ�5�!x഍ty������6	֊�Erz��֍�o����BI��g��`@��Ǵ�;t d[bJ5 �f��Hw�\7������Y高�_)�p��DV<�D�t���z����_�4�lv����+�a$����υ~�#�o����G��5�g��>�����$�]t�,�UK��N�)),�<�'Tm�ypX�3���x�Z���e�ywbL��-ʋ���ʃ�n���A�#�^�!)��l!\�h�������{~m���/~����Ԕ��\`9hZEB8�n�0� Ʃ:&K�������v�h�S~���k7h)�F7�.�x�����S	f~����ٹ��ە��� }���"�C�SH�H�X��*�R�
�l��3ڿ���g&�'�)Q<�h>n�N
i�/�g=� ���A�1k�nU�w;)r��G�\��F:�w�:����v]!:��^��L�cj�5�vP���}e�&� ��#��Ąg=�4�]M�O����;[�U��ZFp(����%])�g��Or���� 0N�ʻ�Sn�,��zج?@(�W����.�_#ҋ�I���57
�)�g��m��v�&<����չ/�e"Q����+�EG�4��-��|�ɛ6�����'F�i}�%x%x��p���/te��CGzm��1R��_ƟybO��Y&}J�ړ�(�0�� ��ڱ`��#}��;@|�vM~?;#�F�F �\��3�'*,'�o߷pO����!���\X�Q��2��� (R���p]����Z:�i�4���_���h�OQ��%��Ơ�yK���🁃�?��bq|���E�草��rE��*�A���b��:\ZZv���
�b n���@LEw���������@��L`��F�����%���Ċ7����;�����
T���*��'Y��*\:�u��3�p�;��Ź:���x���ϧ�m+�{O4�f�K�!��a~�x&K�[����X-�����5��Pl��(w�Ռ��E&��t�?T*�FR�������g��~�[룔d�ێ�£/�t(�}>�V'n�p�*�&�(�Q6��-�:Dϫbٲ�Օ�+7u����X�w���e8;v˫G^	|��r=Wv8�H{�9_�y�>2@��#��:]��\����O�X'�=U�H�D8���S���q�oi���
��R�4�D\<�����2y�g-��.���(��5��hu�~�t!zF�ځ������"��o� ����f���\�2�G���6\�ܨLd����ȖC�����n<��D]�G�����������w^�xX ���4����z�2l��CE���~K�NKB��Ӳ��3,���ћ5����/�ޮjFs{�����/& lF�p֔į����G���]��ӛ������$Sߕ���
oc�?�8N:f��v���E1D��;�8k)S�e�U#��d��t8.we�_D�N�ײ�ͬ�X൅Vҡ!$���#x����u�#�S�,��d�sBؖ�,5�� 6 ]Rn_�71�+���<��ޢ� 5���ɜSHH�;0m(���h�I���␞֌N?�7@��g3��ҫk�V%���?��J]Ȉ�A��[aa����5�+<�w���:��`��6:�3~��4vS�Ѣ���f��<9�Q'�]��s-8l��գ�S-����ը�Ш9:�f`攝�
���ȕ����b����|�8��RW:K��M[H����D&o�6�eH��uni��(�ə=�'^χZ�s+�<�ڿJ�"	�.�y�_?ԉ����b�ŉ��C��@���)~d��+>�Q�ۆB���1�.�P���Uޖ����Wp�I���)tq!�b��f���'������z&d�:�e%@/'�������s��b ��y�ͭ�+JY5#�C��L��?� 
c�����O��լ̋R�8����k�"�a]BX�o<��L'��NĀ��V?&�z��/���?���Ŷ˺�#fV����.Q�2�~JSg�m�c��F��N�gt	m�NTJ
9����3����$T�+˨[�\5J�Y0�Z}P�M.� |(���̸ɮ �(Y��hޅ�z#-迫b0tU2	e�_\��[�|���Q��N���# �,C�WvS��X	�Uj/
ec��!��	I3��o���sZ�֪ ����f����K'�wlc��t~�qa�?i3̀�vwt�?Q'D�lN�Ɣ���	C�a�;���W�b�)V�?��&^M�V@�iÒ�n+�1���q"s�}�'zg���L�q�H�)z6'�@�D��C�x�	���xl`#a*�l�ti&�
���sG�I�~,xė6��KG�^��U�P�{�;�![��S)��)99�%���󧲳�i[�T���C�(,��������(�j;�b�w�CN���W{'�uۊ1��V�C�������XЮ�_��L�e��G���(.���{J��sIL!c��T4'/��,��7�gK�9bY����l�5ʾ���C|��Ԥ���*�є���p���[L:hJ>�[0:�2v�J��V,��@�oDh�#&�N�1\hStx掔�\��`��y��9*�1c�qTP���ŎD~��D<��%N{�7a;����y/��;�x���B���f�v��q��b{c�'���4WΌ��(�WVm��S�+�P?���aϽ[����6*[�;�p���c�,��P0�*�ǣ}�e8��s�0+�����(Uq{���E�I@o>-��dMğ�FP{?���z�Йkl������piV4����S�kd�Ѹh���@zΦ�e�c��9��]�m��l@v��r���)�E�Ug�����Ȋ�*h�N9Ӵ��j��h���_+�>���*�%��;�M�2�����F�vw�&�m���}�/L��n~����ل�)���Y&��>�أe)���R�E�}����ۦC�ܞk��\&�qB BI��R��pj�+�c�g*m�ۃ���[�<�#i�3��5,<�iJ�D�1,��a"&'��Z e��D��=1���A7;�2)խʢ;����;0��k���Ύ�E���\Y�<�k|"/������!i��{����mk�V�Pj�aLC�t#���_�(�Ze�W�̟Y�_1X�6a<�b�#�}&	����lC/v�Ur�'���Q�Z�ٖ)U~�\j3k�u�Ĉپ���3:pﵳV^���J|��(	�o"X��b�%+!�W�4ʭy��}����C�o��\P�gD�"M�s��7��-��,Q�o�����*𿱷%P�U�)G�d��7q�vW$�a+��S����QH>*~G%�%�;�M��x�j��9�7����9t|M<�#�<�|,�̽4�H�U�y,���@4vC�U;�	(�R3���'�r����A9Mp@$e�Ln� -��Ć�X�<�5�E��vp�'Q�q����<���ڇ%��q��mT����7Y%響hu��G'�bd�.Wz�����[+XXm��#���
i��yaL�} ,:_�����qK��[�c�M��i����������h��`���$��W����Fؒ��%N����`H���|C@�^��[�q�fWH�D��	i��3ɂ�-��>���^엃_��R�
��<����Ĕu<��9�暺_�KS���	Ař��6�sa���z=*�"�f�vd���iq)���u�������N����_W��g�UyW|X�������������d�5��D�WW�mɪ>,4��l�o*� f0��Ԉ�W>&";p�P���3Z�6c�c����a��f!>�؆�����e5Z�!Y����' + F���`+\|�|eW�fU�T�웤m�I�.���~P�e[y��#ȂyW"�gC䶃h�iox[sI�[8�������YY��ɒf�F6��.n�4�P���-a�$�斤1M-��i��H��.~�ћe p`uܟ;�K�A��'P�g���E�nh]O�G��\��MsL'zcj�����Qe��K%!�d�����"����0�Ms��]nőfꤊ�_��_���0�^l�\��޼"�ح�v�7��ݼ�l4�՟}~��k�4��
�a���"B��I��yPM�	J��Y�4�ɐE3�ƺ���l�}�<��8�K�9r�9_0��8�/�9 o�����`�5������%�`��j����G&A�i#ScTU�3�^�yT�BuJ�Ź��B&)Q�o�s�ը{dM�+��Iug��].��ο~n����$21Wj'z�B8�� z��f�U �E@���W�^�+i�/��	=�t2�C��H?SC� vS�0O����0:9����D䴰��6�~�J���s��߭��
\Gz4 a�g�a�(�ǔ�{�c<1ڲ<�j�O��y?��8��X7E�Ȑ�NNѭ�	f/�EH����s�����H���u,Õ�$��+M�x���4�t���?�멪����3���'p=�*�s.�uN���8c[%"��U��gMf9��`�Up4ۑG��j�L��&���x��G�#�`� �O�rG=�bC�!�\B1*l��fp�$���Z���<���"#(3Y�ޤ{�I���j�4�v�x�}d
i UK���F�|�MFG�
��W�(��떈a��h�_܂�a�	�''#R0Fc ��?��j7*͋�w��C'E���߳(�@nw
bMP�,�_��j�)����!�wE�k�z`��&�x�e�`_�@��sYC*n�#	o�*.��΁�Ѵp���q���U�,�r�J��/���yغ�?MKX��RE,���|{�~f���q�w�t[g5"@�&CE��	@�e�0|hE,Ֆ1���G�^��I����t�� �U�s�t��9e�zv?�fL&or�����0���_E,*��8� Cnq�-�ϗd���d�E�`'`�7���"n����A��\�����Z�/R�=j�J��@�ܜ�B�=��ڊO����=��/X'�J��%����)3v����J����}PH�Q4]�u3^ Ig�yyw�����'+��r�(���rb�a>?����>����`�&j}ǖN��~�Y��xۂ���ȑ���"�P2�(]��x���T��D�ñΈR��Ve���1���a�g����z$�3�'[x$��Cǟ)|�ڍ�nbq�r}\�<�
)c"����x��8_��ǁ�ڜ�e�9|����D@�c���TW�����$Q�6����x�۫�>[_.���\;D�W؍Z!v8����ذ�]�hُ�3��?3x��S�[u���%�	��SAA(pJa�įˑ_iNx��WS4䪩�5c�{�>s�MiB��I4_'�z
�	�t���'�Yo����V�2�u�|9_�Y!6���ꓻ��a���7G��UW�:���[�_����Cb:tqt��c��0�Y�]Z�Lfu�����ԫ�hIX�\$#f��~�J6ki�Z�B�̵k��rk��Yآ{��^�48��n�j8:��u�)Ѱ%�@�(w9 �&A��?�}��L��H�D�נ*J�]FOFyu��fui�1k�l#�'�~˝�t�<���	�����2��U���Ϫ^�+����^��<�Od�
*#�c�@Qn<��4ڹ���H��^��.?1�ϟ�  �f��6_5F�a�K٣ &<1yc��M���[/�n�.����W޿Q�p1X֞��o�6h���~�O���b#�|FwK@6	q�2��o��9*���4e��~�`ĆI�d�/+�A.�j���G�)����R�	[x�"[W�|���:m�i^]��w)�m�d��L��5^����Aɫ��5�'����m�?"�-��>��xt��)��6O0�/�`ƃc�'���3�C��tC9 *]i�dk�̤+��$�����*�hF��m����㼔�i[�w�Uj^	t�@�C�(~x�|�?`�f�Ą��Ы����;��Y�-h�M�*c(�=�Q���K�z�Ip������ZVZ�2�"��y�_�}���[�p貓cO�3Q&u��^7<����-żJ�:l�CÌN�z)��d�k���g6�"f1�p��vC�HK,��
�ܨ|����j�c5����Ok.�4Q�B+��J��S N�����T�e��Wc߾��* ݿ:�/���٬J����>tT�M�����3U��Pk'��?hqT�j�$åGL��K�I^��J���^���,8���TMx���;M��y�3�l����
�$W�Nv/���U%I{j�6�&êӋ�G�)qZ�w��F[L���@����U-|�'}RNhh��w8�R6�:'*��c�f��f��v0�c����Ú�E/�v��4��	<�-�Ū�������yf��:�������D@�.>e��F�ۀLv`|&�w��'{d��;�A0��*�ǯW��&9�21�������7�VI=���'/&�ߥX7����;?UZ��h�~50s�ݏ S*�#�dP�$E��\�:4��'* I�-n�H�5/:a�8�?�o��dT���\��$B����z2?z�2MEY+��z�TP�zG�n��C�W�E�J7H���,n o48���N��tY���y!�� ��e��̮q�fʭ1E4�%"#��w�i�̘o��uڰ�|mt���.�_T7��������{�!�B�-��:_h��k��ȯ��+�Ȝ�i�c9�ǀ1I�v�(D;ج�l�9�춱5n�M���}i�/�AS��>^�9`H��l/�&j�E�m��\�)%ޮ���w"
Z2C��ڕ�}��}���{�"KT���&�,#�Tކ��5eG�ّgvnW�?#�*��˒a=(��yԂA0*ц�8�,���M�������3k�&�89 �O�ѩ�Mc4�R���k��(Z�aXG�5{��Jm1��3t�}�S�뜿<��
<4�'���|k��6PPJ��V�J���(76#מS3�L�e����-%��3���l��$�k�Y+�r���2��ò��4}��y2�Hҟ�w�A���"s}-�Wk3Pc.���8�(�_��;���U��	�ӏ�f�AE�y�	�k3�w���z��5c
�)�Rr{ZC˛J�:L@lOyv�ם���aZdP�o�x8�Ӹ���.��!� /�yl��8�k�9"S��jb�7mkM=�G��3�2MCnO۫~.J��)ׂf��B<erd�9�
D���<��� �T�9������O�CY[5bwKg�n-\8.Ղ�Ckː^�6̈́L���B 8�ٖe	ö_/�]�G��Ί�X	Ki����m�G����>V��9o�3���#��7�T���I��'��? �����9�"�����	���Yq�t8 !�]���gs�Ji�aY�K;U���Қ�6H^C�M"���C`�aE�R���DI�%L�0��-�.AZ��������H	��Er��G�����;����aD�L"���[� B������^8�B�8^��P/�f`B�1D2usZ�Q�3]M
#>^��z��~лd(_��7�-7JQx���͞��CL���&K�y(�uOQ!�4@jG���)	��oWx�L�����6��ڷ��-CA��1����R�eWC0[��yD}�L��5�70Ar5��h��a>�Aa���\���0NnN�#�a}����̳�$3Y-�����i]
��\�{_M䭸b�������ǣ����f���q�Ux˥�]��� _Le�a�[�:#��,��B���|׽)�~�[ߟ�����QX���,.x�w>e�k5��[�Za�vR�f��B��Ē����Y�� �x���H�Pp
#o��w�}�J��h�B*��a���*�i���@ծ�eQ�^_�wnW�D­'��1�'�`�vx��=���|Ep���2���^�Y�/q��Ȣ���u?G#d�Yd5�ǜ(�׏�5���4���Q�N�q`ڱL,��f'�O�?N�=���Se���C�[v�~�t����AO�f�Z���sG�),��bG7���X��^�`����L�VM"\xN��g��d�2�ql��	��/�1w6�����;p$�P,��H�%*O@z�R�$��L��bC-Y�.�R�6���v{D����T�����r����"�\v��M+���z��N���N�"���]�¡����(���<������X��f�eGH"�zp�ܯ�~xL���n���/��2��	#V��ԫ�Z#,e�>p����ټ\)Y������Y�|�j�FG:߶������ÿBX��1Oʤ���\��| o���d�86��e��>n+kߵ�w�ԃ�i3m�j]��>)�Q��{��fQ�sS#��Z>�<����
�;8��wXr��n��}�H�X0y�p�vt���D"v���6iT}���ҡ�O�A�暨�i-Gab_S�?�^�vN�i�ۭa�M�f�P����nIE�'t~���-r9��FS�D̗�B4���ڙ��@3��tJ^�ݦ�*�n3-9Ă�����˚�a��74l��Ը�� ��Z�c�'��Ӈ��2�E�$��*�c�U�006���&ֵ��` 펼�1���b��7@���P�"�\�'~P�Μ�bg%���UV�+��G���%���Sj�u������?D�����W��!`���Al����!�h@VպZ����/S�� P^:�e�x�`��*���P���9�����lp��1֟7�y�B�
����W�2Q05�s#��\�i��"T�NR��B�`�3�R{j�����h�$t%�|�QM�@ҕig��`�/[|fY!��|�%�cۉ]b�3#$&w_*S���^c
���4<���ީr���ӌjiD�����tMB�+Gw'�x)i���wc�61�fn3H������қ-Xܔ?�꘠�B��NUy���Dئ�mlX��d����~�5�J��7LȾ����x$%4�C���׎}�Wy��6�4��l��u�r����ɰi��n ����ʌ
g_�x�.����;Rord�B ��}��~A=������A:�:����!�F�<p��9�:��u�A����:�GE���ɵrٿ�(�نY��IyO���b��ہz�iK̉�=;��w0�Ʊ����U}����)�Ho��)T<[����:T���ػl��H����i���뇖O�ب�ez���p��`��{1��T����u�gC�'��&+���B���?IB���˟���=LL��q�Q��m��ֿ;D���H��&�v	Q�P��z�ɨI:[�!�#��2i��!��r�/��@�ͬ/cy�H1sh��f<s���F����|&���p#WgH�4��nw$�gi���+�o	3LFf��m��c���څP���)5@k�����EK�-�D�A,�\\�j����P����W׷2�Şr&"��Պ�!�Q���uuM�ߎ�yV5Y�'S��#�<���M&}��B�a��>���l�k�"#UsBz^�m��V�G��`4O�!��/?x�
��S[�����u1��o��.f�Re�A��/���J�Ǹ:L2�W��Ă�O-i�[�C��,ī]��+Py�z�^�֌2^�΋�{b�3OC��jv�}ݕ+3"I8i�8[�.+��*�y
k�e�d�F](_��)lw+�p=Rxs� ��׮�w	*�M۞�z��q8�nA~�9n��=(�\���U��~��]cy���,��٤��)�22��Oֲ�(�z�8��r���}Ac��u����ic1�������Z��6��ާ��5�v�Y�1�54��ӛ���(;&q_�ErQ؇6O��19Ԗ��W�C�t,aRi�$~G��2&�~3i���[� q��_G{��Z0�B?���� ��5�r�d6g޸����'�|��pV�0�cn�5�C��	<�)�C/;t���ⲻR�Ь>s�(��юp:����j+�T�����q<�,\kԹF;�kNa
�/�?�l���8�����2]�r8Q��6�cO�H��Kb(���䣅˷��$Lc��"� �T��2�.hO��PF�������Ґnp"�t?�[NdޜQ���B
�Q���Q�*�i(���u<ʗ��tb���Q�HE�*����\�����L2S�)|�%I��&l��� ��`X��bC���8-�zY��Ҝ�2j����
��e͂b��'��-���x!�U�FG.<C�������!��Z�0p�y�I������~�Q����../��5��}8��Zz�^�:X���8��5�aSJ�(=��8�ic]��r���8r��A�R
������/���� �U�����kX�v��I��)�\��ѐƄ/�r���mz�K>��g[}".���a��y���Pa��4�3������Ty>K�~�(nB�
r�,6t�(�'/�v��/�c����}r�&-���ܼک���n�P�%�;{��P�	e�^B�zh
k��Y�?)/��CS��S�PB�8��(9�[�l}{1�rŚ����xHm�vR��F����}:�4����x���`7�����l�0�[���;^�a��H�9����Hx� &U,��BX�1֢Q�D�vͶ�p~����.�傇q����z����Qs��r��KP�DW��r�/Być��&eM8&�҇Bg�:}�v֏���?[!=��4�d0%k��:�H����B
,_�bTl�e��S�gQҨ�7�iw���*��eq��U�-�C��*�R�N�Ľ�mC]��B�v[����fo�\��,ޞ0�)/������A5�Ĭ,���C�P�W���oaa֯,\Èg�+-����6��)��'�OTZ�[���Y#�K׮{Z�M\sG�k)"����kt}~?{��ުs��\�ۊ�BP����ٮ�d!�0��aɎߍpn�hl
L�{����������< )�����u7@�Z�+9�pu|�b�(B#yG�u n4h�S��l���]L���u�L��z!�����'�iߔ�]w.<�"e��z:�#Ҏ��iW�⨴TD���ju|\u=�>��r�q'�����T(bӪ����	�b���,j5R7���x4��V^�{�)�B6(z�H�� F���J�徟-ݸg�:'l��Rp�@�O��s�M�ʽ�@���y���O�K�g	��L��0�b7n3��Qn����*�H�N�)��h���_y�n��S��W��qx6w�2g�DZ^m�j[��ؽ�VɊ4�J�vs���.%��+�������~������M�}��>5�_��\߈��.�{|�$�ע���ՁW(���o2�e'Ŧ8�/��2��)��:vCg?���gy��W���D�Օ^����K�1�ה;~��M�`;Q�G�(wt���A)Z��N!]C�[�`�rK!-��B`И������>8m�6�����ʎ�+=8��;��L��,�d�C�Y}�s�p)L�{��@s `�� ��&�lw���S񤔧G��ԭ��n����}0�1�֪�F�N����"	���J�K]��lO}zQ��A�����H%�]K�F��r�S#{�Er�,^��iO�Z[_J�A%uT'i�S@3�%�
�5g��\�/y�#h},{��j�2߹VZ���e�h2�A��8���� �>q�CK��W0��_!�yW��<����J=�����ꅷZ˄j��Z��JbS�h�Z̫L*s	r2�񪂕I��]�/��|�Ɏ���w�~Q _x��Y���T0-^�e�� u�kFx��J¾��l����W�n����r�ݢ������
r�/��9�$;UU�M��(Y���m@���Ơ_V3Lȳ��ܖ ��`C,�DbΠn3 B�oϽ�2�+��U�c���*ӤV+pN��A�2������ܘ�t}���%�n�?��#�u��/`�~¼���Jl��w���!g�|�|�Wv��ohxÛ��8�o���z���
�^X�4���8��l���%�������"Mk X6��TdrTI��.�~u{$������g���N�Sբ Ғ�,�0k9��(����.��p��s�U�S:dz� 	�R�@؇1�s�s>���:����ʒ���ϐ��%;T�3�['5+@�
 S�zn�0���~����:�����w#)Q�F{_S�w�R�Yn�{	0�2������M�'N���9�X@p6N���ׅ}s�J����n�c^[#��fYN�Z1��?�VF�>k��8*��2N��Ns;w��#xJ�%|�S�@��^(KL5��N=��8Vo�^S�&�?n�n�lԁĀ;1�����E�v���ˍ�Q7'��J��
v��
!3�iFuٝ�?t]�D��|����~m���\׺G���n�%w�Lo�}��]RB��`z3V��v�h�+T3�ൟl��K�l��	������n��t�A�ͱ��ŭ�Pp|M���N^>�]��ا�R�x���എ��`�5�^���nlw�S�6\O�]pr�w	L�9i"AK��^tѭ{�HOoJ.��1�Y�{�e��l����o�f_>$X�11��^b'b�q{�{@�/��"��o�iK��P�u��-F��A� ·�NX>,b��es�$���~ҳ�G�v,��ct=�Q���o�95ɽ7�k�ƒ���N~�����Qͳ�Ȼ�H��y��O�o��ˡ� ���t��_jI�\��\�)M��� G��Dq��p7H]��O����L\''L�I������b�)���%(g$�l$��Sq���
h��o�1�p�.�*����|�B�4�?��^�߃{>!-U-��j��:���+%EV�{lL4=:a�����-�&��[��bS�H78>1�L�hу^\�f�2�b���U7%��7_�ߛ̝��k�(�]$<�ݛ�g�ucO8�Ͼ�`~�c(j
�<�Nδ�@>X7@�EH�ҹ�Jl��涕�t��fj^p��\�=�&��@��<�DYk��djrJ�(���ی	|PgVE�.#�t��.�7mGGe�風��;J=B�qZ�PX�d�����8(�ڳ��M�c(������(��S*��:4�|U�z����g{�Jǈx��Β��y�Ɩ��a,��)���EOlѪI��"~LC&�Z���Ai���^25@��8�uN􊑺SD&��~M8s���)�Y��XܛU����f=l�A�q'㛵�Z@��^�}��o'�!V`��iƨk{k'#��I�n��0P _pHT\I����n_����쟫s���B:t��垟�ŋ�n���=��*��U����NJ ���q5��P*����n������P?�V�*r8�jI�Ç�Խ��p]g��}�b�.�Q��D�b��Z�m������k�g �.N�����R?y#%�����a<ɓ⼢x�y��8�ҦȔxy�W0,�<[)�2	�K�.��}�Ìt_�]ꕻ�*�-}���xlQ�A��/ʁ�d��.1�Kf��@?]����.���9����e��w�x���P*�ݘő�,$Kc�阝��G0�_�v8df����m�2�k�:�#��|��������Z��@�v���[Ѵsn&�㢰+�CN:��j���n��4�kz��ퟺ�l��O�u��yYC&�"&X�~�����:7r`���Q��L!��!�<����!=r﷤Y~��',G*Mdq��3}���h��ڢt�Z�6�p��Y��B�.B�r	�t�H���]��$H0����h���Z�"�/�V8	7o�d{Al�iC��w������m��ʙE�cHd��ook���m��l���Rf��fdm.U��H1)Yj���g:��#�;��t�%d{�'^+�3Pj�m%�f`(v	pq]�j�-0���>G���>��a�)Y��F��ǣs�n�P�hN��F�fr��w���.w��Tk4�K��6�L��2ݝ�ӆnE[9J,��Ի���6� e+J�޳w������@��LY(�.*�Ȭ�G��BӆrH#�C�8�ܓ�DB�6?&@55(�=�C��&[��	nb�"g,��
\�\׾)[�(g}�M[�E{�\�	-{EÖ��>	��Z�=Yӆ$Y�mP�W�)Al3��i�G�0��6�E�7舠��Τ��˝��N����D+Z�)�GUS�Q0&�n��g�Ċ�^e�4�iI�y
&�o�>I� �F��l���v�H46�C�7�6F�wE�Tyf�KX���s�գsBc��e��)��؁Ij�ķ��}���!����<J�lI'��D��؈$�l�O�E�6S����Z��2bt�je�iX�N(�B@אէ�@.H�
�v�[N*����ϻl3����!O)<jƣy���$L�"�������y��������Tn/�il4e 3��v���l��]�j�U�.���M�@����5dy�䁒�_�b�����s��2Ŝj=����aF��ݛ��6����ɺam�x��q�/mMwG���jD@�ލ���K���՚���j
��- H�%#�R.(��[�Xa͙�Q3b���aHSZZ�7��V�	͠
��`?���?���kxU��%lW��BFd|�prƨ �ĩ�*����DI{���qsk��&��C~�K�i꼍�Ϳ��6�7S��q�%�`�ȃ�:g$3����$g�.9D��;l?��ysK���Yu�nms�r�yy	L4����A�l b�=��r�I{��̈�M�u��%��;��d�ǻ�D�Y>߸�gF�O�O^� � $Gmj���#;<�-�j.	�k�hoê󪽔��������ͦ�̙�����w@P�ĝ2����Z��"%���s)��P�̾1k9��`}e
ryt�[eAx2:���Q4eۇ,)�-�*	�Gc9�0ۅ#8Pt1�	�%�N��(cF9�䂉TA6���||b�'���ґm�&�\�����7,bV?[Ҏ%�1�6�A;Db�)E����x-g$P��:���r�`���"Ĵ��;(c;��dO51�_����Y�kth��������������Jz�Ǆ\��l|�D�%L��e�$<�٪a�H3S?�7S���ѡ�u����(m�>����]���v�5NDa�-�p�w\��ڒ&���;R����ml�R.B4������]" �gE/���00��W2�Q��&Ye��iuY�Ef}��l��2-A��-����0T/�!w��!��m0�.��!�[����K���YS-�Y��M'��B�eR����i}h�c�|&C3'���z���.ϼ� ���9ʇ�׃~W�ͮ+v��o:uR�m֚�A/��G�;Ȥ�k7���A�"��숆�!�Q�0+K �:�n9n2�珧anO�:5��%�`�?��~S����J�p�	�q� ���@�g_js���MҢ��6lR?~TAPn�Q�45�w0Wf2Z.�M��W�P�L�6 ��i��7Ā.nTRz�z y��T�aF�;*(p}@��
��]]���ƒCq
�?o�$�I�jƭ���G����q�`���=l�0��Yl�Sa\z��,c�x*�����Y5a�fHo����R����,(����]�v���O+z�_a�_O�f��tY�@xқǺj\0�X�[Y����i����`�b�̱�ht�lp��k�
���QƮ�L
�:��m���JA�f�9�k���K!FX��U�	�A�Ntc����I�D����P�ǚ� pm������?1W�%r#[���?�m���V:���F��,d��ӁOF�1�4P~Z�ͤ;u���#��è�ۑ;ڲ�<'�kt6��;�uܐ�ϣ�]:K'��W�4]a0�Gw�zi��QN���^\�Yt[�Դ��0�\�ȅ�97U2E6�b2��gD�U��{��^>0bxVL0�Y��I߼G�RzTgd��W��7�&�E��+/j�R��,XϤ�_V���9܁n�	e�v��K��O��:���=�Hds&/9XF���N�L?�iޒ�|�P��c/V &�d��^�K�[�_R,������^����ҭŌ)|����L�0�N��\����q���S}�Q�a��l�Es△r��C*�g51�`8}�`ܓ^�����:f�#�C�_�n:� ��G} �Gcr0�Ő�j������J`����idE��Z}���� $%Ӏ���HA�=-<�TT��O�U�A����d��_��'S�hg�]<!X�*�
o�6�~�1��|@���<�V;WN�S��ۧ8��O�h<o�Y6�jK�)d�o�!�O�µ��l�=ENV�e�T����-lyu�r��V�CϚ�x�c_]��m���d�caMG�u�P��!����i�7�ԯ�jW�]O ������ �Q��J>���N�����D�D��{F�E��<\�&E6� {gauI�w��6��)��Z�m��"�V(\{M��+��E��C1q~����8�R�ƕ)�2�W�Z�=_��\K`l�����;�fȚ���TT��1a�'��"��;�}��:�o-��s��w]s|�D�e��*J��y5u�B// ٠L��@���!޶�rt1�}PǠm�~�k���'χh�a��z��X�uKh�;�&�_u)LWtEO�y�3��5]	ɶ;��xІ�;�;F�;f���Q�i���%�m�ɞ�r��楃�L󎅢
��m���G
[�}_Jz�Βj�;�h�<���i���^+�ծ�V�a��C$�6�IG��a1�C�D֏֟D��:u�T+ qOA_�-�Hi�oBa]bo�B�n�}����C��8A��jDלtdH��S@w	��'�7�74�c�:�@�P�>��G��Iѫ~J�U�SI�
�1��З'�����ĳ��ؗ�!�l�F�ɳŒ!<��<�L�WV�ƕ�;U~V���J�-��J��
r����ws��̱���"��d�� m�cww�#�qX?���f��h�!��WV�q�6�g@�Y�`p) �wa�^������h!M]�KQ.��X亽R#ʗ�i� C<dQ혖Y�h��zQDlKz6�@��@q��챾TK��K�<�Б;�%e��;T��
e�f�O����
����jT�I�⃏��Ʉ
�E��R�ίy����
����F�q+�k�d�� p�:�u�Sd�*޽D�Kp��SV����s���_�)Ү��h������h�Vc��p�-(8��	[�@WMY�i�?'(�q�iq�;��{bԵ����!R�O��ՂE��kv�M�m��XrB�o���:'p�����2\��r��]��;:��<A���I2*��
�,�k7�� �[5�+�.�3�7�Ǐ
e�6G��RFԖR�)IG��������������o������b0��i[�{ک�+��1�A��9#&P���=�Q�K����^D���4b��I%��<4�
x`P ��HfD�,O1��gY�~���AR�^�b(^�}�t|g��hA�An�	W�����֨�5�p��'��GR��H3��X�����J�1�B�-���p��W��n^��A�����v���{!t����F�xa0��@�%-����Cs	x�d���j�9��>#��?M�l���'y�2�ح�]�{e�Mu}�j���?���n2�Lf��'�{��M�B��en����l�CqZCq�1�������-�	�7`q� 5�����SoK{|���q�)Q���]��LH�*&�:[$�y�����@g���/Fv�H��.y�J>d^m�\-w�3�DbZ
�K�{��	�!i#�{���M[l�.[�`��CP`�g��t�4�e[/��1lB�:���+2E��lbk��|�Q&��p��U�{B�P�n� yAI41�5�F� �79 ����.]��8�����a��Q��/�	�:L,�����[����P����M��媉�u��e��׸�?���t�`��b,H�9������_UZS��*=�b�"ބ�9�;��I���E �@�MBН"�3L�'���w��݃O�~?b��0�R&o(6���*��7�����۔��칶/^]j����fYkoz?+,X����x�I �F�xb�p	�q�x�H�=p��[�,�N���>e��'��K)�Iju[]*��%��hK9���8v�D���(�s?�֥�>4`m�W?�yeS�+���ޏ)g׽��n��
z�%q�///���x)�#8'%�-	=:m{����TL��{�/�cN�6�nXj���<kc�V��rD�8Tl���A����#٢����~R����V�~~�W�P�F�W���	��>��I���@z��U�4��	{�6W#NCe��zY �.t�C�)���Z�q���M	���A���n�.h����(j
k�`n���ޭJ�-�X���2����RL)���Hʫ�.���S�Qd�ޑ���W�Zl�F�w?h5a�`�odH6M�;79Z:NlWc�d��2����s��@��]`���p*0kU�� `d�o��|��;��nb�^��IЏ��biR�f��T*F� ��L[�����."W��'�i����`ō��$�`��M�	��Kw��i��}^�����ti^-���. Zv�7�t����Ӂ�J�!������7��� ,����p�:��s0�[]wV��0)�1��O��u;�	+������n���Xհ���X�{D��������K�q]̑ߺ���l���/`-�c�l���p�K��M͛H�R�f��ig핮ma�a�h ?���\��j�H2'O�C�\� �FԸ�C@>�TYa�Ζ����瑞�	�N�ÆuVU�_�K�Aؐ��W^�~����!�<�0���*g�خ2�']=����SK
�:4���6���-��lu�,gB��ڬb�k�����Z|:���sV���Qq<�Z�����p����f�*s:lI�2�O[��'O��7��"h*J*�f�dGq͝�o�:1B���@��s;�tE����5�b��Y�T�ę���B��u,~���9�I�������/86]LM�F�P��Z���,�O���i�i�d3��
D����}��Υ���`��G_��@��A�dcUL��#���n����&��� 2NM�/
�����(7$�l�xs�U����A'�]I���H�g�B=x�Ҽk�*�DK�}�@TJ��t1%t$��X�SC-ؒ.��b�8�o�*���]׳�(�z�@��Ҡ�*Uv�-�cĆ�A�T�G�~���Ƭd�Co��>q��ae��w�h$m)JruIb��y�����E3�P�nR��E2Vk��}���(��!%�4�PO>��ʭ���z�Jx����n��|�'LX��-�<bH;�mڨ�b�ũ���l�M�?P���J#W� s�������h���i%�v��$ʊ�-�gF�0~6��ob�h�P(-9 �|�q-՝Y���)A�&�PCm�?�%t�ܦ�f4�09�lo�=2�za�C(�Yµp��S��c����nA��EM����؍yP�i��m�őW�YS֧�i��F�����㪙�E�Xf�0T�	�� ���C��=��M�Z�l��D���x�u`a(|�]�	x��<�(� F:�@g��?U��݋_t�����6��,�~k�	�1�dHz�TQ7�N�`��?��~oY,��=�6���0k=�wG�ĉ1i��lo�1y��hC��?P�uE�V���D��k&����ȜX=����������bڝ�����0H�)ƻ�T��&�icvƕ#MN0ld���!�k9�@���тz��ȵ��$���ͳ��K��� DJ[m�u{�����T���I�sg���&���һ�����<5���p���5��'	��dNs��M��۸���4�b1Z!N�ݭL�2y�ۘ ^'��Z��yò����"F��#"�t �����US!���eh�ܖ��w��SI�B*���-f)��Px���~'\���+Wkh ۵��°|[�Jb�H��6��6r̽c��y�੡�sLv3P�v-P�2�nc�A�	q:��=��!��,`ss�<k*��1���x�K�q*/陆�2�������!�X�_�|,���Q�$�|�'u��|i��E|'h9�������?�O[փ2tX�d���= r��`�fF�FL�p�E���i�gr����H�г�F奮;\�,�4�u���],�RB�]�$��;X^F�V�e�����}Y��ԏ����K�N����~q���XyCf���`�(g��Pv��o�:��z�x�� ��u�}0)M���$R�]������_��%e{�ÞR<�pB}/&�p�0&>Xw�&�x����p��N4����euժCRmí_<���må~tY���T��ߘJuQ��5�<�"$y�t_A2�>�Z� bN*k��N4�4n��pf5Hi^�+v]aA�l����NN��8�H��$PT�5��"�ܑ%���o*K���6�aN�r"���R�72/1��<׉+��z�Xe8ag �ՙ�f��^�m"�Nc"�?���I���hW�߁�� ������']&���S��DQ�meY��{�~m���w�O��\:���EI�,g�mxY�v�wJ�������UW��>�	���W�"�Њw��&�u:�-ja �뻕M��b��7�Z�a)�Z�~�M��h�-���5HB�3 ���M@K������$T�Ͽ�|'��E?Ǝ���F5��s1��Y($,.�[��B+g��O�P��S�df6�~q�>����jn6�Jw�lb�$a˒!�a��F�����Rۥ��C#΍����M��
�_'���tU/O=Z��9����{�~����3�;�^}C�Bf�ҙˎؒ~���m����*���r8�hm���./+!,��Q�8�l �I�v@_�l(� ƞ]�" ot�`.�\�>��m�j括�I7� Ⱦa��ۏ5��%�ޣQ��h����꽓���$Rb�׵[e��w���P4Iva�'nPt4��G9�%��۰U%�fJ�O��JT]���� �&;�6��ʯ-"�_�����M܋�,�i� 
-�a�:�Y�߻�3�d-2[���aqT��p�
����kfi���c�-��`=̫��9�/kf C*H�:G�l,�X��Q�k�O�a�~$y��[}9�?��)[�C��]�M��j�l���#���A"����A
�w� ?[�������`$���g_��-U�\-;����*��gv ȭchI3�N8HV�k����֮w/�1sa�X9J{�����a��?�h�����$��,�1\�����T��Y=�pa��`���Rm����!�������� ����X�e&���ؕC'!�c����|_>`��c��s�6�p�5V��7A�-�_�|��}O�����+g?�2$�*�ȲD]�];�u֢�ݟ8]<������Vb�^섌�3��n/ƣ��5	*l3�([ V�H@������J�Q��-ml����O',��Qx�坫�}�7��x%`���B]`u�y����P�Tr���/�5<�r��W|
���ߡ#��)J�E���5�]�A���X�Pk^�|��e����?�vY�4n��6#�gqIQ�r	*�#{�Q�rZB�Dme��e"���R�`�Z��Ȉ�;Ho�_�\$=��C0��xA��,��~s�k��6�إ��n:��a#\CФu�j���YP�Vn̦�ˢT���_�%h_�����6}�;qZ��]ݎ�ߐpN�y��l�2=�`�A��������#��I�H���e&t�C�n5�y��&�����)�x���q��Ww�ZY5�ld�X��u�5���W��ֹ����'����2�Z���Q�;ϑ)����d�Y��)�W�M2��s��?��6h~��ί$���^f�E-i~���f8��ùKOO�#��O($��9�BeV�_Yb���t�н�������2⮍������0Y6r�p�nZL��^i8�c^�a��#6�G8ݚR�uw��|� &1J�	ؾ_�$�[8��+n�� �5��Ʉ�* x���ry�q�s?y��z[�i�NX��p���jE
���E����t��25qH�]`�䋣R�_�j޸���
���A�OɊ�Tm^t���4�t�@\�t�*���r*)J�4�����|c���7��*��`��`Y��H�gV�����UV�+��+z+�<��y�������+�W�t��_qDi�$p>w�~ɐѸ8f:��ُ��iű<\�Cb"8�c&X�O9�J{�#ɂ���c�(��v��gO
�"�zoJ��{����&�� D9�Hh��d����m��N��p�A�/�;�L��|�ĆREg:�N|��&�Ѷ�)���£h�C�];q��b^^�#�Ev;��شI�RҸsO1���{�T�13<]M�ا���e9�u�haL{�>�$@#ܮ��)�U���S�{���l�������kR��[��KuxQc�q�Ʋ�6�"L�3���s��,��u�w`�b^ʽ�E�~JVO���O��m_F�E
(%�p�%Y��L/�:�K�1�3�<-��A�.uH���i�v����|��G�6^ԃ�X�_~~L�>��W�)�
0��?+�c�^��} �;��p>����a����������k"�k���R%�W�$08U�P:�@��@b/�;�0���4�Ƥ{4e�3]���y�N�N����l�t�V��l�{�H�� $�2���h��X�W6��r w@icNt��O�f�Ǚ;�֔ҥ�W۔�w1U~,�$�߷]��TWW�|�@��J�K����JZ( J�X�*�����!"�88��ܑ<d�Ā�Ƃ�Յ���G����+��D�v����$�>�]z�cGG��y���G:t���He�>�0'V[��~zҁ�D�>�Kz���,�K�_�X��e�>��c���)X�&!U/�Q-a��tg1�OZ��j*�
1T �\��L�r�j8��N�([w�B�|ya-�i��ڑ[����������d�Z��� S7qXL������kjE��"����Ǿ�S�c�I~����dQ�T����-���M�E�������7�֒'*5("��k�":m5D��H�j�LLw|���(�JцW1�r��!)�M��	����n�B�ՍF�^��^}y��z���8 G��d�N6O�=Za��8���nnIXq!3��&�����A�3`,��r؃����!Љam	�B����_(����|����b�i�d]���F�'��BK
$V�7uC#En�qm�o�&͹){U�e��uA�0	�Ymi7�*�@����
$�LC�Nyg](��P��ӪR�ҩ��u`9=ۦF�o��Cl���XP��j�_�"�:Nl)J<�ҹ�_�n�w֔�	��\��6��qz�r2���?OMLk.��+�!��^���:V lw� ���G��q�ؘe��n�p<F�c�j�`�Ou�o�-V����q���� ����X�j$E���n|�)�J�����a�^��Y�I��+�L�4,J�D}�c���a�t�h �L�� ��8CUG�	'�!�z����Y�V~F[|ht/o�1?�v}��&[)��Z�;v*fٗV=
TA���%�nⱋ��sP��K�K�JZPD�������|��#62���ժU��ꍬ
��+���-�}���J5��2'�{��Y,'}�}�V�h-+��z�춒�L��{�+t��6�Ai�!���V�*�=c���3�x�X�T��T����T.�̽2�!,���?���h�&�竽�<.��Vsue���ʊ��:2��epjO�3��������^�O�ai8������d�ށ��0�-�� �R L���܇"���'���%Dz)6Ow{&`�p�	u�0�1�
v�,~��(X�&yKX��E�CjS[g���/C4�Gn�Hz��C8����wR �X��n���Qps�#�a�$�KO0v�a�LlnZ��֯���:ʽ��@�m�6�����u���^�h�7�,U�9��n�Z�	��G�G�v3��LjB�Ag���-��W~�]H�??���D%���&�Ku'��HӔ��P@�,���~�MZ-o�),;���f��QqP�aN.��b��u���yi���E����9PR���Dŉ��\��`]l�z	��4�b�vب@�f�Q9�xƇ�7�eK� ��d(�C�,8弣�}�t�r�h
�[p�Ȃ �F��O�)�XM��R���x�j�R�ۛ��՞ȠI�C��k��T�#~����b�'��!��b|�ݠ^���p��-�`�v�v��\�6u�h?�	�@㤧�ɿ?8����DmѺ0a%9����0-��̙J,25*]�S�9����:W��u������@�U�K&�����6�(���D" ؉(v��y�*�_]�&�q��D�Qy���[�#//�����RsL�+�G�a����҅����]S��r�Z���$��M῏���0���mՀx�\��a���G��:��DТ��b�!a���v <dSãK�b)zj��x7������-Ʉ����]gi���/���3'��dfO ��R>���vA�Q|���_91�B�x���7����Wa@W�
����6��,�oP	��}�+����ܶ³���G_>�1����V��w��'!9������1.x��$�Ef1��b��bk�ݕ@|%���tp�`U�]���{}:&	��z�!Ʀ��b18�jl6RŻ�0�"y:)ߴ&�	/ Ӑ�G(����l��]��	�=�m�������d�aQ����0���#��n���6T�mN���1Yİۡ4j��O�{Pu)���zz���<�M�[�H�r�=�!z�?>�#>�_6,R��Z�>X%�T��-�+S$��Uj�v�:��t1YX��F�M��7��R��P���Qݏ���2h��"�:�@�<����>T\W:�4n��MT������
� ��5B�%��NV�=��?f�k�����#ɳD��|3�B��<^�+iL!-�B����e�]K����.��q��M�nV"1+8��
��!�E��`+W��3nRs�D�2� m�H���C�b�}�a�q�c|�c�	$C��!��>�=�X���/�G�۵�&F*�ݻ��s�ރ���PJ��h`3>`�T/+ǼEj돑�6���UQb����l�t:h��,_��B���Ȫ�>O>p/�����Y#�8 �1Vjq�+⢦߀!V���L/L�>��A��`�;&#�|� �u�K�����RB�x�. �N{��nfxڌ3W>#P�nШ�mVx�71M����3#\���p�[���SF�Җ,���M����؎����:B�b���b�Nt��R���n�w��ˏ]��jG܈��P��(F��G÷o�g�/ȱ)�,��i)w�:5ϴ�.��It�7�l'���J'*�*����6�
�r&�5�!��\�-�lPk�g#��ќ�Iy�����p'yM��4����L�_�K�s��[��![�K�I�9Uw�&�*�z�44@���F+�b�I�a���|���\�R��:.��r�@c�rX�ᘹ>k{99*zY��V��/y�Jr����k���DQ�'�ܞ���\�{��k_�r�`qsU�ڦ�L�74�=�j�3�����/ZPLH�<����%� ����N� B���fds2��fK$�F]e�V�T������8�\����L��^YU�P!+�'� jݚ���;'4�"�_��D�;X'@7��������׆��VtJ�<>��*$O�n�3x:�AI ���F܍�?�U[¼�O�X�;Y���W���1�8&�6�I@gD�*�cm���C��;�-ACH+i��h���7hˡ��M儭<��(��ќA�������(2���7�(��4=��_%Y�tV���
��:ľz�j�s'(7v�	�`d�'C����2`��.�* (u:ؘh�׀,R��~�>�#�U[kH����	o2�;A]v
�J�Ĉ'�u�4p/���l�?�Y�	���>,]�D�6�"Y �6`�Q0��T�pB�w��#�E6]��ET02�������Kd�e7�D��[�D d��m���r�vU�$Awc//?��n-�2+��7�+b ��sf1(�E9�AM9Y�����ފ��~�����G�bc���,�{̩7�)�`���z:nN{
�A���$ogt��>j�N__�eA�t�%D����@�l�67���ذZ��+ҥ@4����nm��A�Ƒ�p�i+�΍��Q�A[Ϡ�I: 6�p�E��^�h�,6�3;~p��UB�����i#��t]��rwޘ��G=�lMGL�O~٩��}�=��<Fӌ��o�����R���b����W���R��w$*�r�O#J��x���`�#���:�T�cd���$���s�Q�ݚ�����0e��y��u+�"
F��|����ty�Iq`��/���.��ԆpU�1ܚ1]�1Z���b�Ө6J���9t]�g�K�� �L�a;�$��wQ��=�t�9����bQ~�e�2D�͙��J�D\����F+��R(x��&�<��BZ�����Z;ס���
���M��Ϳ]�7��-��.�?�/���5�o.� :szɿ"ݞ�dҋb�kFu5�����_�m&I>A08Kڳ�]�9�X���[�Ն�c\/��|�fpѰ9�:�(�I��u�>(�ݓ2�ʫ����%�Rl����P�pO���7y�{��`o��6�O$�PFcݝ�qR���b0��+�<rq�����.gb�K��\�.Ϋ���)+�?�H%31@��s9���=�V�<L�e�=�}��Q�Au�WLޘJ�3��3M$�4(����hҫ1Ϊ�ypgi��E����:�zJ��jΈ��m��H��	�p+�ğ�aY�c^���F�����s����Y�_��O�9�,M0��n�¦����t��e���΅Sx
�F#ݪ�i(6�#O�)� 8f�yV�ˬ�+[h�nh�z����JA�5N�
�-��Q�v��5wĄy˓�&�P��~1ֵd��\���Wz���o�[�]�mG}�	�4�Y|'7�S-�D.Z�,�]��:bdaAG(�6�&dV^�=������Od�����n�եW<���#�>9���%��6�4è�G�s�hT�ϜW�rE6�ċg��02��8C���*����n�da7��igP�<й*�k��I���]C�����2��Hlg�����7�����!������71�
�N	��+
��7��v?��w9�֠}�*���Y��]C�]L�okL͗���r��h����*�4���E�����;��~��`N�8��n흩+��G�p: ��5~���Wm����0���ݪ��d����g��j�g��"fA[S*��՞���B�Fī^^�D8��O��s��#��+-AM��dw�����z/�;2�w��N��Ԅ�z[�riB ��#�$&T�`�&'e��G��}�]5?�TC�������.�rGK'�@��_�������9W�$߱〥��g^���&�&	�m�T��I����黂0'HE���(z�)�@Ef'µF:�JBj����F��=�U^k�'�CS�� a��I��k��i����בw�0:�?O�=8�������~	��N�[*�¢�"�d�?���.\�A��@_K��"��T��XŶ3��l����iCe���a"n��չDL��O��p�Ӎ/bp'][׏� U�Z�0cQ�*.9�����E��������U��R���i�����e��9*��5��{�y�D�q0�@�cI��T�t;+�K7���8�NZ�P��;ϓzk�}M`��\����P਺��c1�X��m�]�g-�N�>�P���t��=�4ǖ}H���/�Z���R�61J
�
�Q�	lGA�LJ|h��k��#����@�vԬ;�#����ӷx��e��"���b?	�OH	y���z?�M� �������ڂ|9�;,{��ԕ	J��F4M*��DV�z,��җ̢����}ާbV3eӣ�H�4�]y��4l��Am'��mw&R�t�?>K׏hͿ�yk��ʃB�|�{�����?�p�8<$z���G�\�Ե��urMK�s�'ԛ��,U(4��\�����������H��"*RD ��(�4����:���8��W�Ž�ŐB����P�A�����uc�/���Hn����ɖ�0xY�yϨ��BU` /[s�l��x��㴦�-H`��[7��0����r]#�d�S.���lv�چ�������jn���v��&���P-�@� �o���_Ҵ�Ð�����\ɘS��� ��r]]�oV�+H�c�(Fy����(��<F�{�坲^�*{�Z$�UT-\��L��S=�-	�YE�R�\��u��q;2���]�'��Q��#��h6����H�5��k"M�	�H@��b��F>3R���+�c��a�����������1m��]��=�8��� �S�QL,����3(VZN-8��Qlh�l��9g-�h�9��H�&R3� :�b��@��=-v�0��c*����̅�s��"�#�6RǏ��(aSˁ�<Q�Z }}n�A,�O���{�w->�1���/x���J��0���X�v�m��f�9q��d�D�!�e+2	[�i�"���a�$M�y�����Ah��)>����������	p{M��߼������ˮ ��5Tp�-�ci�;ƞ���/�dB�_5�m��Ձ�V���=]���#I�ա�jM�6OZ����J'�c(ꚺ�hA�0��R1�_��txFʉ��(�~ ��xͥ �ƥ28ā��A�Tߡ�F&�d��J���
�t�G̀�3|�z�:)=�-#)ͩ.)OՀ%���>%-ӥpe*�+L�[-'�=��1=�^��yJ滣(���'|y!_�_-;��b� �4aPm��Ww:/�Ѕ㾡q�I��Ȓ8ZQ=� <���=8�"_����n���m92���ȗ�m�������m�^���[��-���!��J�F����qq��k:i�3�!}�v1}�X�X��/6xe�bө�rF��j�;FUM!��Aa0�Ez�����z/�ṳ��lQ~	����Wm&t�M����n��P��m�!⍉G}UGl2d��
O���f� ����v0g���;6��(䎺��W�KMW��1s�O*)���>@*/���jb̌ݬ;& Y�o��T�S��.I���<����X�׭NwC�25��o�����*�>��kM1����>`�\��?�f���q��2�N[�Ő��e6+��4�(��G�S&�	���|7[�r�ؓ
��
�^,���0�\d���{x^�y��{xT��Q��qq'���f�y@q�i;�(�n�s,�p�x�:�,���UIxb�WSݹN]Q�A`�$>)�Ÿ���
YT�9��tQ��-Q�ʧ�5�kpS����o8�-�"���ڥ�kP�W��o�X{���(�)��^�k��O�?.�!���(����ǜ��߰j9�c�t�C��%��(����$u5e#Q�;�"x��1'�v�3C��s��[q��[�+5}���蹃0����V)���d���s���!\�"�Z��w����Ld5�������� �FD I�ib�0�\!{�p!�@��"��G��1x�[��I�]�J��A��r �D}�~�2���w@dj-�i��{2e�;V�����K�0FjNՙ��6�c�^J���L�0��oH�'��m�8�5Q��G+���3N~4���!�9�c!�;ރ����渌���-��V������n�:1pR���RDӥ���9r��������񝰚��<j�i�s����P��G�?�T��!�{^�,{r�p��.�C�O,ʄ�G�L$&̙��զ�T-�ą$�PF�UP����lEV��g������O	�J������@",c�e�&�ӓh�
Ƅ�"}^^�˒��K�/�f8��I2�60�E����/���FS��[|��{��m���H���f�k��+�!7b��qS�&a��pDA]{tZU�G5(��V�	{!��JAD6�X�xgOO׀n�}�+��#P0�)��2����'����˧��.ı��y���E`��Ti�l�ϧI�l;uWv��?�]��ىwDu�v��Iu�
;࿚������vahX��\��b�}:�P���8?�`z����m�#�L�kI������$���3�/��·e��,E�6�2N����׻���׈��D*���b��G��c�r��G��vȪC�����>������hc	�����{|d�������Pr��/���*��7��!Og	B�5VR��ϼQ�	})l �iV�C���Y�
a���V<��`�����1�$��RA�(�ws�2(�� ���u�	��rą\#~?��.�RpPr�&�m��:���>�lJYуYSfQLwD����	�7�
���],��90���/'��EvƠ_�(z=��s�ե-��F�b���[�����D��2�4(H��Y�`6��Sn0}P��IP"������Qjx�����渕 н��1	�r�|���J�9C^�0F]� �(�b�Ӆu��9j�<�G�J�
&���z0��[�ݰ��3��P�F�R��T,�#��V!@,��	?�4R���%�m�Bk7��s�4��x��J�콆��̺���c�����ė�=>���r�J��	vhq_{=&�d�$��n%���/����lZ߹��9t��'@�(~�%�Ԓ����LBml��q�\q�sr̫�<��cC�J�^�CR%)��]��J4rj�٦���)�<翔y��$+Ig����hz,���n$�����bH�R%:fI
�U��M�[B�a7��tŒU{�oH�y#�g�cP�� G�X�bj4�N��r:�~�Pd���,���i��B�$f	���q�|О
��l�f�����<y�=a�=M����E�������Vr���b��~��:g
�v �(�];F�2�xN!*%���HU�D���~μ�|���^�[��#�����*қ�[;BX8,%�>�q G��HlbZ��s��~�=az��7ԫbI�9�G�F]j�ѓ��r"�q:J���d����qy����Q�f�d�,����5ǘ�J�&o+�V��y��s�� 8APU���@UT6q3�:���lp����+v�+�����&��?Rܐƭ�2�k`K��M}��T�q�]�fJʎ�;y�(u�+Br/�T�����bM�c]o��-�ϑVNl���WW��q|�z�,3$G*�U#�iK��9"H�^��l���|)S������)`.�Tr��z1�����3�B	s,��`!،�r(���d���J�A]Eee2��9m)J�������7v�N��L��_�ƚ��I!�ݙb�cDiE�y+*�hA!Z���x��g��g�gf��pyI|<�7nߘ\�K���|R���O�CL��Ջ�������?�K��E�N����@��t휓;�"᜷-PYTcXvI<���B�g�����<n���(��� "�����_L*7vTg�Uv�����i���P����������~��)�y�Z�!�C�2�t����XC.W����T�^A6�x��$rDbv� �2%��M-8��Hc�����9�J��A���=�fW&x[��`���؞A�4�4|�pvOKmT�]����)����5qjP��4�E㤂�v���2�UDX�w��SK�/���B'k���"��Lm��G��W���Î�h���p���IE}�y������!d�*�N,��f�P��E͡~�{���Kʠ4��PN��>9����֢��B�.[�J*��O�\>\�H�謭>���piR��2�Ӭ��Z\���iC�3˷ʼ�;�.
�b�P��K��&[����A��k�z�N��_�m��b4�"�0O� P�[�I���ҥ�Bh��ӢeO�<ݏ�1$�_ͤ/J�V��rȴ\�69��1� R
��E�D)��S��C���3�g�|n�����9D%׆SD4�܏>��q�\n�W+�'�c��g�8I�߻_�ǯ�٭��o�6D��y���3O=^�������@ſ�� yG碴8���)��<JM|������S���֛�esG�'WV��/�����דW��e١ 9^t�Pu�EE�k�'1Um��1v�K2���4ʜǼg�.���}�{x���)�Bӧ׶��%x)}���L,ܟ�>`�5�$.@����>�%�E���F��-Z�C�]tkJ��6$?�s2Br�T������t��m�zK�ӣn�(*�9��0����	��ɕd��ӧ?o�~���ϡ�T�E�l2�yd=-U�����8�+i��8��a}5���;���Ӣր<��b}�"I۷O�h��T�#Ν�����E����Ǔ_�/� �z�v�@V�Nd�>�ߏa_6�H�rJ,�hX��}G	X2�z����km;����}6<K���钟�p!S*�b�n����[�C#�^����y���Q�DN�[�a���5>�_�O{�?���b�ZŶ� ��2+@9^�ݢ�O���+xf�RxB���Ǭ ̓I�0,��ZH�\��Z�9IO���
1,!=�����`|�/�;9ÜOC>.�XL�fE�<�6�V�Z��}H��C�+��2i�9ѕg�0@��^ J�J8�B ��+�_�f_�����PA���8d��,��D��(#��^�v�N�/ԟCr��?V�k��r�،Tl.?K��"��ɕ��;1���"Sܖ����g��(1`�u7����5J�X{�ފ���S�������uަ��
����g������\��ס�(�.��Sc�ѭ�0�؜��'����`�� I%��6%�$��}�m!&Nm@�i��\Qw4�PSd�;��/��I� �eѾ<�&Q���ps&C?�?��o.��e�T2Et#��=���2B�&z�Jҫ}���5?ks���� P�Q���9l��g�eF��:`T��R�|�Ra7��3ޮ[nCq��M�zLdw��x��E�4��b$ Ƙ+o'�ۮi�Fo�����`����AT��T�`��`BW�}E�h�#*ov>:.rK�ߌAj��B�h�����r�qV��$��;�B��\������;uң�՚��p>>ԩ�Y�[%L3�[�"uO4b�O��qW���.u*��g���:\�x퟊7O5\�{/T������l~,�2�*��q�nY���??X���}P�l�[H�%�\��dS 5�g�_o%l{����0�����3��Z��#����݉�z�UU�ūS (;	�g�#��[3C����I��ed6�M@�`��/�������E�X^jP ��~[wZA�!�w�s=�A�����ˆ�ϣ�Pl�EQ.��r�L�T0����W���x|+u����(1,�Y:l�d��$i�:�`��A1{�ʈk����2?P�4�L�����~x��?n_�;��ɘj���ї��Q+�cg'�˄<n{^N�9�fVv8�H#�n�T��[}VAF�����JE�`!ϊq�u,�5w�.�=f��yt�L�B�aS|����t��]D��e����3��o.��q?���kg�ߨ [O3����p)���{<�P����g���֚*<�o�Me�q�y&|�S���
���ϐ��&4;����X,d&C7��̲�����%�����>��*гt�{ѹ�ǆ3=L`�K/�-��M��ڀlnc��y�1�,�	��n���		��ne�����r8���cTJx�M�^�4������^Ro��M��h��tan76}_�@Y�v��Q��� ��I��-����%oF "Po�C�^��4�2��pв�HU���8�ӛ��<JĿS}Ɇ|զ�2fhki�ϯҳ0͈�8���|}�0������%b�?%�ߵ#@���.��x�p�QWK��e�֖@�Ն\J�����enL1�Z��6����;���zF{h���B��y��eKyjh���������D�S����"��<�>9������^�t���nD������s1H����S�/C�NZwvq��5g�B�����dN�� %��}8<B�B;��D�P�,GX^�8SOK>8��")���B�YK ��f}���%��Z��7�p�o�!S�*Ф�7#�n%8�E�մ�O�w6nUt `�Wַ,B&*�v�n�6�4[�����ΗJ�b
W�s��`[��j�'��{�v�F��������q����k�W{���G��"Eu��~�t�Uy����)���������k�N)�,��4�5)�sc�Pu_un��:��3��<t�����,0��余7�"��흶;�Q�zu7�S$���tu|)/�t��@\
�^c2UJ*r�+�ii�*�u�v�����/1��C�x'Ck��-�;Xuή*�0	��1��v s��B�0�$��?��K����2腝����Tm���W	~_�P
��
G\�.�?���2�7���H�g爁��i
ĭ�����P��W"{2��@d	R�Օ���K�
�]���ŏ�[�&>��҅���KD����`�Al�&*�R��Z'\�R��'�{�g��H�*M�k.���������	�)�P�\�O��2�W!�����4	�-"_�l,���ĵ�1�6𷌶���Մ��Ȇ&u	moQG��ٵEυ�)�`�2��z僇	�G~dRI�ϕ�O����~�����0��!�4Γ\��Y�e�X�l�>�6C���K�^�$W!I%�=MB�_����&XB�^~�L=�6Q�g|m��LO�zd�Ô_�^���7�䊓[יT]���%�c[��l[yC��ʮ��@�l��pi�v
��Ʉ�|��=�Wu����J�K�:��P ?�� Xd�:���Lg����h�"ަ���h�.&2��r�o}�"`�S����(�����!Q��N|z���!\ٕ<��7e�4�cZ٬C�=����r��}�a�'�q{kD�"�.@���"W̗�̰?�g�`�scp�ۄ}?+��z�-$������~��8In~t��	�ȁ�2e��+cc�с��ukN��,��FP3x�\S� �9�Aj��w*�ԟ�)�P���C/(���	��P8��MH��^�۳!��u"���q�ͥ�Hn6�m��y	�03�	Q�Cv� �k�ڗ�X�y�R��`7-d�OB�ͷLl��?Z�1Fi���̳�m���׹�4���J�[b_
���IE��=yN�^~{���]���R���LtG�8ȇ����ʜNݰU$�'����A��r�Z��A�I���d��W��|[s�'sa����r-���K�xKyO>�)���ߛ����r��+�/��r��p�a����M���l���R�FFB8�v	�D�[*�~}S#�|��`��$|:"��iD�
�M��YU��ߵW/����%)S�S���#�U�?�.�%�r^R�B�1끚��d"ۯ�����?�@W�
2N)�?1�)`;��|��zi��2��[��u��ւVb���D���$�x���$)Bn��ݱ	��ZQ@'6�-�Y�F�/ۓ�~�g}���%8"��H��'Sr$��j&Ȗ���i<�(������P8dR�Q�wX��x)n����̀EHaN��F�e�X��6\Oލ��B����*`?���9�<_<�wZ��҄��b��8��ky��.��?�r���������ϰ�ҿ
�e-�=��w3s�R�F�$Z��N�QΜ�M�V��D_�6a���5J~|ԏ��)�d���W˺y���\��?��ٝa4�8��/��e!D��a )���B�_J����˷�l�[6�<wÏ?�I���H�p�H���W@��Pʎk�^�ӿ:�yI���6�%�a�bM�h�iT�+60�]�¿j��㘷O�&T�E>1Ľv���acB�h�2葋!�d4	�M��F��0rZ�y���zz�0�5��\0���d:�(t��;g5���>Ѿs/hhZ� �T����K�y)��#��p�J^h94PV䛢��`��J����Sä��|�٬����ny����X��kl-~�R��{2�.:�����=�@��z����t7*B,�t��=O� I��OȳM���z�0��t|.�^jq�e�IZ����dc8�l_ZG���0�	i�DFM�Ď 1�B1c��#�*�k�UA��,2���gY�g�"�1�;�8��&���(���iM���6Z�7u��GLۍ����V�c�4����D���]=��"���;���G��]0�2��m�'p��5�Jy3J7�5?�W�P�/�G����K;{�`{|�bL�nmz`��%��=B�ȩ$�ns�3*E_�f��]sC���}p���*�{���ѩ������中�=-s{�i�'_<�CO͎(5��.�m)�B!al��]�{p�sa�:��F�\�����nq9þ]������Ŵd�����,��%���k[�N��9=	��J� ���� ���żz�%�z�W���VV:�eR3� ����]�!��BEZ�ߤ�9M�>�&��"���b�,�=W��.L��8��K� ��-�d,�������Dc�?x4�Ԥ60"r
� ��&�F I�We-�8�	��`��z.����a���'����sG~��9�󻗇g��[�>�).Jt����K�j{�p��ȯ��e�KȾu?ER�_,�����<|^���v������z��Z���S���0���W�q��(Jh�"oN�=8 ;|�p�f��Qe-Mq0sJq����I@*���Ѓ{�4��Ș���Xt�2��v�ż�Iŉ��GD��	Q{}���1�9v�S�Y��ۙ��Ŷ���k� �;jgž�Q�f�Q�݋�!��B����*�,���V���l]	Js��ُү���(�hwd�h���^^+��=��*&Uφ�]��9'�5�B5jBz��H[[��In�̴z_���}BDLѱ����@j[�xg }�#/`��'��SO��e�w�4;b�z���{�;�0g�gY��l,#0�k� �;���Q6+>�Fv�^u�xLW_�������'�xCXb^j��W�&L�6�E�He��?�nz.A]�d��Rh��+����YD�.'�H��)��lgom�H�G.�Z2��!@�h�����֙���M�d�a�^�5����E�# ��f�g�v��~A�v���暇e ��ҧH�Fs�'TKG�{ɝ�/�g��5P�~�&�X>կ��tX#=�U�s���PvO��$] #�f�h`_��r-]N����B�
��js�"�=�|� <��&�Gr�����D �Ú7��VϨs�O��`7q�|Ͽ�&��$��������k��G#�"@�?��+V�J�x�y#7�7?����֑g���!���gm���N�/�~��:�pRon�ᒜ��I�n����cM�,ݙĭ,�`>��X���J�[�16��~
+j�������$�GHg�v���.����m���K��
׺A^AחAW�-<I{o��w�'�0p[�U`���<�'�rx��zѾ�l��i%d>�j~� _2(8�5YZG@˻����y��'��v}��­���@�D�/Նz�fM#C�7��F���G=0��7�> ���3�u��r��^��0��������6]G@D[��9������H(2ŚL]��zD�8��0��0&C�_����H�:�(\N��`��r���Ӣ-w޳�0�g�5��#��24��t��K8�Y��a����z��ajq䄻?��$2��j�͹�Xu���r~N��������tfe.�����$�JY��r��=�w -��W� �IP���=�V}t�]�g1�6,����؀�(@�|���( �p��'�~�#�W�����pv��ʡ�LBWW6c�)rPcIf��˵j�ü<�[Op���׽Dȅ��MRk�=��X
]��P��lK��W�����G�co�:8˔��-*͇J�����݀��/�q	q�m�͒���y�A%P��WQk�k��M�yB.C��L�'9~W����z� �7�9�jz���,��Et�眅v� XY���#|˄l�fP\�d��DW�R�01U$��)��aO�ܱ�"��r��}���O
�	���h�u�jHң�bm��k��_��΢`�h��_�ph�EK�Z���/�R�Ac���n���PheP�4PKWPzWTOP�'����`�$�=����%�A=��;:]���x/�_���ô;�8ᑠ}�m���!�%��ּq�?#� ������Eb X��:Jt j�$�10�� vZ��M� /�^���`G���Ӏ:|�y��1��|%���ơ�%n�j�`��;��q$7g�[�@����@��F�HG;y7Y,���G�v?���58�
�{���B8���6u6�@�ז]�f�ց�G�.�2Ů_?��l�9���$p}(+j����z�W Y��6X`V�g8:�x �=*�BJ��@�XH<�z�n� �E:�W���[T��!�V�<\B�7� ��5$۝%���Z���ǐx$��7{���rRn���|����ȍ�s�I߆���<��V��Q�[_	kNO�x�ӓ�l��uv�ј�"�b�Ԑ�2�oOD��ϴ�k��]��87���p��/�Z�4<x锭��ٻs�%O<�+�����x[��汀9�Qĩܝ
Uq��?�2ʽ}�(ط#��D���4v�^p�Չ�}wfe�J�5[�-W�{��?�����̓p�6z|��KV0���|l�%�y9��E1�W�ٛ���p�>D$�R��H	��4 ��v�G�jv_���� ��r�XU��9r�^�����C �բ�Yh�
qK��l=M�3Y�TZ~"�{bP-��Z���@'��m�=�x���7x'Qm%�.LQ����/���ۢ� E��/1����kS�E�v������V�r��pAL�n��Do�͘����}�!@��S�76�@�@T.���n'P�m�O�VB��NM���-#c/�)5�R�vCfU|�mb`|�e$���a~�~�kh�n�1������ۊ�g�F7��rq=���=���xt���]��!��a%"q\RE{�w�*���ٺMg�+�j�?l�d[�#���B�*�ל,ߑል��u��?��s���m>k���Qޢ8}!oʑ[�o�m�H�+C�~�g�R�n����T͝�]K��O�mʵ���L�F�$��\�d̗�lJ��^C�/mvq������*x$e��e�O��a-n�vU���^�>�mC�<I{�{O�g:.�D��������t��m�� �g�؆#�"3����'DN����t����e�o 2&[�8.#����π�K����g����Yf���6��-�.��b!�!�����S#�X<���׀I���%��,=;�_�����YS���J�;��W��YJ-�����_�����`��o��d���~�U��v��[C�|{����c'�s�'M���ι�M�>6����ƞ=�������f��[��p��I��S�6��:��/�y����֤<�(���M�&Mռ�Tl�s1܀����i��׷T6��-C�Z��W�#�(��o˅>פ@�x0���3l�5��۬���O�3���u;h2�}��P:�u'Tsp��-��%�v���iM]��-�u�~��z���$Ȧ��¹y��_*�B�;gx��MI��`E�ݗ�:�e�x��-�?TJ2�d��aç/�f�����(���86�7����ͪ����(��Q�8�J�:����a4��s�V�-�Oi�ܛ���*N: ��Q{�t�Y�`#�Z�(�w�?5)N�t��L��B�RK��3�:�	�Jl]66e�{3*3�0�&.-�_<��`�dx`�Z�� ���q���OL��-tX�+g��:J�ʤ�n:!�9�ǒ�\�[�}Z��uF�2�� �=����u3؅�8�`^Z@�����h�[8;xn]�u����<7X;	��$�r� Mn1v��{���/���}d�W�$'Z���o���4��ovɐ�<),���Oċ�S��.��y�ꋿ'A�s�jB�썃�Zh���a��LQ:	s`�����R�5ggB]��S�ݯ4-���9��:!q��qⷯ=��3F�t�()Xg�����r�&*�]�������cB/)Φ��k�*��t��`����E�/�y^z%���B
-'�3/l*�+��O��3�:5iV���3b�y��A\�!�E�0"Q���-F]�|��%aM�J�̠܆�Y��=�z4bp��˙΢���g@<����w�u�.U�tu�a��z����c���2�I�Uq)A�=Or�l�1�"�Ċ�0��R���.����4��x��ƪ����7�T�KnQ��[�~/{`�6�`>5eO�*����O��|�����Q�S�J�I�������?kt��ja��F��:�$`z����i� �b����#��C
n�	'�����Oc)��S���ӱ6ӵ�]ڼ8����+Tܲ�v�X2��G������L+.�8-�N�>�;}���}0˛/�8,T_���t�5��R^��6ϖAȆ����e�I��P<0K��M�i��(?ؕ]+�;"�,�0������E�ɣ��|FJ�OE��T������ň ��Z�CuԲ�	��z��}_����^����CVFR@)�r�S5�~��9�� >��Q�jS��Y�ҧG���#��@��ΐ����aQD�~���a��G�Q��]K����v}�̶���>4#��ӣ��wq�Ea��wf��A�a�����@
|���݇T��G���Hx����Ȁ.�=#T6I�Y8t0/7Qg+6������K�V��s忓6��iaz&�]'L�������C%��Ӡy[ܝ!�>2�O!�?���{�|d�.�?iJ�Y>�pَ)-e�<3l~��z��X?�y� f���[�S$��X沙�8A�g��	k�qt��xy��z�������j$ݥ]@?{&��(9^��J��=� S@X�w	=����
�+#m�����W��z��*C�(E���Z�~��J͒d�pi��p��O��	�<�'�L�*��� �b���M��a�rZ0�5���N��jh��.�śjc�/��u� �<�a�5u�6���✡-n>�ɯL�V�  Ug�*3�m���?��.M�G'{%�y�49��R����T�H		���5x �0���`�M�uD�Lu������b�N���Kғ� ��K�y=���/��h��L=S�(�5����J�S�~��c��#��|�&pH���NSŭ#.e_[���*ӑ��E�جo|�2�hB�̨� c��{C���??L@KOI	� �p�
����Y��W�4�v6o5ȯ�7\�G��9WnR�1��5�*����L��!5�Ð8l���3�fj��v��/C��k.҄z�6��Sw��zoّ9.��Y�0*���(#"9��`��� .aS� �I#�]�l9R#��*�T�ٗ��-�@�f�%S�.�H�nIk�'\RXD��۶�f�9��C+�Y'����'�4�f����!�P,��׀����U�Ȁ��������Q��?���]�\�V��:��l���^�o�-���r�lw��w���n�(T+��-d���˗n�|$'��+��
D~�7�.��y��.������T[���+�Q�}�܂��=�n�/y�Z�.T�.�ߙ9/��ѳ�5J�R���J(O*x�G���?a�$[G��
Lԩ �e������F�,�g0���C��4L&Cɘ)�7���f��"nVQ�Ί��J�e�E[�+���J҆3�<�����.�4z��g���w5`�nz���_g]���Xĥs�pg�GB`��y�Pj��ob�Y���\�G5�*Il���Ë�J{MO��J.���ՏY,���'h8U�K+`�����~&�9{����D0��uǈ�8b�جi�s��>Kx0��M�?�>M�Д�����f�MY]�#�%<v5�0��$��E5�r��p�,=��^bܳIq��� �AOw=���S,��0�.':�#m��:��ܰu2v(5�l͛GU�0���Al�ɛ�S�q�5c�pR49�5�E�&/��=@�I��[ߤ�-D�Mh��scX���!F�{�ëGaV�FEyU�<�^Y ������*� � �`Oϱp6z�1�g.������T?�oNhd=S}�=�Z�*��B��:�H]��� �{�
s�Z[�K>���r�ѣ�Ȕ��Ó�$����%��tJO1��k(
*K�'�l
dh&�<�������T9�hF+�GD�N�i�D����CIRd�?�#tĘ�ǭ`���l��T����������[}�L���N)�[V���������L��o�/+j�>(�RY�˟�G�/�7���w�>�_�����~���l)���p���ؕ��'
��_�M�@���4+N�E��	�	z��φ�٫�p�(�uʹ�72;�����]��R����#�|'�(*X*Q=���͆�c�	�8����D畜�,W�2��
m2C�q�ׇ��s�������$Q�C�ɀ.P��G}6-��JI���ݖ���+�9*w��S��&��5X=A�����3W��9�T:�7e�]c�:pq��d�!��kf�a�9�x"--��T?�F��h���4�渑i���1�$M���^���Ӵ�<�rӗ����B�+b�#��m�>߉�>��[.c*�ة�S�4��K�W�B�-�G�?��,�@���yB���0+��)��״�x3�:����T�\�n_�� ���\�H��5�nn��א^�����췳��=<�ݢKJboPt����UN5���nå�v�va�)�0mv��%IS�,D��W�Lo��Q��y���5�@yn+{"�ڔ��sDDHf� �g��7��q��R���������)�y�vR�^��T<zQ�gZ�"�!�1�sUH��!Lϭ���7t]q��9Ĵc����<�I۾�x*[�9~�RS_��&�r��)�^�,���.�v����͌T�ha�����@VDx8�������)ʐ�&�3
`dLɾ���΢�,Z�]�ڒn���x0$,a�;�t̳�+�N=���Y�K��%a:�pq���1���B���C�T\��(�I�l���;����_[@-&	@���s�����;!(:�7�U�P�����3
��9�7ޣ(�"x�lZ�����x~���3�R���N!-mP�Ph�}��K.@,�ݱBp-�l��b�a��ht�i�a/���8u��2��X�'��<ݳk+d������;H�����{�
��lR{&�0R�����q,�1��iiL ���� �����65��ԩ�°=xl�F�N�d��� �h�H&^*��W�*p�� \U�>J�A<����]S��e�>�p��uI���MP�PH��g�&�4�N�>쑯�c��4v݌��N�$琂��u��Z�8�kd8_�#q&�ݑ�o�-��)���=Ψ�o�r�W����h� 2�N:v!�gi���WA�_�v�ښF�ٹ �\jJIs;P�S]o@!�󅗆&*sS����G��|��g��-����H��|4���gD�';%Mι����v�u~q	uG]0��r)��s���s���:-��4�/ͻ�B�-7�S�絥ܢC��홎�ڣG�O�;�?vV�D��Z�mi�I���&�b�P�er��� uy79�h�NZ~�$Hi�"%[
+��*�p�J:@)!��ʞhXp������,�p~O����]L�u�]=�j�6�ngX񏻷)�2�@�?j��\"z�^v�H��V�N�(��7`��8�B@�K���n�#w�
�C[���M��C�w�6��Z�!�*�OL�d����3�U��ҩh`U�/s�R�Z!ԋY@�ư�TbI��z,]�������;H��ri��8S���|b�+�r�0�=�4�Q:�L��Ǜ��e�&!��nk5�\��*vi���3��)e��y�4
H2g/ ��a#��;�㑢�.�+!7F�A�>d��PQ�5����6����ă���_dYt{E���E.�k���T���߬F������J�r5�QJ"�ܚ2���n �)u�r$$���J��"��
:�e\;�4�\a��1�|�:*�8IW;��y��u��| �a*��~0Ѩ���i��Y��]��EBlu�0?|
,);TM���T�΋3x`��ȧ�y뎈�挼���=q�j�:�Q;�COfg���u������v
���w���'ؘ-bb�ƭG�D'�r�0��;���xb6>���X�.��Q$�˚&��:�����a˚�ElQux/@<�����v�+hh�:O��K��ډ���ۤ���,*0����kh=~O2i,aԢ��T{���n�]��������#1�{�dh\@Ԭ_�$A���S{�ǯ���B_�����;L� 9}���c�\g�7j�TX��Qt��%��:�)9xP�.mouvpw^���[�,X���t�	f�ؽ��������y