��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�!��
��%Y l�׾���b������o��ǅ�}|XBi�v���Ĭ���DT�7ׁ��X/����J�(2h�sݤ��E��]u/��Jb;�A�����G��}�n�:9YQlX�,��K��:i��d�����I[��1���DQ�!���p6Щ�§���Mr�<`����=��Ece������"����"���]��h��ɱ3�� ��T��S%.q�_��u�-�F� L� �E�t��)��0��{{����cpA��k��z|j�9�� c_�y��j��}4�F~��U�·H��x�pV��i�߃?Lu�v'W�_nb�.�a�SL�}�����&G>�c�
;������6`Cz�h�,Co��ΐ�7|'�o��ÖF�[;��'�?v����O�_8X4ZTo(MF\L���S$E��� f]�OO�"Z�֓��]Y��ycW$٨k2�+��ܱ|A|$6�頩�f$Ί�!oU���JH��$ɕw��Kܚ?�$4D�r��C�����f�yva���=|�J?���i-�*����i�v�`ͨ�	yA��&���C%R��l�[������n��	Rq_8J
ڮ�Le��?�`��p��5�'�!(`t�&�oZ���;�iR�"������J������{�F"V���t7���x�.�¬�j3a��|K�t0�!��{�k�z�힩�V���{O��E�Qع����i��΃��Kһ���o\�s#��¦R E�-�i����'��P�S��@+c'On� �`y�	V��{/�B|��I�~,��DDK���SSH���Ds����ґ�� ��fv�!Z��?�Ih��_�<�x�ʣ��k�Oj>>c�t�G�*(i�k���Y���+"H���,�m��-�?>O����.]����$��TrE�ĩz�׃��DN�䕵�b���1��%��<5�/��<E�5c�f	WUB�.~j(i�9HDTe�[O�f0~��8ƀ�R�����.Y:M���R�!�B7k��Am{�N�i�_��ВL!�����C�Jsn����u�\	��r�M./N�*��8��޹b������������������g� �����/�~�{����(Z�m��<��y"F����0�!����f"D|+�6Z�w������w*��DȔ�1̮H[��Hq}��,�,�u��ې����.-ّ@xY��|N� ��Jf�'�?5>� <E�V44�E���:��$_=��d�7�|z���f/�} �{��2ɓ��A��ը��	:�牫Ş6^��kd΄|��vB��-�����Q������ն����,@Vo�<�����5X���\��b��-!�f�c��9TO��֡��`)�v��,8�٨�#��J:�>��Nq������H�}m�@��つD�O���O�� �Y��l�� ��g�d���5��I��N��D����5c�dj���n{c5���sr6d �ZB�����0+��ɪEOt��"eo�[7��.�T�Ђ~��셽�OK?�XÇH�R��1VRA�qm��b-�� ���;�]���;Ӡ�L�k�Z����"��S��3%[0�
_%��g�?���H[�5[]$��3�����F���KI-9T�Ļ[�s��`��(o�?C�6}{ Q�T�R�nX�`ZU�8�*���v�^����ߔ�d��|ZD�k(5��7R����}fgna@�vDq�����N~����MF�I�f?.dQ���ߩ0��=��N���qsa^���7��n�����؀�	�5�!I����JΏy2��ͧ����}G���r�������a�a�z�����#��.�IN�!�٣�w�).�����"��t3`ji��g�]|�Y �0��>�l�ّ�:wɅ� �D�W?H�
�M�ڽQ6%�i�V�-��Y	��%����oxEF���)5�QB��S�MK����掆���_�zH}��/�����T;3�;h��Db��}�+�w_{I nx���1Lk�T���	�vn�K<1�5֑�p���0�W�3�Gx�V^'��,�.k;��WBa1�� �ŗI������-'z�ہ�ɇ�s��Ƶ��ȣ�D_�k�+��/��@5�IGM�	$����#*�((k�o��������}:�G��l�%l��B�,`&\\��-�8{�*�@UwRL���FĲ������P�룓U�2��3�<��<�0c��#�D�VF6�=�lO�YFD�_��;�Ob	���L�w>���f�	ݶē�9->���+��xx��p�qp[P.�ZX�/ >M�^I0$m#�{��t���Y�N���B9�Lc�9L��,ا5UvO�$����Z#
��_���}*s��k��P#=~�^���NX��}R��q���!�?Z3���ZQ���d���1��Ԓ�*l.윧���b�3%J�F�� D VD�!h��r*Ɓ�''�<?ɮ|,���(���x[B�,��L��)��	U3D~�^�2�A΢������^��^Xq��a��|�de�AC������<�	���M�a�xD�zH#��`�[�^�)�ء�N�#��?]��i���GD�!�x<�2������ڕ�ߙѰf�L�l:4���f �aD�E�V��)C�F`������GC̤�P$��P�2L{�w�&����t�t��tg.Q,��\p���a�#$��\!�O4�
Yp�/�)qL��5,��{����4�bc������<J�).���Vn��c�m۰�{i��6�Op��P������9�g�7	���s�s������~,Dts(��9�	g+2�PfuzOhr���bsSS	m���ZV�3�h���B>ߚ��k�5��5�5��A�z0�uMO$��^��pTZ����{&uB��?���tyj+�3^�Unѣ	��Ag6oA�X%<=�ʺpu�W��
Q�y/�:E�-�Ŷc���q�q~M�xs{�쁔��+F��ɺKb��͜{�1��Yx3��c�����������6�6*1*�n͟Co=��t��.N�.qs[�kf�����۸��a}��֥»��_ĸ8�60����y��s{��}5]�A�?H�)���c��Vۅ��Uz�
)d#uǐ��ς��n�vp[�廽�oǼQ9\dQ�t箂.�^�����hB�A+]<��>����}"_�DPV`����� ���#L(��uw�Վ����u˵�I�>�x��B��l����%|ď��]�V��F���w<Qp���,�,f�K��2ТI��R�/� ���M�O@"�/�m���Y�Vu�\�:@�Jtŭ!�w�ߞ��|�`'Ų��+�nVPԡ�1w�I1ԲoF���i���/!�/�L׸���BF^���CY.�._��	�cl]�L$p���Ԥ����( �%|��r���iX"�z��_��P���A9lk+|��#�$2�¯�?�%�S�=��k��ՙ��)���Ն��4��ٜ��6gy�Y�j��-[R�&��V�p��&͇6-5�_��k(ʭ|g����h�G�C�e$3�;�G�8Ro��H�y+	�~��q��[ك��,�Xf�*J]J�R�oo����Y�Z�K���u�����2G����j����k�[���KRb��g��)�d�E�M�AA�٩�I�_�m�hY��[h����qn��0#6���'����������}�I��Q�Z�0ݕ �ӓ�c����8�`W�n% ��u;������(n��'�K�`�4��Za̱Q"�$�A�x�4-����Y����-.���g�K�����}�Kb$H�t����J#g��Z�R|��u9J_�4�a�)[��[T��ZF�s�����B�{ �P!H�ܝa���w=�@Sxr1yG�k(d
�޿ԍ����S��n-����軃��kT�O�U�8[��'&Y���*�)�ު&x�c� 4%
(��E�<�I��J�%��
~����x>�D�)5C�(Ğ�ý���D\`����%1q���fn_���m6��� ���%Ae4b��&{�wfxǁ�Nj�fJ5gO	�&	id�ԏ+UwJPG��!��S;Đ�7��u�;	s�n��	wM7g��(�n0G�^���$�H%�u��A	ؙ��m纃��)&B<%��Ieo�s��2,9OQ�����]x�}p� *��hÙu�	��1#�:���cɐHwr,v5H�8|��Nݖ���,�[&<x�R�nk�y�T�$�'��8c��k}}j#����������B��'m��Z�u�	G�������f���g��z�T����hQ@��l�٤���mYkb<�/
N�����X+�^?*�56#B�g�������{eNmIß�
lD+2�1��-�:� �p�^�v��m.�z�c�G��SacN5�^�5.�>���o��'$p��U��"��G��?[{7�Ȏւu2*��9(�N��;т*&8���nqHܱ���hS��t��L��ur9��H]�f��R�L~=�-~~0T��:T�����{�zR�r+�9qA�B��"O�ԉ�=bMt዆�+�y�,��&���5��_ȅO@TT�Ǥu�E�8H�+��<]���W�*L�)�qPB�l��y�k6����t�\Q��#6.��Ӛc�E�	���6��2�B��NS��2��֩����$54�L�z�tT%�d�CDj*3����oDs`��~f�� �+��'�:4^4�Qზf�z*�4���'�K�du�k5~���Q��Z8����֠��X����D	(��K�������H�́b�'�)�<}\L�v�W�؇b���c��/h"0x��T��[5t�7Yp��wQԫG��@�~R��b�G�������kj�+���]˛�7�IK��f��!�ǭ�2h�u��{0�sߕnǡ���oR�)�dt9�+-������/�1W#c}���Xǹ�V:X]7\���MΡ"qd>)��n(B������s�TO[��Ӏ])���y=c��3�V���~9E���O�!hmLt�[}������Bv<D��n�,&GxQ�ٟ'6�Y7��qstb�/Ip�9����ş������k,��a�m��H�>[Y���n�%3l�U�(͍;��V2�k����K�ˍ
���5.��ǐ�2E~�>I�1���c��	B� 2�o'��2�i��g\�� �ǂ�����Q��P��-Q8w~ab
)��yLa��Z�,AEJ�OE��{���k[��S$������D�?Hݽf��|5������&1N�a�9&$@U��=Y����+wӃ��D!����E�k���&��f;���@/1��<2�/�(�&.��_>gy��ڝ�M
.��(����0��/�P�ܘ���q� mfc��ㄪ��'�9l��T��~���2r�A"�՘��;A$+�ٶr�_��k��b�}ŋ���i�y�(���X
������꟢l���Tܣ���~��W�����Apa��ݒ�YcVRZc��nf6���|A�����N@�Y2X��hdV<�s?)�93DLb��Y��oN<�k�s��Z4.�48Q@1*�Jg>�����g���g (r��0�F�^!RX�V�a�s�3�,쟠a`���m=},)���Y空�_���*�g�ݶ	O��YY�="�vO"p'C�0;���( ��)���.��"��ֲ��2���oJ�
9���������o�*Wepp)��eL]��8�:�(�^�*���>�W;+$r��-�[�Ƒy��]>B��L.4�xÖ��ll��</�3 �F<!���]��j�\�ك�g��t�-��>��h��c�^��N�9�m��	':��j3Eb�߿��u�{�`�N�ѝ���̞�5�y"�KJ Y��S�Ƀ����i�IH�ôS@�EӐ�$��ɷ��6GZ��MC-�1E�m<v���A(��$O��jG��&�5jt�B����&��0̀h�W-p�Q�L9�A42+�<�
� /[e��D\�s����(�B�Z�/*��)�}l�_Ւ8M4l�6����=�6�s_p�vf|g������9l��Q�w��L:~����&�y6��|��˙��T�Nf�Q���
jnSG��ۧ&��O{q�1��!n�ҼR/���|T[n�LU,�X�u���-���v��I��⭎)����c�]I���_Å�qB���]�9R,��)����*8�nf@{���d������|axz}���@m�����/���\��Nf�i��<^�|�Uƣ� Xrd���š���@��j���F�^��c�O��[����ƾ�s�n�s�pK$�9�O=5
v9�a�.��
�d�n�-3]�&���x�B[<iD�m��{�F�ۥ�EV��ZG�Lpߤ@�p�;�M����>���:1G	��e���U͕4|�6��L�aG]Y^�����]�ܐ�h`�NkdB?j5�<���%$>��9��̗�t��T�?6H�,K򁙳ih�-9��<�rmK&��q�X���[4��qO�2YӃk�{I}�-��5�>U�b��e�Q.��j�����6>1/������������4���4׉��h�����=!�q�VGK���_��#h�ُ�O����7RYߓ�.JC�a=F2�s�e}c� ]����ȯ9H�L��u���"�w��Ց�ʒ�m	0�-4(Q��m`�]��@"�/e��( o��ꊿ���b()�t?�7�t��Ix��LG?�a��ݡ�U�L�8�����h	��%��P���J��U�n�N�Dh[��Ω�$��#�$]��z���;o���zl[��!�H��ZP��(�Yfo�rL�3�اw�#��P1�O����У�9��Z��5��m�=�<t�pr3��o���p��A��A��Q���	��+�+�c�?�����ٗ8M�/�;�+���4_K���)����$��3Um�Jت�I��_o����? �A!\��"���g�$�pv�H��L�@Z"f�7.U�埆��zGt�,�N�s1�X£�^���Ċ](~)�� �dڕ��``D��ϓ���� =	���,����
YW�W.
���+��b0�=�i7�,d.����L+Zq�J���0܋t��(� ��Z�5��z+V��U�Q�����`D���`X>Z�m�T�G*eQ��Y��m�p�ҁ���#\��RO�j�[v���$��d� B"t�A��~��is�3#[l��A�N�@���+��f}Y��`;�{P�aW`�Z�$�3��Қ��V���|�=��G�h� �əN>��<�� �{d/j{QL��mc�H�^ ]����z?�)uw�5�Xf�،�^�@�6���;�oZ���|����������H�GxWޏ��x5���$6S~��$����a�$�$���M���73c�	���<ė7���
sI��#���e���4J)m��ғ�r�H1k\Ʌ�L�^s�D�Ѡʧ���0<���W��<+Gg�mA�=n�2^���Q�@�>���`�\��^pQ����Қ�d;l��5oz�H���\2����,6o�$��I#v{N D}�`��l�F4g#@զ��.I㟧��6��Dlhѷ_+D�Q�!+����eM��뤚��d:��'yT�U�|1NƷ%J0Z-,���P����=u�����i����W��Um���[�SR�����)����qU��2�ގ�VW}��`�3�����,s%6v{�֔ϐ��-�U�~��YoF&}G'DJ���Y����g�j��3N�����!�DhM�}���%�.��x�g#e��Ӌ��:;y8�3�8����E>�w]�&�z�?��߲��F
P�[���)J%%�j_�-2w�����A,���<n�4>\�F������$B����L����4%�$�Q.��ye��/����P�^�1�O_>x񥮆�"��^Շ��J��>�Kn4Y7D՗��Q=�Ÿ'fݬ.�V),e���,G�	�5�.�"��
�7H�t�3O���U�v5IѬ],�-\P��6���)������'C�;�06lySa[�H��B�:���{� ����v�,h��%3x� ��ƣ����XC�ڄ�4����B��i�1��0��:���m9��?�-Ķ����:�{�DTb���1��I ,�qq��j�`��
m�!77�ݡ������I܋�1+��Y���)�haZ����_|EZ�X$-�ⰷb;-EB�������>ϵW��/	j>#����]P��o�r���p��@��	l��Z���nH��d�,�鍟�Xb�ld��a,�$�v>e��]�:mg���8�v���y}�o 	i�o�ҕ?�d��$�D`��~�;�h��kg`�毌:����V
`�Zn�IC��[?th)b�e�d��*��^=��@�R�Ѡ�(��\S�B\(mPA�Rk��E;Z����Wl�	��a�ح��O���'s��X~�ˣF��Y�� +��������}���U�h6��K��φ	��\aF𪿋��Y,��^0=n�S�w�9<��zc����+A~�~c�`�W���Rh?~n�nU}Ð�喼V�}�C	�Ƕ��/�dh�W����P��4��D8��P�d�2���b���$������p4�,m���l��[��K�]P�V���Œ����2���0���:�����p[m	T�$�1�1��e�m!{A�o�7�2�}���L�@J���m �F�8��B����q��wy���O�nptb&��!������u�!���"���\_'�º$�]L
!�2d5A�'���B]Ũ��+>]p D�GF�2�A�6�Q6o��Iv�1��^�2"��1���2�#��j�̇�&�7��<�q`��H���Et���Nn�)N�6y�3�3o#v/�y\i���8Q�S
q1���Fo���)T]|>!�C0^�(q��Ri�C-����?H<-P�<���^�dvA��	�(9XOe��c�nS���t�_�ք�<��%���6��Ô��.�$%Dg�>���>�:H�� �>E�Q�tm��rx"��/�yY���w�r�GR׃b ��\�7NG7�N���3�MJ9�\h�۪n��A4!��m�H�˽�o�~A�Lg�mu| �(����ځ�t�5 ��6�C�r�p� ���S��鈈N�@�])��~�(��S�m8y�E�i.�����&jϬ1
��x�{9�Nn\`S�^'J&����s��x�@7���B�|s�I���N�``����H}y�2���~fs�Qn�F�b�����/
Z��qlˊ+@F�m��쎂p�`���U)����`����m��������g��o�I��"����6�a�Ԡ�M��1S��<�Ȗ��d�����s����� :v���~Z�G�Y�����T�����E����,ȹ�3�̟��)1rx#9!bi[l�]�>�>Z%���oN�s��:����UV���(�[D ����׌�1�8���2h�6�b�\UY2����tZ�5\��kX���%���:�ؕ�}P��/���/}J7��ۘ����{��݌�~��4�8\�	�=� �5��eȈ�[��������&��m���hX��mbH�-މn��'l�;�Js]�$�~��c��F�K����m�\C��ɝ�`��' $�Y<w_Y��A�D�4�!f��-Li"(�$��O�R�mldU��4�L�����<�=��/g�3V�o�w��5�z��
;�4�%T���i��F\â��q��6�]oiU�9����չ������@
uq�Fq�B+n���L���m���v���F��H��<vD�X%��#�2]E�Xi Ϗd�j�e}t�W�i�;¼��[�E�N�E��l�um2;�����ɵ��(�`~b�o�4om8|Z�9D�C�Q�cc���QZ#^}�[�ܦA��*��v*Gq�L�����@$Ɏ�p�!��)�,�xFhfZ"6���V�L)p��e6�����
$��|�'9�yI�����>�)��a���v��6����B�x�!`�A#�����0:\�������q�6����)��%�ݑ�� �}���W�-^%,Tæ}l�"-}�A�x��4�ͩ�M�#��1h����_�Fa�8mL�tf�X�T��<#5�3����s��9D+|��V�Y�~�`V�0��i�p�<�~�oh�)z������Nĕ���ՠ��
PY�H1�.gp�"P����3��?]����S�3OX�a[��\�z(�N�V��j*f���|Ř��"��^�w&{�<�	�O��:;r��i�H5�#�7��� �<�-u=7��fI�j�n+e�-y��6�;e��ޞ+�t�����m��^�V��ϧ���{�ii_����^��Qҩ�4$�@�{œ:q�3� N&��]�=\A���>�.XME:�^U	m��FRa!'�K�"*=��T�a��K���#��kl�K?�Z��31�Y,���q��>�u$��8��=�QPr3m;&,�D)�k(Ͼ. H�P��t�F��؏��X6�
\8����Z���e���v�U\�P�oe*��򓘄*�ϋ�t�,R�A��QB����iV2�N$Q��wp�p�[�C %*�/>��˺}fki`>4�r��¹�ϼQ���9�[���1�b�\>[P$�6��ro [����7f��`,%���Hcm��Pe���sG�����_mc7j��a�N��i�n�� G<ᣧ�����J��Zd#�XVSޢ�a�� �ۖ�����A���埻Q�[�xHsgJ�|)�ى5(8���)�t}#�}�^��;g@��Q\��2J�(�C*g�ͳ��r.j��pǪd�uZgM<àyZ��t�m�2?ayr&Wma�@��X<z���0S�D�Q��#�框�2)��Ҧ(c���bU����n(u��t|UO>���$�� �R��Z��l?S�Fi�{d&-Q�U-�����bh&�ؒ@c��'�|�=�y�i?χ�_˛w�_j'���z*:�$-�0s����Df��w����F���&Y���#��gjX��)��8Հ1X?
�;��p4LcJ̬ē�yt��$h0���Ea_�D�dLcc�%�&8�b��O��:ֿ �����s�wa�&7�S��Z�Y#���>?*��X�RqI���'�=iT]`�g{����{eE���V3�-Y[�7{��� �K��X�@#��˼�d����<$�xZ%(��@��@�����O{ZEj;#��څ]�^�T����+����2�`��{E�D�zD�Z�B�T�H�<��/�����ª��_0��H^�jW�}�8�����_��?F�ZxY�����.�ю?"�	���s�E�&5j�[�'����smi��UR��3�CS��k>��i�o�2�3a�w`3�o&�
���r菼2���q�KA�G�"i-�5)s"s�;r4�	6�N�?q�����Hoj;Ϊ�q�JA���5�l����
0Nջ��� ���P�����
�p��9;!�7m�Ս��y��n����vؚd=c���o�b`}��#J��5G��16��S\m��3���OG�3΃�����A�VzV�r�eC��Q�3�e?(�EҎ�v�3�i����`�a�Pã�O���C'�%������&a񙛬����sS+ �f�Į�;�t����u�TY]~��C�D��7�8��zX�P��$W�R~����-��g�zh���9���y��7��'jE�V�+6����	u#��ߝ�Ǚw���Dx��;���ZZ�w�;��^rg4�X�[��_��I��B�/�,1հ�G�`�q,h%@v �.�U~��ͷ�&�@3M(�Ot���߯�d�PM��ڌ�����t����#!Zl@�N�>͑x����8oX�[t��$q]�&'��� �Ї�����.0-Ηh����E��NG4 +�$g`ڕ��������Gz�ke�dc�P~�$E�������P25�e�_e��f��ڏ6�@qg��&���if�Q%h����-����0�kl�{p�6.�t~��^��ף(=������`pj5b*���hC�ա_�hu.�a�tQ� �ǨA�HM�t�:�*AT�mbҁ�n�U&�;Y��Wd,35��@���JհAO�r5�t�	9�L�
(��5msP�`���~4��ď�-G��{���V�_��ڶq����&H���Iʯ���٠��a�����*���N������#��H����K� �'�0Mz�.v��U��9K�P�3r�}����+� -��M��I���.��98���C���s��%;��xU��HI}3�q�o�v/����>�5^���`��NI�:H����k�]-P�&17�S�ë� �m��%�PR��<)nK�'L�ssۗ��ux��Z���p��#�t0�nZ�5&
o�x�,����q1��+��sU{��g-Y�i�!-f��_�1E��%�4���Lg��������#��qg0I
PeU �V���*���"�H|���)��b�f���)/����Ҭ鎋�s�f��	���)���¦[v����qW��J�W�z#&�L���^2��,�"�C�u>�m3��|��^g|��.a'�ia��0��k{��Eg�I������ge+�K�����m� ��V�����9d1y��tܥg6��OTx�a��@��aX���94�(L*���N�Hrٺ�k4g�΄:�ǵ8#؇l�����T�{F6�zwX/CR'�e���;�~V^L~:M��)�E�'TsI�/��+��#���=���;�ʙ�Y$�7D��P��.t �)(d��������<�3����6�'攅� �k�"�X��@,��ro��n�X�������A께��ӏJ^R�e�nyK��q�zr��o�F��;�#	�#�.�ڻM��s��%`<~��I[����8z���Ԋ*H�o>�;���g��#g�H�z2%��[SR���@Շ3�48��{ n�]��9�;l,m���&���%�Fy{\���u�=��B̆-��+xA�B�S�y�W`�R?��c�rF��#�7{I�y�ݿk�Qt������R˸��|m�D���K�i>H1`���E�&�9�v�;�р�h�؇is��i����ZZ�ȿ�X��&�"��̳}���!��?rM+c6t���g�q��☍� �G�sk�A�N� 3��K�$j�#C$D���{EáK\*x �@Z�V��%�./��D�'���H����q������>,�����J�S�8�P���W7�y.D�F� P�����89ڡ�$�k�~��L�˖��y��l�:�Sf�ѷ�V�Nk�ɳ�Op�8Tփ����D��E_G/z�բ�����}�+_��eS;���	�9�áD���I���n�X���ya69�)�[��F�D�s�z�6�*�Ȼ��z�+�!��0�1u`�MB� 1���S�b�N�U����:�- ���X� ��X�Ǳ]~��ό�~�A�����{f�S����Ŭ!^1�n��k���K|�8��W}�\)�k�M5����M