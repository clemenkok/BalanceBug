��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�!��
��%Y l�׾���g-�hjxZ�bs�f��H��"7�߫�,�y�z�%C���<	� �u� *h"9��/=N��S%�v�zew�����`Kgޑ��wA�4cYI%u(l�d�������i��l͇p3��26.��x�`(b�o�ٌ��!{, �`����
e+V&i�pǌW���������F�4(=�	��"�Wy1GŜ�9��'gS���-�铥�٭�i!{OL�q�.H��COݵ���� �M��?Jfy��v�v����kό�.9i�X����I�j�7�!GR��-�a`"S�G�:���u�2{��:�Gl���^>��j߳1��W������.�j��7����u"�F�%+����������囔O6�!6�S����G�0v�q�D'۽�?��{/,����I���f�Bbl���.�h\���no-���5�z6b݊�2�N���5%�jˆi�1��|M'�J�[���@cY���'99�<U�1�+0��{�uB��Āg�v��9�u~�z�l����*�MV�f�$��i��ֹ2��i��Oa]�gte51��eA�[�|�߹������7@a~�<��,O�a�|bu�����̈7p����G߱i�k��鷃M�5�hb�Y������y(; /���<��ޙ�E��*����T��_��T�ݖ��\�� ��K��=8��.�k�Uˋ��u�1:g�s�7DG(�t+K{[j`w���
2	�]�1I1$v�6��ǧ���B���d��	��s
���qaOr�~ڻF[h�����<]��-���E{��b��Lp��jG��rP��jݷ��L�s�����Y'o-XF``�+���vk��*bjZ
���4�׬�zmt�)cMn���H�����C���QR�fZM��F��J����W�PB�O�	hb
ґ�;�6��XzbW겧����.��1���A9OMg� �s��gos�ڄ���ra]*��ݬ��Wh�=4_��S��#>�&�u����Q��/�6�Y�h<�-��4�LY�FW%���O�)����:��6t�p�.T6c��/�wYd��;&��h$�JP����fB	�7���\��7��
��J�����5�΢�:�Θ�@x|vۜ��H��B��_�=�g8��do!����ބ�C���]�/F��@�"ӻoO�P����%`5&ݽ�ɈU��j���E*�_2r �ܖ��i�?�W��Oǎx�=X���Smu�{��+�ь������(���M��
M�H'�#�"�ߦy������o��8Z�����3�"�����:{�<ލ�j޿>��N��$2`�q$ߞ�ְ���Ӥ�x���ܙ#���W{��-�KF��9�H6�ڑ$nZ6 l@����[���X��W;�^��&"ը5�0(�.�G$�ӕ��]���i�*�<7��+l�w<v��-��Hr O�����E���]fa�cV@��"L���+N�_�0�ME��>lZb�3�3Q�]�/�;IU�%���a�
����: <�x���1\���<�8Dk�������NN���lN3���"wo��h��x���/��0܎#���o��rg���o���n_0���gb�(i�g�y��Q�����1�F�~XL�p��z�KoII���?�1�' ����JX�^�\�?}ė2챥Y�?�~�,ܬ���(Ύ�W��Y�d���؅���&�?��ަf�z��"�⢶3�0�Ps|w�5��(�U�O��`�Q�ORW���N_�|bPe-��?�Vm0�w��I�ނϿ�ː�)u*9>���WY ���/!>����R�r��x&z&>�Vh�s������j�k1�}.�?���Δ��xD5�/��!WDDK��|37_+a�M>�"�����e� ?ڹ?�?7��4X�T���=}����43���`:�?���U]g��MU9����2y,������p�r.�_F��r�k<l2�m��vZE�]<���9}�fY��|9�q���C��v� �V��xȿ�I�
g�d��u�;�{Ơ�${7�$F�t��#N�Gm/������@$��/4�DYd.�(
��������قy�ڏ�t�U,s�/�����6���b�U\f��zU�g@��W��1W$C�}N`������φ�Ɏ��V�t��V�tt������ˇ�ؠ�^;g��"��@H͡��u����{Ǔ����po��&*ͩ�u����U�_+�NN�U�y�+�&+�sM����Xqq]&N|�{ֆ_�|0��<���F_0��d�{Ն�XR�wC�\!"��t�`�K�Tm5ba���]va�`$�2�a�o�2a�Q)�;GQ�x
8�Z'd��y�l�B(�ِ�T�����WQѭ'�uG�GSD�g�~"��/â�~�Y��t����h�b�4�ٶ����)/�9���pa����9���4�,̲e�q�S4�1 %���0�;u�O��5=�PD�RG�]*�����F���_8$i�Ӗ	~�&ICe%���F���1V�:��l7SBF�����	�#Q�[�p��Y�6��F���L�H�� d��`y9R���<��?Qd=�[�*L���ˁ$=�0����'��K*k�UY���1��&���<�z��o�7�J9�	ʄ�z���Qh��LgK8x�Aw����;������NW7��SҶ��c��GC'���^��mL�����r���t�N��<���7YШ �c� �I��yҮ4�l@�z���(|�c%ora'4 @(�zPw1b��/"9Ne�;��>�>�BsA��6���A�5��B�����4UÐO��}0=nIn�C�>B��0g��L	�l�m�uQ<Ǖ���sc�A��"O�+P_�_;(�i��t�캲������(鮓��V:W�[b)�|/��`XZ������ˊ�q�(�%>�D�QN����Ж"%f��#�r��~�K�dRe��n;�2��kP���<��XY�����d���؟捛�����8��;�u����k.�Ům��2	P�f}�ψ~�x3*NE��bav�j�16T�..�r]bʞ�'�ԝa=r����J� �l��e�*���Ƹ�I�tx�|�E��%4���{�T��SN'��B�V2�\f�l��n��Y,B�.�ZWV�Y,��젳�n���=�Y� �θ�*~�2���kPO��!z��<(�v��t�cŢd���ى�,Y���E�� ������4��F"��x�(.�z�N{
��P%�v�C2El�Ñ��a�i��9�k�~�FC~�g@�	��
Ӄ�6�MヰǇ��(Vm�ߕ�o  ������燹����Ck�E��߆����j�h�'�m�;�� L
y���A� *f��G�.�g�\)aa�yS�WB�7|kj�8��HXT���mBĨ����2+���酱�G7�A6nQ��S�Q�ۏM!�07�Y���ج~A������S�@��@[��vw~�6D����[�f�U�B]�}��#@
�Mӗc�����`�?��d4���eE��&u-�tW���i�۟��vGiR�M�]8U
 �������q�
�����.�@� �پ¼�(| �q���=���۸q��d�0M�"��QIH��¦k�*W�_Nk4Gz��L���֢Vq!�*/����;�K7F�@����v��la��m|O���,؉�����?��yC~�v��z��g�$( ia5����֍�7�£����`~���sr!��+�DK@;��Ԉ�A9^���H���ǐ7`��z��K$�;ІӍGY^�����8�S�1Fh+��wڂ�SR���$k��b��Hz�cH3�Pp">	�sxK�Ki�q��4��(�Q.�wp���X~9��<2����$".� �؜�҂�\B��/�t?d���|�|���2�6ݣ&[��n�![���4��t�0Hgb�����*������/��)���3��%ʒ����orY'�CT"�;$�M*�'p6Ic��H |� ���Q޷�F����*z�_UQ�Ef◫\��j�<l�*Nk�wW��;CF !���Z�� |�W��CB�'��#?��u�A@��A� �j���O����b};)�paZ;#�
.}q5�H�%� '��3��8lbD��(�V ��J-Ӗྸ:=MF۰�?�JV��LC�+rG�ip����:�]���U���Yc[� ��3�7Y"9ł�Ż�^Չ�X����j}����a#�`k�F��'��݃�[�۞�>"�����88]\���ŝZ[ �|#�6d���c�RR;��P�E��hS7�Rn����ʫ(�
���c���ܲW���HY\2 o#�zߏx�|��/��άo��Ϸ=���O%�,�A�IZ����H���8Q׌?��.�C�w�5,��7V5l��G�ߗ��;���@͗Y:�\�
e�1�:y���y�+�.s_�#��֗���[�kS��;�yCS��y�U����iSt�Q�@�>�~c��~�F]k�MQG�J� ����g[_>S�׆Q���|�QKHMW�b�"0������q�f����dST�\���ٚ&#���7���6����M�6L��9�� �J@�s�N#`:����6�x����UXc�%�S��ziX~⠋΀���v'.���dO�tG�!G������l��H9́�ǚϸ�2��-�L�\3��['�g�\?��ŵ�������i�/
r�s��Ӷ��P�ƒ�A���!g�
���Ӿ_Ob���H�� �D^].�~�m��8�_hd����k1�]
���D%��/�K觩�����M�B"�hCK�%�	E�+a�dSn����鼁�![��U9�s��Y��f�����������2���o6-������CQ��3�\b�����s*f��	��%����rF׌��@�Q�	|�*�t�+3���g%|8��� �����	� D�f���K���+E`��V���?���wѝ���T<�6�2�أ��М�?�Z���W�Lg��ҡ�lA����8e�g��b�<M�Vw(5�n<���7��1��TJ��֭�`� iQ�>Sd�W�>��֍�iؓ�=&}�P&=,��v	�g)�pC��d��gu�]���$��FY�����I���~s_� ��A>7�,���_[wFp.՝��kk�Jh��,2�^�6��#���t��_9d5��bDɴ������*���5���_)xm_.'n�e�ۇOͭ�}�:�G�r��h��{�V���o�����F�@��K�ήYf� �����SKq;��p-oIh��P�h��Z���4��U$�TNd����:t_�� �]Z�ͺKe���
�=5��J�Ȏ�T�y'�)5o�:\l_��	?��	� �SVXPs"�~Sp���蒷�Tto�%C.��w�m��2�I�^�1CV���#���^ibW*Z��t��!�,YX�mh���l
NXE�tLi��v'�.%���>C�����9H����>1۳����E���JaI_T��f`(�"�'ԩ���@�ǄC��g�T���D:j�[^i�m%����*�;�XU��OvG�Z�_')`�	�^�,�-�KG̈��do�j�V������-`���:�9e��`�(��y�O6�i�lLD>ҽ��ab�񉡻 �����-��gq�-���C�~^q��g��&*�q�&[��̥��ģ�zߣL��}U}��Ǡ�qu9ݻ1uv��SCJ^��:*����y��	�x0��eϼ�P`����O�P����>�P7D��Z7���:�4Gʞ�5h��qi�L��r �Nj@�3����Gq&�b;(��naΔ��O�^�	� �)Y�HJ/! �u��w�=���Q|���,��͟W�~��n:1]��Z�a�;��l}��jP�ƪ�uxu�9���Of-B���ť�n���?�� %��m�cm�$S������)C�5CMq�r�K�˓x\���t�M��Ю�p�U�w��k�R6�<��(���k����M}m��*���dZ�U�EU�N��7&Y�z㟦.��؟0���{�txhݳ�=�S��6��u�PP:�l�ufl�4_؏�[h�J���%p��?�_ �1�g���lԵ)�~g�=�H�"���l8l�6E�����AͲ�N�j����[WpYя��빊�$�S�s��fZ,��:�!7Pǻ�a�f��^��㼕�k,�<X��-�d���-�'^
�=�E/�	۰١:���д��6}]�l���Y��:1�q�*��S~�QwGy>`��]>�я�6"�ܢ P�x��j7i��C�F?	�w�cҘ�9{i����3;h�!p�;��Nz$]U��K_(�}�L�)�(9�;�.g��[�9�z(!Co*��b�3��?��'q�F3�\�躣'��z�y/U��v8��6mt�uА�21uT��օ/QN�����?\a{3��,�^��p�u��)��~@'�dgyVVuO�������)!J$qj|�G-���}��<��W�)%���^	h��75٥��&�Z%a��[��-ξ�=X.
/���"C�lEW�R��pԛ��0T�0�]��������!�p��qܫ�J)GE����Cu�۵�-����\�g�ڦņo��`�(1���$T�a�w���/`��h˕����\��uf�ΚrH@Od{����,4��d�	)L��q�L���t��x2����R|�'�F����p�����;����s[��C���2��7N�l=Z���!MW[����H")\W�_uJ��!xJSU��lM�o�dKF�®C0��:9-�>P�\݃��$ڈ�Q3��w_>�Ś�]t,d���<B�ζ>/$T,Ǣ�ӀC���|\ �ד�?t��V��VR������A�oi�P����ߢ�ȩ!�K���&AZ���/���F��T�|�`�A-�C�;����@3�~eO��6nf�}1����I^���)��%�	̓`)l�?��T��.ܔ��U�����LQ�O5�4�9��8k�<)�1��l:��,�V�!3�"��ga�����b�<�Bby_?�zW$����	bA[�r�:^l)&wf���3�_�$���UVw�)�#J�/cc�Ru�5�B�dX߄�O����K�c*G{�9<�:��_>��~��ɞ�����E?�d(��f���*"�Ӹ�)��z;v�<q�2�2� �u�#�w_(�ӡ��@��F���)�Pщ\u���pF���I�0��>fT� \�:��b���ī����'�t���"�%���.]�Nq���7�qE�ũ�9�^s1Q��=�	��f?m�K�h\l:�����m,.��$:LjB���u�vI!g���?�����Xu�j ;?%4�g#�r�O�&�#��C]o�v�>��P�	�m����3/�Ĭ	K��a�9�HV��f����f�|� ۙ��9��Ѻ��L�ʹJ�cfY�2�M���'}}m��	@}|	��G��Ǘ��M�?s�@���/��z-8�����W���2u�앆�B���¡|:}Qf�[,�S!��=R{b��}�G�|�h���b����~â�Lsr��!W޿�;j�m�'�	���J��}�Vx����X踣`E�ā�4r���P�E���21��o�mL��ni`�-Ԇ޸"�#��>}+pX��q��Q˗����؎��#�9�5�tl{�r�Go�v���G&���&��qӮB����\.�:�ھ���)�]<\�Ή�{��RRj�g��H��F��-RG�;��R��k�n���[`a_��q��p�@i	�ҹ^��#�5P�
`G��V��BC�I�AH��Uػ�~�5J��<����t��g��b���<+�x�6$~)6;e����k�0�������!���18�?�u1�ĩ`̾��*#�>�Nj��@ŋ��"t[��6o*nQN�UM���.�*�_�K�bwf�����J�����t���~�(����&��ab3d��q��Fd��e��j)�3L�72�~Ԓuǒ?{����o*]a�X�	���:������#1ba��K�*��js�b�wb�:c�tX~���'�C:�U3X8���Rb���Hw���]ZGG��8�d�H^pg�ӥԹ&�O�c���⣮���� ��v��
�6�2w�/ˋ|S>Db�fl�o��'�ٓoM�#LnRz�!�#��(��:uY(���>l+wW��}��d�Uſ��n�g��=����D��{���n�W&b�R0�v%<_;$���]7>|�+T�d��[X��V����(����^�]v+����i��*�����K�xe���:���yw	��~�<}���^f��A��}M��ϛ�E.X∔`l&=\�gݯ
�N�<>K͑e�� 5��ZN(�VD)K̢A�T~ǂ��N��cq�n���fJ~�T����}ז����=$H0pׂ:kE,�1
��UZ�zܒ2�;c�V�w�]0�<Q���tGL��\���Rԁ��t��Tk���48�i2Q�0q�{����X,ޭo.n�A��RMW�0��_v�C���2��ߏ�n��+��'�j�~���E���Q��B��}���Sq*�Y���+׏sQ�X*�b�И�x���w��C�.=�no���꾼G0��;� �p���M�:1��+�o��O��a�	�/���O�1��"c��_�-3C}M�U���s��&^@+�A�u#�D\Y3=<��1����Zjif��{���5�P�v��*S��A��~�a�r��{?��|�u���y��X"\Q6j�P�~T����^=�ʐ#������Z��h�.���6y�m2`?�]�$�Me��l `*�9����� d�E��3�`���	�Ai����;�.`"PS�ç ����4w,�x�̦Q� JTT��'˟�I�}w�ќ(�J���S�HZ�˚��Rl�Xha#|܏>�{�f��j��u�<�Hth|Az ;V���A��䚳�"�k��\��&�t%Ծ���4u�ʸ�L8D�󾕗���.�!��T��w�7B	nUJTT�@M�,�j�����E+����ן�v�ޟ0a�*�^����!�XGT2Wa��J~���K�'(����lo7���ׂQ�0�	1X�pQ�뗑P�?h}"��}Q�Ad��'jYϸT��@��qf_-��s���r�2��Ff��|MRQ��7��6M�)����Y�Ym4ӧ��sU*l^^�	�HPšV.����N��6,�v�Ĳ ��r~&�9�2�2��,q�"�m�0�� ��w�A3�a��{H]��ٷ��>�!ڽ����K�.e�!z����G��a��2��4�>Ĝe8�����Hd�H��/;���8�a��Gy1��h��H�x��y�[��l�ݬ�ChG��\n�H��WM+��ɓ��GF6��ބ�$��Ns�!%�����n��A��bQ'v�1�K8�a�.���zpۤMh���'�c�t\=�
>�L���M�5ӸAO��D2E��1�b5�M�r��`��&������b�D�p��˙��K��v;Uڅ$B,Ǫ�V���D{fc۬ať ��c�Go��֥�4���+��_�}hdQeH�,����!>����T���/���`��������Q�g
�c�l;�����퉷v�of���ǿ��g���7�݃c��&�wa?�a��r;�Tyf�B�*�����g[�/1ޚ�3���'R��{�KY.gҿ���o%��_�5��7��lSOfѡ.�٪c�:�D4�AD!�>��R���*k��B��q��o���L��x��`�w�|�P��j��
��5��� �sD�~�T��H/�G��g��N0K�7�U�a:�{�`�5N|�y���������8{d?����//M��Z�#��aH-bɛ|�x�:D��m`�Pg�7��09@�<^d��B�^�m��B�?��Ƒ�`G��b��+�)�'\��KL9Sm�� �(�
��5 �+�%��e��:��C����2z�� ���y�rP�B�2�� B
<��z����E6��H���)���,��y7���f[�ɖ�-��_Ʃ�̢#�r�ɛ�Ķ4��ﴱ�����w�t�́,�V�����=�;��*�R�ԕn7�?Q�7���:��o}�p�|j�#� ��-Y��3�z�+I֠�!�t��u�o3��c٫2��7�wq��jSrT�k�N�3M���?q����).�|
 ��X]������YN�}(x�mgxX"q���3��k���i�KA>3�/�ό���"bw]�~:T8����hw��A*��������\��#���Sh[8ӫ�o^����o�'�P��GǼe:&~�m\��R�'�j�������y���*WЎ]L��U��?70n=U�0�
O�����?�;�ք�{���!4�ȴ\P�%/b��wŘP-e�j�8(�ކO���7�4��������9[��"�?u�C��D$�\lr�
��$�U�@�n��K�	E̺�m�:����"y�T���c�G-ȓ�0�B0W��|ͅ��<������N���&VO�:�������v�(�L���yJ��5��,!؉[x�0�2[A�)�yTk��|�xex,g��К|{��|E�m�rm��Z�L�	���m��t���v�pC��M�I>_���Jx_z������c+(�?$9�)�\�}�݌�i���|9�����Qom���E�[c믑�b�.����{���^�HA�ؐ)�/sza7��,|����2���s�� �eT��&�94�e��u� �<�:��ˍ6x�al��?tP��R�/&�Js�7��R$C�SpԜ�V״���(�V�0Ko%X������I'�eǎ�v\to�>����x��K>�K�$ú%ם�ƨ�US�|�1�\��<Ϻ�i@mH��]���=/��2L2�M'�}|!V@R�xk!��a�R��| Y�QY���&������9����pC�}���\P�0��'�zf�\L��7)�r�GX�Wvgc[rK���=Q��˹u�|�h�榼�\r�+���7��E�c�p���R�y��P�4!������T.1��[�HS��'��A�U��������O�^�����.LU1k�Z�{�E�+��A���%3�Z�e��W����!�/)��0�Kn��K�`�sߥ #�\|8��fsqt���B�M�Ԅ�$!J���=��Y��0�|_�H
�.�� 1��rZ 1�k�u�'�<���
p	7�t��op����Q�}I��Ѝ��-��X���<Hl�/��G�Φ�V_�jB |Q��𥽚�ިƑ�1]u��u^C�6���:5i���듵E�������s�`����o���էƲֺ���Ұ~
/�#(ğ����k�˄I-��N��)���a��y��[7ZEQ^7����Z���ɺbET��7���G�~&�P����}�2�$�0��`�ٷ�v>ԇ��9�[zn�

䦽���ȍ}R�~H�hF�p�݄�!n��Ru��p�r�??��ɀ������5�Q	+$pW�%�%�H_T��#Պ�5?��U�/|ѝƹ�𕙇��=<���#^��mµ� !��$�#�$4O�H�]�:�o�gG
(�sB�77r��Ѕ�8�Rʢ9�F��r
��6\*����2�ص\vQQ���>\)��s��0�Ù� ae���?vb-=$~w��5�����V	����[���k��fE��lj�zg�U�+���l�DfAH+�*w~��]U�L���Z^G���`K��#���گ��� �K;�k�5D����=���������G�c1,k��#�,�>
�j�t!�Y�B�6��ui/
���6w|�����`
���vߖƺ���e�d
3���_��qC�����z���R�>���R"+��/O�z�F�ןu�\���ҥɁ��Ƣ��^��K��t�k��I�d�K�jk�T�:î����jo'LE-�`��Z����WB�(W\��u���B���=O��$e��ۨ�>�rjo
�0��
��sV'�qEG�4W>;���0��V��m��xP��SN���J9�>���ߺФ<D�j/�ny���*�n���WcRP�V!�dA��N�6D"ӛ�罐z�}�}9�m��BU3Xx�$���zBr�w�L�c@�H�	�Kj<�Nf��˨뤩�D�ݮŤ�|�$B��S�u��Ad	O���Đ�ĄQD��;3z�m��"!���ރ�E�3�O)���.�r��d�c�`w��
��9��
�^�m�@M�bǰz/�� �'K`��"��nq�w��#��$1��(�zᬾ��Q:�>ų�������O���uJ�R4�_%��G���[�u���S��m2'k^�a���ka
���#V9h�	���d�ا������Y�����b�<͑U��E >,��p3���KyԹ�Fv�q||�έ�Su�r���+�ZF��ᨊ��E3z�rz��G��f��Bu�=rTOT�� S�#�@��dXi0O/a��s)�è/��,��,K��J]��
�R�1i8��2yq^�
����fi�|ѐy��J� ��v���/e��Ҕ��kў.�aF����<�d��ր�����00��rX�����0K|am%P��ߎ=��5@29A�N�C�����ۓ�1�C5���W~X	,�Sr[YN��bM���Kg���0;��2VCՎl9jt���\��?=� עÎN���i% �xH�)��q=�p3],���g}��6�O-ͦf�1=��{��ZW"Kn��?��v�0�i�~lGc�)��Q����+�هX�73n��\s��:��l�$���=������s�˸��=����N�ë-`�!�Wס:\���*$;֑��)O��'MR3u�G�L�.���l���r �S�t����k�g�$kcY��^�R���T��k�]߲��9q����'2�З�.jd�ق��Q9� �\��FM��>� ����v�a1�bhu�z�}D� �ȵ���kn�(\#@vCW���i�N��=�=�9_�7��C�7|��N-F)��8�3܅���dl 9��i��Y�(���$UI�`�>�l����\�-�IbNgy\�H�:�魐�_D:��a=9S�oу|���z�<�[+SyZ��Q�A���Øt���] YUu툻��r|�b �MA~�~A�v���Qm�QؘQb�ck�A��^ɖ�~�P�l��UB�
{8]��;.�C֒�O��N���ݰe%��2$k.F+7o{��:Z��US�Q95�A�����֬��i�a{k��y��\,$ʭ;��ms �����s�?9�q�N#*���r<18QZ����Sw�;T�����c�"��&D�2����q��v��FͰV��+oQ@�aޝ�?�=���`>������c
n�Pe؟��F5t�>�H�=xMT�ȱ3��S�L(SUn&��ڷy���.�'�2�]uI"���h��kf��q���=�L���MO��l�B:_B�����b�����o�a�~��VL��Ù�	^	�+�bO�[�#�b[~��/b8'�gĂ8�X�/W)6)/���]A��q�"�F��tP;Bd�5ִ,���Er+�y�,G��b�4}��"�X;�@i`��w�L�#�[��R"�k�$�j/j�:�-K*�5���9I�I�:�sQ/_����vY"���ɹ4�R��qX����%\�yv�4	���k@��wx��b k$��ɁS�rD�aVA�2�"�$�2���ιc�2�t����< Rܱ���q��2^���;)�R�b@�JDs�?	�5KS��*�#�FWZ�$uD�$vbd��?#+g2�w���sjB�4NЀC*��Nz0g%�O��X���|�͎��b
xM{���%� P��E��<q�]R��c������Y���$�,Sk��*�I�N\L?w����47�GD��".����ٟ-�4Q���ak��U3ʘ�V���F/`��{K����o2"C���nG}(?�t@򇆳�z�e����ZY�_p���0��	*���6�lZe�a�0�pU��%��_�L)%V��N���CY���r. >�"f��^��ߏ	�����n3`��:�݉��|������)��s��bRc>��ڴ}j�$M�Wƅ���T�lI��=����2���WBR<_\D�PII �_ٯ�r[�9��8�s��?;�4(��=��?�N����E��&�4T���qԃ1�7���qeJ�pT�ky2W*&��b�S�ԏ ���>�;� ��gৎ�����B��cU΁w��ˈ�倰䐙1ym^ъP=n�eMB�;Ud"%��G[`i���͞�Y��d^���>3L��*�5c���W�.�ΐh7�59\��2Y6Ϩ��(Z�ǡO�P�V�"�����~�+`NX��*;�ΰr��ş/�5w}Z��`����!0�PşH�I{�̖6ȵ̪&!��j���<�q��F݌/E�	EGp�X%]�gpӠ`��3��gČ>�K߮���נ�9�ʓR����vs�&B��l��y�hDp3v�f)�.�RSȯv�	����х2�)\n�lt!�sY�7�d��h�딃Q�>�3��+[�G:�3�&�r\!� v���e�}ڭGM�^�X9,������p��]�ݳ�hǼ@�b��^C�ԣ�#�R��BCXKE�f�ŀ܄�?I�OeEO��?%�=� �H7콷�s�Eݐ��s�[�?�|�>����~�wg��'���rT1�^����W�ա��&����T灼�L�t�wG��r����]h?�5�g�Yռ�#hl/��������t��Y�ҁ�2p_y���t�Eu��S���C8��!�	<eq�bV��Z���am�Jf��5m��r�ó�D��"_�ǫ�N��f��
��{�μຎ[�9�/	�&�-΃���h)��:��hP��Mw�zMNS�����/��o6_Mwq�1{!ҫ��0����BA���@6�-o%|o�������4���2� }��b�[�Ff���::��E�ֲq�0{�_�w���	H����A!��il��FB�&�L�_��V<�|T*�n������k1L�Xc�M�m��kT�ut�x��<�o�vϖ	��v<�������"0uEJ=Bz+t�Ԕ	".����G�_E�2�E�&�΀ZJ =�C�M��]A$�нlL��	��ΟhTw�B᰽ۧ��:9��!���N�%h���z\�49�7��D��
�L�a�J��9o&:��=ͱ/]��z7�X��6
��6�2���Aז��|�D�<wv��n�gՀ5TiS����P
O�S���qs<-��X�c_q�ԋ�0�t���N�[�E{�uQ/��S��7��i���A�� �_<{�w��d��Cߍ�!����k�����$؞�k'�5�OP�萀MkN������KxO1'Cs8�U�lDԦ�\� I<�Q߇���M�b��3u�sUG 7A �vq�Y�v�_�.g�h�p��u�}��r���T���m2�M�`��&}�����]�*���pA9Ύ���\���DO����_	�#�h��	\�Sl�M���ɔ\�k��xU����Fd~��Փ�\d��[��q}&�ʩZ�!7C��	��#v��]G���J!Wu0&._,�d�
53�t��^��P��;���<
��{M�&��!7��33&�մ���R�ռ��6VT�4ZU ?��w�e`��9f��ۗzj�Я�ũ<OM�fs��o�`vB��'�=��2���?���e��[^�����X�ѡo�z�T�ӑ������ԫ�'o圛�G�b
�@M����o�t����PF�,���)|Bݺ�y�^PsH�{0���4�b�������zz0���&Ŏ�(P��=�w�Aj��}���4֕��! ���l�
�%���5I�>0��U7�Cň�j�V���c��,�K�?�����i���Q���So�͞�[�C9-��Q�]�jq,1�?\�Xជ��Dn��Vw�W�x�i�%×Ǉض#��~s ��!-^���r�Y.�tò>O�$2�Ӭ��f�c^����*�4�.)hOv$+�@�`����M~�[��y��oH�A�+�~����
�Ӛ�a�j����Iث �P�E@p}����Q��'�0ݎO������x�J���Jo�!��9��|I�����'�$Li�^��fr���~h�Q�DZ��)�k2�:<ԋ�6\=����@c��z��^�_��"R�y���*|�w%����1�a۶��>��g3�<H��X>���j��m�ڎ��z:j�Im:D��y��2>{�79Zhs�F3ؼ��E$�s#��@�k�� �8���?��yP�2���l�-C�[�o�L���P�{-��6KC5QG�l��*@]��}f����c�Λ�6H$홖&��>����oC&W�zsA
@���x����H�"��H8i7���r{�r.�Z5�����i��~�Xeh��0��X.��Q$�?�f?|�4Z�V���+}C<<"�7�S���w�s�VLZ�g�9r*h>���v�[&���>ؗ�1a8�e�e%6��w��e���z������,H��{��ȝO ����+"�St��4��p1�%��+«����K�:$�#MhzcLS}{X&_ ���ǵB�����{c���|u{@+PQ���Dg���lRr�r���c�4���N�Y&
��)�i��\���$�H��S��5&�w�-� 1K�܎�L�qD��,կf���p�ی�,��@�y3
�"�
�B%�
�N�@t!b%��A�*�)�Pǩu��k�>����>/�Nf ���%��@��Z�G+���B�QU����� �l.�{j��
���/�Ɯ��r0L�Q��1�d�z���|���$��=^���-�	4�1�䪟/��6��!"����k�6jQ#��;��`#ݚ|>.�w�'��;_ҝ)�?NR��VE�XEU8G�)����~�*��V-��j�H��X�Os ��5��o�`ؽ�.��z���|��`�!��x�j`,\f����XǞ�ǳ�r���G�w�)�<���<� �pY ��Kn�$�x�du68z�08#��]�'C� ����p��g�h�uB���9!C��,������#��C�@�̚�W^3E��{ը���L?N� /�e�������.�]>���L�9�#/.T�e30��r����	������Y~�E��CE�Ԡ�O[q�3&P���_��Ȇ�4�&�R~ ��.Ȯ�	���Ѐ�nf�v~��}X  �CCES���r+���K}������۶�?9��'D%����r�Zx��Ƕ2�{*N��\l�f"�Bq�v�DT� �\u������+Xpy������B�i�1�A.Ai �~��&��g~�4���6N|�)]��?�$1R��%	�X^;�#Ea?G|�(��+9���VrV�L����ǡ�5�ʷ��@-I�N�۳{=�	Bx��}����^C%e/ԗ��}�di�e��K���4��i�ii��L"��ʘ�e	��hH��Xtmp#�c�1p@d��jz.V��ȣ!�S/�k��5ap1^�����π"ɫ��L&}�<> )�G`������4܈�ᲜH/!���?�d���]���%��`��<�����:q\�@t�gI!��L4�W�@Xˋv���	��oq�}�v��D��=<5ؑM$��ڇbRn~�)+���\m�0��=�]����Qz��'�}�� �2�Q^j�$���T�g�1�x�8�H򸕞���fK��W ̈	?�b1��`�P6����7a��~���@���+���s#ey�b�3|�` 9�b��P��O_9�|Je��]*�.,uZ>�e���ʚ�&���i6vd09�����G�:�o|�e������2	�4��D�/�v�:�- ���W��.���p�!_�K��3)�-|�Ď!�x` 7�>�	���f7�m@X:�#/�6�fٖf���[�˓o�|����ϲ����f��cl�D�T'�-���W6�� UL�gŨ���7��D^�������}��m<TN���3�����m�,���O����"�MCl�jšx��|Ϸc�Ѥ�{&_��� Nj7��͡��V�y�3��>�(��icxk��]�r���a��>*B����,��
z)��,� �8��˅�W"t�6��I��?{�w�Nfi��n�����̐J��/ȟx�����i��7"Mb����9�o���i�a��� �%9j���NJ����m��N�k(b�̎}����\&m�R�j�m�b*���J�"ƐB�
|��uҔPY-k9'q �K��j�t{�Ȉsc	�!��h���y�cb�\fy�2�?�)LS'u_w�����]��{��>�,��Q��d����ڕ�c꬜�&ѹ��BZ8�\����^S9����Rx�:r$	 EH�q�WB+�̾%�vL���Qn��G�b�b�������"/Q1����z��IR'�eS��/��	���A�*eĥ�ݦ%�R�H��a���FB���O�vO��L�(���Ѡ�}	���@4IQV��ͩ����d���z �7ckV\����=���>e(2�0����[/ǋV£|6p͋,���m�	�I�BR���{�4�{YnK��﹒�O�Zk	�%]>���+Ј�?H:j���������l�O���~�hV��MtԞ�\�+���W������r8��- ����S{�@ӻ�^���lm�N�>v:LgJb���$G��C_��!�n�c�;�,5���P�8'V!;���ފ���_�]�|�@�����KӸx'�!��hƑ��2��E�����	�G����	!�F>�c_�ߪZ�S_��ϻ��d0l�:� L$�88�+�J��-�������7Q ��KU�d*#+8�t6��u��]T0%
����v�fҲ�L��O<�Ǉ�[�p}��0T3��/�9�'Ѽ-�W�H���_8A̶wl?+�?�.X����n�`>�����.�8|>�����4P���
�l<o��9��c��a:#��������
t�fܧJ&R��"�H��Z"��"<�����pk���Թ��fnp��r�;��'%��sT��;!�sanf��5�k��T�<�M�R+�i��jOA^czFm��CZRS�:	�[�x`�a�@Aq7�b�J5�d�������H1~�f��B֖��N �C0�:ݒ�4��x#q҅�MP�I'�l=���8���qt��Ҧn��y�x!��I�;�m��������`c��3��R��h�����N�>r����`Wʝ|�"��X_[rC"�(+��L&�����)����g�H�k�z��X�,q՘D��8�`]N��~���p�B�*D�-z��/�@���5L�қ�\R$5,�~�~�D�=N�+>H�[��o�ǲ�Ǒ0���wi��fG�{m̚dM�����yyyg,��'qc,n4º�% �j�s���݉6"�/�6�V�,{���Q�<� lc�?�I�K>D��8�{�!SmZ��uΚ�5���:���"й���G�qx����і�*���O���!��K*pi��Ag.�^�tbJ|6����s���0��\W�O�7tm��?�\l��G�8�jm"W�M�2{����Xaiw�;W�	�Ħ�QVuLwN�8ʚ'�&��dVH>k��ҳ����5�Z�)4�2��}.Ln��(�x���S&SS��f#]�^M��'{��Ɲ���ܰz���Bʬ�S���%�/�$��K��#�J�b�^��E��U����X����@��I���@������="�������[��I�KYD}����Z<�6{e��_.|��g� �B�r	��`����$~����y�Z.��;9ʘ�#�b�"�DU��,�N ��5E���~6ɻ�έ�-�� �����d�O��;�M�a��_��//P�\ ]�-��H���#�ƀ��1����FY������BQ����,	��f�������&�g�����R����7=����{����o��{b
9�>wq�I3�������x�>G���I:"#��:�\��FK��E|E�n��27פ�ௐ�l��#�Bz��"�C�Q!�g��O�.os�Ms�[�L 0*��������������KM�P����R՜!c�Spb��X.�~%��S��_&��f"hs�$8l\^��@S�.ףI*�d%�b������o�)�����/�3֠ _�e	�<R�-I>�>���9������4�=��!;b𐹝�T�B��5P�CaAلW?U�i�����pu��QvQh Z���4��<���#�!v�Ne X��,4�r,oJ/���>� t�¤a]�]ݗ��TT��E����O�.�y��h�ڛM;��[��#�AGH�Т��Mk���z�H<�22ޕrg7�SB.�˫{J������K����~a�[�<�P	&V���,ɫ�/���0��$���Y�6���a��P^��dޔ��5��lsm��P~$�}Y��L��4�sN���(/��eG0c�-u��ʆޟ��>:�|Q�]%
�VWW#R� ��:'=y����`/ Ƞ����%O��6u��gN��ix�	"/����$7�}�#PZ�w�~��0���Jt;���N v~.��"#��I3��A��E�R9�\s3\A~�����!��!���=��
=7xS����HY��WȨ\^,��aV��������;����`?�?-�8gg$Ȋ�m�� [g�_�yCY���L�`_Ү�(�_c��V��˱LN�y���1ϊuů�I�$~*�r��=�����R�|\ ��j~���E�%g�.*�J��>���7%#A;�&Q�+���`���>Q�8	5D���Z-�&Ț���8N�7�OY�)�#������P7,7��M��{���܃H����W6;_r�<�-�<�h3�}�P�_���8����߁���Q���<�,�R�`��j/�&�o�]t�f�,���dӡ�:�3K��r������|�%���Uq�|~���&���͉x̓��#E�(ڲ�֒\E�u
���X�coA}�lC� ��h��?�ƪ-��K��H�9���O�������M ȑR��7�6�$'y~�7	Ѓ��\�|�,lm6�t�ͬ]rV����- }���H>�s�qA|��a�az��Μ����W�,R�T
���A���������s�aJ�Q�!�	����VU�1�HalY
����i��h�R}޶�41e���$����9`@�893i��/���^Wjd���W���p��r5�T�C���&zե9�p�S@�4��iZH�,�������l���� �A��p�K��v9�F̳�������xt��|_���얨Zk�>�ݠ'���[�H3�_��bh�Q�=�B�S���2zѝĀ��GGյɣ�?���>�l��EQ�R�*�cR#|J�=28"�����l.�_�����JP�A�6/R�O�D������X�+$�D=�������+Y1�}x�:odɘ���ib����l�Nj��Z�xmK#�.r���N����{�K��c�����B�'B�R�62fߚ�A㹏�)�[fa�ia��k-yQ��+� �Iރ$jϏ�/��Y��3R�;���txKd����cr%�t3����ef�Kh���"�! {!����m>�J}Lh�#��@���x����>��Y
PR#e��J9�ul����dYe�R�w�&C�]�B ��T>�ҭn�;4H�E�K ֍K�J5����y����o��_�/���6rF�C���5���Y�t+zE�QK�oM�o�
����8�9z!f�3�M�c��7^�
W�q����eFV#ތ��%�`�f<����I~_�z���G|'��D=M��)�5z���^/��1��Z+�/xd���GD�"�_�E���?�9B�G��e-�qnq���Y�D��C(M���$%3?v�֍�������pcIn�+��a��z��z"����0�>�3B׊k��*�.�-;�p�n���r��#3��vM�݁f�Tؽ�4ϣI��}�}���nV L�+ƅ�~s�1T���*ҙO���H���I�@�JrB}��q���V��e�O)�
��Q���|��y�	����ɷ�/)ٍ��\Z�`����jۜ��V�Y�¹�DʼP'\���#lgϑJ`�b�����*�D~)�^n,K�ǰ��2��6��i�F$�.�n��Fۈ)��'�k>��C+4�
�WOyE�%�s�`���d�S�=uE��@�@A�6����"�������?����vI�C@����:��V�68����Hvp�5[��<�s2�㷑�W���$b1;e���TC�p\����F�o�� �(K��:
�-�5��ڨA�������+s9࿿0� ����Rf���R�Sv��m�u�
T�P9