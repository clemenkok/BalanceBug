��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6��&��@�l�����[cC~	��Iq*���8��%�6®l����PT/^	.7Jj^][�F���3p�}5���tj��L����W��v��*4V3XԊ�	��cCE�r��6�#�HL�UN|�\d� o��Q���U�oq�����s�m�?��oA+�eQ٬᫦�v!6�56Z�E,�*�s?���( ��I�|p7��xO`�^��BUy�:����I�=+e�,�#���;�pI{�Z��u�Y��h4)�npު�Y�NYKT�H �[D�.� "T�bNa��Fj*9�3������Y8�Jo>xH=�U�^0�����ɚ$�6�4u��H΃9�
=�(a��p�0��0�M)�3	�ֿL$aHK��=n��H4#3��kd�d�f�k^s	g�a������F1Ncv^��ǁ�'��ص��,��V�wR6�ڢ�¨1�9e�
�=X:v���8̹S���*���p����Mb�]�L5̭G���EhJ����$�U<F�X5�^>(����eם����Db�>{�Љ3R�*�T��nO� cO�8#�;���9w�~�v�V��@f����M}( �{���V3�;rW�OTcv��gS�2yh^RϞ���s���M�i���+�T�7:e*��pjv��FhqL�*_* E������X�p��H�]��ē����Э=����YD�5_�>_��63_n m�Vdvyr������׍�+M �O
1'5+j��7n(��A����ɍ�fP�w�|���Kj���%/�~͘����LR)�i��~wh��E�'}���vj��	���e7֮`� t���VGQ�z�
'&���%T�)X�������D �����<D���<# ��G3�����.읛q�_��6!���e��dd���ġ
{@��뫺_M�Y�����y��}PD�˜�Boz���Z�'�l �m�v{i%6�7f�kI�F�.�:��9����-����Վ��́�8�?E`8���F��$�����_l-`W�"�z�,�(0D���l�d���ZH�=K���)��?�%Z�I�x��a�D��(��#ܕj�
�~�/���M�B-���X-~֠����,V�3ywӗ;�])�Ɯ�j��F�IeF�
L��e��Ұ�Uh�$���TH�l�U��A�� �a~���eJ=j�K<�;b�i���Ҷu��{��ٿ/�UC�Z1[XF��{1%,�Xr� ������W�%�kb�+�a�t��v'U��K.b�²��C���ޯ���B6���I�'y��q]d#!�<LdY�'���z{_t��ܖ�u��N�̺0�x��٥X����W^�?�s��{�*J�+l�:���]�j��<=:z���$��#��V���#�ﻻ{y�ud����Uq "b�%�/�9�B �&	�'� �IMQr+A���P���<{bI�����=�n�0�/�W.t�RV�-zaa����ʹIQ���S ǌ$�L [f�p.�[H.����Y|f��ą��`���]}�����Mwp���T�m͢���/�P]�N
 �����v��!5���]�{���v�O�F�|�3��䡙X/�_t��9J�FTV��<ǘ�p�Ǹ��j3�L�Z�9��0j~xU)u�3g��SJJ s��8V��9��eJr]��̎ސ�TK�o �&֛ן1�4�M��_����	��Rp�e�e*E�������
r��z��e��%�e��-Ba�����+��/�	�_5[�vrH�yW2ϒ��M٦�̰���~�]2X�?HA��4������3�x�>���j�Rh���8*TN�♲����=Fo����h��{(ا�5r�cX�R�7�{������ֹǗ�N�o��ý�� y�{ا�9��!��DH�8�a��4M�A�f�qH�F��bcw��y���E�TC������4^����Ҙ�U���*"�ZKq
F���;��:����f6Zu��s��>��Ѿ���5�FL�8-�@�'ǂ�'��Ƒ���n�T�[�l���V�p�C}������#>4n.M2<��s9B1��_j����Q�o�6ˊ<B{�a"�=��IdtjO,��!9��������f�G�;O�ED����`�t�a����H��pEfy6}�໯�l�AE��H���=E�	��0
�kP�����G+,�b����RT��h�)�~�Eu4�#�ξ��3N� T��xgK칣�Q�1�a�`^��kҖ~x\�?�ܭ:�8���=�.ۉv]Q3g�c�ד�UP�C������CN)�)�l�J����?���3C�-ц�ЪN�F���3��ҥr�
}�3H�%�D'5�L����C���s�6��<_y�����n����|c��K�ErRh�	�?�|�ZV��e%���R�z�a51�g���-���%��-od;��H(���^S�8"g�
���u�l��A!���'��Y�DT*
/	Mޮ�bf�W�f1
#IfY��J��yDx#�h{�_�;*_�a-��x�i�R����s��/��7�ҕ��sĎ4�0�/ѝ�֢�Oj�����t�Eӓ }��=+�*j�� �<�h�x�U�u��>yy^��V��t��)�tM ��KsV3���kn¨�������4_l�ր��gQ���4v~���[]�s
��}��R���C�30��Г��J���LX��]$��n$9�H����*1�W V�@�9
@�!��󖴟r� ;Ǩ|�OR3�i4��9�9�3�kۜ��~�L�`x�s�9)�f1�ni��5�:���0�ײ��v�6�dR��ea��6�t*[����X���ΌG,nZ�>B�=!'�-+U�-��\�=���H.�Z�%�t��f���xL}e��ZIH0k�S���Gr�V�����$�V�c��?��#���Z����3��}8}�3��D�-h�M�<M�n������5��6��kZo��=Ú�WH~2�9(�0x���!�R�' �[Ӎ�	���\�mv�@��=�!�պ�q΁���0��y"X��=��}�
3�:g^� ����QW��>B4CK�UW�[A�'�������;+8v�Ȃ��,~�a���k�%��оW�|��ql���gU���$#��Ap��A������dd�����'�y��'I�F���V�+���0]#7��.N���5!�5����A�M�;�(�q�͠�?j&�m̝�{�SU{%�%[�m�V��|Y�}!$��m:�>,���V�5�6|�d^�K���w�A�83M��wr�>���uf˚�J��PeT�B{�-K�Z�y��*��nI�%���?���Cm|����?]oV*P�|$�s���g�TL-�3T#9ϋ?�G̢�����7���>}���L�s.����D������F6�z�P9��S��5�;�Jpb�[h�ޣC�}���R���ڃ��D]�����b#Wmjī'�C�M�=��/No�
�a1#���AQ��s�N�=e+�"�ڜ�8�fd�8��|��:�T�G�&:�M�S����~�R��	Ikw����.ָ��f47J��s/�،��ƞDg�fdPC3h�/S���v��m>�YZ���ky��Pk��w�i������� n�Q��(BA0I{���Y,ekG7]���ا�7�;��c���Y�M�*@�G9d2j�[Ԁ�LAb4p��5<!¢�5/{E���M{ �kVazC�ׁx�VJ{���$݆�j &Q�5���~�혦���v��0Z S#�e%Pd�����L���{�Ӱ��N0��w9ps��"�J�/�GR��3m�_���!����'��K��֗�(��F���ܑ�0�y�_��aK���NA+�A��S�����v�W�Ib�1{ �"���ោ����ZF��$��W�IA�,�%gly�9A`D��b�;d�:^֜�e�~i�2/�=LI� S���ǚTW�|M�}4�iL:�[����'���9)padEY>�Mi<w�(��|ݼ	�>��	*k6�$A�T(g=P���݆1�'3�:�\箷/9�
x�E,�p��6�j��<�r��a�,����76��7��xB3���߫>c�8$�~|ox�!�P�������r�]DD�PBA��6�.�u-�Ch�j#�3���Ylu��c85(=˖uc��/�ב�s��<\��]�Uug�r61^K��rφK0��x3���'˪�/�R��)J2�T-d�5eX���2�.��К�C	#��d={�k�3�L�x���7.ʴ�{'_�vB�o7P�`�K�?lt�����W�~��Lz�����|�vB4�h�Ve��@���<$�@�-M���[� �4ŀ��۳G�)��b�>ܖ�O|Ҽ��N�uw��F���==��ZHӻ�_Nb]w�n.�HTZ h�aZ���3(:]>-��,��Zz	:l��x�گ���8�z�uWR� ��']W,��iM���&��vG��^�77T)2����@{|Q�m*�������h�_$���^�&$�����Z/�4ָ�����Z�zV��"�>U�k�B%�G�*4��M�I��WQ>�q�t�	jD���v�M7Ȫ�"�R&�3��B����ͅ2ܦ��#4�'[z{���	�D����-�vԄ,Q��:���3�W]��c�L�K��W�����aEP�RPq��)Յo��P#�8:����U���K>���	ϖ��U�܉N���=I�r�el�	�?c$��S�C9��Ҝ���Ib���P����c����W,���d�������RȭnM�ܺ��!��jU^�M�y�\�h�Xo:^��c��ق���%`@��7��}h��V>3Ж��Y��b�:����d����8[3�Kϳ��e��&Y���y8]�t͒	./ş� �|s+�8^ډ;�M�X�9|���Yh���{R:���O���Q!�P�(���I�+17�\�S��)���Փb��0���M� �A>��SV:��Q�`��� ��T�����W��(�]�U ��q_q'�-���d�x����o�����o��
��=R�B�Y����g5'zƳ�^���Yc�D�}0�F+�>���tRFU�i� ��#4��S����N���X�L�Ĳ������DNp�$�e�c�-�%r���Ѹf5**њ(�k޼T�f	܆nGt���!�����τ���|o�r7+sg�m0��ж5xK��ŜJ���Ҝݹ��6��M�u���4�1g5��������B�OK :Z�4(�	Gv����n'�ü'!,d��Q=�!��y�pA �⁊�r����q=<E��F>�8uo��f��Yl���e�LFPq�D��<�_��SED��$i�<���u�+KȌ��ʼ��ɑ�/9�R��*�i�A�7y��O\�K�$'F��1�騞!��~Q�ە��JvFXv�FG3P��v���y�z�vg��E���Fz𚬏�Χ*d���IN�nmCŏ���6�4�����v�ZJ��(��+"a����^��@�+�
�[9�$��{�����;�A���_����HRݔ������d��{Vk�����z	�'���g�>� ��ΟT��:Ll�i^�{�6�h:	���rM(�k&�B���/��_�q���r��1m-�:όz���a����*MĎѶ�7o�c���`��`.q/H�.�}=$��!��$�����8���u�9w�,^z�a�Tu�
u���J>��l�y�r��!6�]�r��p�8}T>خ��������>P��i�⋦$_Hk��PY	�=;�@D7g1[�>���ۉ�����e���`�uE���'���n����>{}ؖ�P�?V��n��j���o��[��8#�X�Ν�ݗs��c{i|l�D)�to����;�1(������_��2�.�2�W�|ӑ��;����Oo_�B���k�4�~x(��{�^���;f�Ъ`��z�D�ʌCͩ�
�c��*O����ў�y�U����zl8ے���枯��N����#������*�U�F�b�W\�'�����zIFH�*u�I#{��
6�e�z�����>�{�HSaj��|O8�
�PX�K��8Q�G>���-D�5�R7u-�u4,�.L����V���l����_�n ��^�²ǧ1j�[ܪ �V�=&@����ף16����&\n�\��L�K��u�j��r�N8�_̨ތ{D�WeMI(�˛'9��
9k�Q����"�^����� >�\�(��-��^��I��
�(A9bǪ�����N �ը����=�l�_+^�P�p�mB�s[�st���㗕�N 52�ob��>�_a&	ۭ�i��3@w�+)}�kLŻ�4��ѐ�Y��kп�΍�V��0>z����w�G\E�$�h=�4gYȥ�E(1��ޭ9�/�C�~ n9���f�i��]�㡞d�[ruE��un�	�e�$�ǆJ�s���aS��K�Yӓ�I��ׁ�Z���T�M��-�Y��p�JOH7�������c�MA�� �������h5yj��"���L¼}�����D���# Ujލ������Ǒ4�� #�T�?M�'���g9iY�:-][d3D��W���`����e�S�:X���)z܈&�ǘZ��8\��)a�|���y�e§u������2�Zr���t��RB��������R�L�o��^�ǃ�#�0TW�9��"&w�\k K��%������k��Qݣ�d�-�Il��c���B�tj�q����ϭEY�G�4[����;-��gf[h�Pw��65���q�����4%�cit�'��8������#������,�P6ciӰ���b��c$�D�t�= ���kD:V��ˌ[
s��߰�z�h�c��VgŚ%����mфl�k��~#�ʔ�?O|}>7_7V���ə�p�C���	���r���1�����syɕ��s���?���˚=��O
��rc?�
�׹
?|+�Hֿ>���,�X-���+�Z���b(gX"a�R���Ko�6B@ <-n�b�6ڈ���Y����|�ǈ�\�����F؅-�uc<_�:�$Vh���I5,s��7hXr#4��*]�P��h8�z`p��
u+މ@�d�2���V7��g
�>yd��E�,�6�p�����Qp�G��I�9FS����C��)L�i���\��e�u�W�9]��]��?se���0�P?�=ىì������)�}���q�|��3�2Ҟ���zxMF��X�����Ey��>t��4d��A��Y��p=$��%�