��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d���麍�Ks�%$����+d7��/��������ߔ,���<�E�]��&��z>��>�X�������kW��B�>��N��e���e+癃v���"��Qv�謒X�<��9Ff/�H��Y�m��{oݜ({l���;����{'W#���F�`��s�QŗS�'��[����7�5G��Ξ@��/6����=;+�Cgt�ܫ����ߥo��yqa�ĝ!�G�F#{5� �E؃��\il����A�E�sƸ��]��i��Y���i���	��'i�6�9U�x� ��n���}FA3Yt��SRJ��UZ��	����\�\�t[�oA��g��m�o�I��뚑	�u�!y7� С��/wn�31h�O�3�8w|?���oh��m�&��}���Af�m*tH��i�U����W��-�JһS����si���Z�v�x�謙���FMW�K$��r��R����-�OMjK>I4H��;�a�3�a���D#����X�ç`j�h̼!�W��V2?:8�k�������%�;r�N|S�v	:�$��Y2/
���������K;%V����������:��*�
g�
fIRG�/�J�G�jM��lS�H�.4�U��W4�:��:1�*�h�C&B(|�y1;}��?�L���8���9g�afP�- 7D�.�^7�D'�{���>�#[W���J)mjY����٧j���M�D}{���پ��z��<ȫy�a����g�`�y�}��D��m��)�9Z��l�6~o=�C��p��m���ȥ4�Q���zX$�^k�E�ve���r5����Q�0�2IL�Ps�3j�v��ΰH�\p��}*���z��OI�"d�S�؊��dd ]�&�����.M�'���~�w?�2o'��9|������}��#|�D 8�ւ��-3!T�ڵc�ݓ�Ȋl���>r��蕵�`ümى�ʓ�W��$wӒ��aM�Ɇ�5��ƴ��E��	����Ӹ��A�Q�VJQ/3`]��(�d���R���.��7�ȩm����6:�'|Q��b� ��\j�F���rk�fKF��޵e=�,�*�?��Q{^��9G0���F���K.��j��0S�IH�Mݤϕ����~;X�jp����<67��dM�Z�f$e�l�����Ǽ6mI�e_�Y��p���*�6�����"ľ��$(2�#2����@�)�`&\� g}+�v�ˉ��DUy�����q�q��� �����E	��0�xO��NZ�짔G�v��ή��l���>&��;M���rW cE���OoR@n/��f�;�G��N;�.xo�c�Ǡ^��~|��L���^���H����=3-V����ÆR�'��]��`�]q�1�l7  �G��S��!��%I�+��<zbA^鬩\��>l`����;m��
]_5~Ԩ�u��i۟̉���F8̴��2��@��n8����h���y�E��R�,r�,�
�4K���vDY��H!Ds[�テa궶gN��ނ�-�b��G����ty]�|0e�������+��D��_�^�N��U%� 2mXJ�9��)r�ȼ	��C�0�~���%Z +�@�X���p������QA'c@  ��'d^���%���w=��I�o,�/��^�l�t�d�~fK`G-�V�G��+��O
��������&Ά�}x�#�I��}'| �Y�<�?���	P^��(]����E]O���'VL�m����N�h�k��F�� U�T�� �P��;!G-��*��8	�a��*�wK�0����RgP�bm0ѻ3�l����9��C�b˘�h�!qd��.�J��&���(i=�꯮�o�P��PX��ȧ̰Cc�|Q%S8w��	|R Ƥ�O-�����@7���9��*a�N��副/TQMݷ����'J����6�7�\�o��2�:�3VQ�vi8s�uK�" MdU\ǎ:��÷�3�i:�Nӣ�$�r��UM����U:ɭˤ0?�t���ngq��N3��W���}l� D��5PM�	�r������Y>�k�e�1�i���s��yc�M6)��{i��,=Ԏ�%����9B+��4�A��p��{+�����6JZ#b\6��������M��[����_�U!7�Z�|>�3D30�R�lE��a���[���a�۬��lvHmAn�jx0��9�~ju�,׮ǟ�>yf��l<��[r�2	\���)I��=�7�sn-^P=�D�.�G��#H�~)c��1��1Jx��=��������f��CX�8?t���j8&y���NA��8��P� �B���b��������TnL�����o�ހ�^�L��y�}X�����	P����P�����:C�w�܄�h��b�Ǡ����+�J�P���ƨ�����'���K?�"R^�jT)~�:?*�@!��WLm+@�6�T�j����ÄT�-��%4A��Vh-�5��2P��7�:z	V��5w����:�k�G��I�:�h��Ge��&��� e����YW!g�Lψ8Y�Jg�;�)����p�x��3?��a85�)`x���F��:e��g���������V��}~���(�˂��;8�0�/�OP�S���;^�*�Rr�J���$�+��'�H3$�]�$UP��)��e�p�C��' ןKf�E�$���2�gRu���Bc�s�eϛzj�Em,uΞ��BU����f�X����G �S�\j�Qn^�n��[ο�qb�r�Y��*���,�M�fV���^�����P񱆴E�<'�'@��#ӯ��l�����.����Qf`��a{2�c��O	]|���ҕE�	
J~f��u�B����UV�P@��[�f�'O�l�)�~�vτk�ӒF�)�뮚T �S&�(�~ǉM6�#�5Q���~�ޏ�GF��������oz�t/J,6Th}EN åϝTn��sH,��vz�C�{�js��[�|�^'�xw�<�ћ�ړ�2�-`Dg��igj�Xqɣ}�w�wbO`^���f�1����q��0����o[�)�27j�Lm
>�dT�<�s��ɏѡK���آm.��E^�U�'�q���dɁ����r���-l�����lˏ@��-�+�J�$x�.7V��@OCe�f�7���h��/Rt�ձ�L���<
��l]�$��X{4�m�0C��<��[*�y��52qpQ�E���]c��|G-U�8��T����nM�H�Y���_�����y�o0�� ����5z�y[�v#��{ЎQ���ԕ�l��<�Ƙ���V	v�7Y2%��[PdԊ��PQ����3���&w���ܲ�ټl� �J�:�o�靖�!?φV1Z2ʭ��x)��h��=�`d�V�(5�MT�� B����4~��z7�zp��&:�+�ؘ��"�ޓ.%P��~��!x�/��s~\��C�bSTm.�R�͡�����S/_ܭp]sŲ<��3�P��*��Tg֝����:Q|:λG"��-כ��1��7�E����oQ���2"�s��v���� �c!�b`�BqOb�K�ZF_�9I�����_~W�}<��}�1��֣в��3L��Λ�ɐ�����T�B/`-_�A:��o/N^:EI��b-o����Rه��ĪwT����L�|�@n��|]�w����&E�zZ�[NF�<��5��� ?g�#{� �?�)0X�_ozK ��v�3l,� �h�.����#(]�a�T5`�~_60g�ɦqNR:?g�E�&V@���F�9E��SBY��Ѷ���7��%C�7��N��r#�r���_˾A�.z���k�-�Z�4u����N�+��w�{zg��|?��Z�Zt�ߠG}yԱ��4s�ed;dn��ښ�S�Wq���X� ��lO���=�f�h��V�?p�����(X�:�R����
/k����N�J �m*��_P�<G�?3֛ʘSHA�e5�@(ݼܩ��r0��@C%�����_�a>o[���[�$r���'3i���OϬ�p�4q���ʝW��$u(ȳ�PW�aD!Rg�$���2H�]��M�H=�?fw��`k[�z�� !H�J�V�t�&]����q ������3F\�2���
��p<"�s ��ƫo��pa�l�7��eQ�a)�-�?k��1R�Ef\�2Di%�,��71�2zA���gg(`�A,7�U��E\I�C���}��y|����J�iXt���$��������w_-����\�&��8��#��5D�B�ً��?������,GFN(�H��2ֱ;̭��rq8�P�;�A[�_V���\.�t|�nm~�q�j���>c�Im ����d�v���.�Z�����`�̆@
�Ô�pk�o̴�,A_�BI�mK;גѣ1H��وFɞE]'�X�bTػ����>��.���������3�6��t��n���Jr��;���n�s�6S[�5�09~����<CU.$�ӫ(�;2��Vj��>��~I�Xd.N/7A_P���IT���6�L�KY�wx|�ʛ)L%7������6��A17��y�#E��M�1y�){������UL-Q,{� �=���K�_N�"����� ��-�\{�Y�OٗL�����>>C�W )�Q��	l�oXG�Y{�'U��Sf*��Wh�����Yف&��
n���P�8��C��@͒�k�&�-gR3>MZ:�N�����1EN���9h�Թ��ZN�W�b�g�2��,��,e��h�'$1����e�N:Ôu�k3�ciy�`c-��nt�� �B���s��4}bb-Sh���t�<NNY�\<��d�)���$S��	|�H�.Kk�ˊ�*o=@�TJ��O+f��E?'��dz�m��o	
?�W����ʢ�f��Z��N�:X�^���.ܯ�X�8�ufFQ�'�Cb+��!S�֌s�n���uE�
]of1����p�sr�-^N�rcBDD��ǳ�˿��p�s��*?����0�Z��%K�խC8y\�[{�8��Kư�v�r�^�E^L��~9�%oBD_iK���l���������:׽!��0�H��=�}�:�fr��edeNCz�TJ�$)��-��;TP���?7�쳶�̏1�I�X�{d�TAs���Ƭ���.=tv�`D"8��K@��>I�FɷR~ ���K,3�h9��|~gHl�9��܉[�Oɂ��[�G�о�s�Z-4��\ƽ|
���}[�l=�lé��v�^%�uwL�=�	b����Kj������Z��b�	��J���� Y�m�94�zJ�:�T� ���e��|�;�	�5i�%��e�M�A��F����Vf}�<��I�y�ȴˮ�-k���S�:�Ha[�NU���3��SV, ���2�;D����rnAq��xHg�$[���� ��h�_k�J��	�C) l"� �:,@�~];����F���#��P:�,Q[��7g��h�wH�rqN�:##mc��r���Gܹ��QQ\;���������i!H-l��MQX*{���6遅�5�>�+'����������C+�2Ow�U�\����ϲQ`SG�ɬ]�b5��V=T#jpV����c���]IՖt��շ5'ǤG_׹�xCˏ��_SFp�X�UP)m�B��Nw&w=	�6��T�]Zi���`�_�v}Qge�,���v^���Ϝ�ޣ�v6���L,�*)T�X����Մ�!����	V��n�h����{���.:ε�	�K��a������nϧ�O�F���Y�]az�O��8'�jQ�պ���]��H�ó�3�Dl����y�p�)E�dE;��hQ0��7�&Xʷ��}�5�\O�ST��8�ގ*�sco|-
��ĠV!��\��aO8Je=DM�%�	�7�UHk�$�Q�+o6��dd��F��Qy�x��2-W�PB���[o��*�)ҷuU��De�Һ�c�#��>������J"=� `A'��Py���_Dsx�O
�1?LQ�m���J ��Ơ�\���C0����-���}���gQ�]_&NK�D�=��	� ��H�,��Z&�3M<����x���iw�����"쿝b^v{}c{�E��|�N�xՀ��RJ�>��/;���%Ň�*}����[�5Z{]�l�RyQt��qt�{���B�W��M����ɒ�9�ܷ�T#��(b��3.�]+zXp��g� Gy�d�@�/@2�fz�Q�˿��5��/1�(z�A�*�Xb�2�4@�����z$#IF&�-'�y��=uZ$��������#��䤅C��'�
r�����ADv�/l���3�p�%����㈫��K�J�3E%ng��5�"�W��N�|*ɌǦP\+�R9������(�u�1O�Ÿ�����S)�D� ��0ZiaV�fX�~��+���/ݯ�_��6���.��ENǩ`�O3]/嚴�Z�̔	�'V=���c,�C6 ���?q�	�G�UQG!G�ߎI��z�ۧm�_q�Z�U �.���뙁�,�Q-q���ZTr(�r���}ñ�bE���/���1e~�e�����8`�g� �����s�?��D�3o�L��y?�1"�Ͽ�(�*O�7ZRb��o\	u�܂^�Z���/Y��]GF��|�s�o��x�P�Zc���Q$
��&,ؒ`RmJp#�Z���K�����u!�L#��qF1�bDW/��NcTb-��~XAS��WKJ��s$�O��/��ϣ�nW���pj==t���j�����s`v�q�yU,G�f0�uj��1�۝%��u�����B;�#'0A|��k�n�~bR�(X�d�N�$���)!˹�'�+�mTr$��w@��d$����Cn����k��7��콌Ш�eDMN�xB3]��ʦ'���U,�~����DZw�� �ȣ�?G��:�ʈ%M[�#���6������Τ*��K��DC���O�o��|l�c��mYA�j`˒�.����񋮏�yG����q8��<����_��!���c���1g
=ѧz��h�k��HY؅q����\���q~:�J�����hӶ|�o�R z1�J%���O^'P5�S�T�B�ԉ���d&�;�o��lY�Ķ�q�t�k����np�E���}R�`9������8���rd�?ߋ(�m2\16e����2$G7�rC��J��S
�ʏ4KV��u�����ҵm��[�ۯEU|}Z7�6�@l4�G���J�+�����<2�#�]@�l9Qڲ�C���R3�x��w��FV�U:7�2`N�7������U� �w�#���. Ʉ���Ι���.X�0�,t�6$X���Kp�k�y
醢�+��(��U+.��gyH��Rݽ��)�֠��R1]��w��%ƖDm����c���ù��ݵЯ�d"�I�JH���ٔ�m>w��� g�ҋ��"�k�
��]���Aq-�-�����VX�=z7�l�_aK7m3�o !�-/��4���~Y/ek��F����m���&��=�����g2Z5�G4Ew���F�WѕJ�
�2�c��R�c^�b���Q�Dռ�p��g����@hG�/�{t-h�h/����R�6�e��jBAg9��-�TTA�V�JΟ�n9U�ķ��o�7�)ị�<�.�R	�YrP�~����k�g�e�����To���#,>K�Ik�2+AzXf�%�D~#cS9�"b�4
�*�tÿ�ü x��T��v�5��x/'!'f��qƓ�����X����u�Q�g�����(�D�^�rM6G�Y�����]~�2�u��X���2|b��@"|}�X�_��/F�8_�8]���IH&���-����C�X�ĭ_u)�'����<������͘HQ�5V`��c�m�@!�lY`\�d�!��|�C�_��e��&��q���YL<h����=E_�s�wXז����cE.�$2ȸR����ofw�2V������%��]��
�����tm���B�$*���3���3IN�9o�`���J ����u7��B?7�C��k�/��~��\��-e�Ce����uv�P����B�hG[�G]|*��R+���f'7i	ns��T4��	`v=y��z�����pCT,OQ_v]]�&��aDu�����X����ٰ�@��U������o����>}��>u�	j�&"Wߝf�]�:�Q&N`f0F�a��+&�������(z�:�y�b�����P��z����]C b�\�N~F�ZO�S��3��͍�3D��y���Z@��i�0�2��:���F�ob�R��$ɤ� �W 2���7]�{��V�#ELlǓ�k]�oq�R8�Y���� .�kY�2�Xg/U�єt��*f��=���  P|x�9�ZLn{�Փ�j�ʏ&.Mu�D?k;<��K�`E.#8�$�S�R<�]�i�K���G�����3��!��wrM�P(�UM�ٚ]/ڛ0.�����\�b�� ���dO�S�o�eܵ�#���5E\����?�ֱ;�k�Ó]%��~�<H^ax��*��Ϣm7Pc�'�|f�g�Nh�G�1,����(�B�m�fy��5�vH<m�g��h:�wF" �g[�� �����1��	򕀁���%P@Y�TB�h�8;W�t\��eH��)�xl�����R�PM���a9M~�3V�R��گ��4�����;t�7�b��$��4ֳ|1��V� �,��8A�f��D�@A������m~-��v�E:*��,�_� ��S �g��2K/��Z�	ރ�R�m��D�d���r���GfY'|�Π����X�rk3�(�㎶c��@Ѹg�=���� &>����1��N	]o�7�[���xǄ����tg��%v�I&qӼ�	oމD�
�L��kSt7���d5�s&��
U�Q��AK5�Z��� �1�nA^�$�����Կ�۞�v�?�?�4���.�	�w���T;�J���"|M�~�������`��o���ڭ#
��z�O�?�{@d,�NkC��x�U.�r�u���p�ڶl��ao�C���n��垖I(�Lfi.��gYpB��zt���}S���2aՌy+�x%�f>n�� ����0-@'�D��#v\��w͟������韨3[�U^�,����p�apM���k�DZe��@�� P�̍���qAA:�N�<�x�����hCUo"�;��{s����6�Q;h�Ǧd�s*�e�a�`�W��e�=�l�C?�����5>^ί��m��̽��;�ms$�WAe$���Jæ�E)Uy��V��uW�=�Y�|w�\�$��0��$��r����Ѧm+A+'z,L�pF`�tk�
4��e�A��ʤ����o�y��-�k�yY�g9S�h03��nVփ���u��b�,�#�\���ͥ��*���P��/
�v�A?����\JJb��W���F9'�Mʨ������P�f�1igOKCQ ��Z�~��?[��j��?&�6�ɬ���@�i�s5�#��j�� (Y���j�;�Nk0�Q�%ܘfd���&�7�,��dUTn`X��_�xd2p�<��K��K����uw�< L�($�c���/��D8$����׍B!��g[ʕ��|�2��n%�P W|�2����>}YvI�.${H�_�G����=������ͤ�9�o��C������fa�	`�����7����%(n/]6�>���Y_�}L��J�*.����8��h=����!������O4�x$e���(_�n�rc);�l�Rz�R0�J���ȝ���3�!����d�eT�!_@��H-@��
�$��>|��5�*x̓�vv;��g*����h���CxsY��O���$�*���0�[����q'�y�mz���YT�"B�
m�B��{EUK!��tAG&1کM�q����@���S����X��]2i0F�+=^��M}�B
���ݡC�޴�2G0��[8�ς��J�ʉ�<^�����I�F��_���-�9�E�����Qe? *�tVv��1&1�~�zV��^J������J�]M)!9^�n�]��#�8w�B�\������oDP7B	Ǎ�\/�(���&��j�N�9l~���-�rc\�;��N�����D�[���8B���J^KiVw6�}����⪷߫b��s���
qT~-Yt/���D�!�s����/��w5������d��epb��<�g������P��������V!�y����2��x}>�ض8u�tw����L�F=�"[A`���@9�u�SX�м�0��鋗R���1����ro��.���)DZm��gC2�)8 ��\��h���n{m�Ү��j��
w����]�,��3{s6x�5���j;�	Ц��/�3e`����{�O���ΰ�)�UR��8������YA��6.�rЀ|��LQ��%��&��@(��8�lN��g.bܖ��<1D��s�������] ����!5Z�_J�P/e��~8U����"D�4���X1F�t�{I��ܞ�Ǘ�z9ee^�5�n��γ�k J<B"@#�]�@�}����' �_t��AjHQ��%@�R����Y5�uM2�E���`ZQ�ʞ ����s�	�Ȋ�~�De��&�
$�|Of� �W�$V�R���do��H��q4�y��"���"��Q�p���ʟ�ny���D�-�W�WkH#�w�d���TSYE�U�K�)�瑐�v�+f���lȫ]&�*B)��tj%���a�5)�d	͛�#|m�b^��3��|��9�J�s!g�k�Y4�)w��=*"�+v�"�a��kQ�;e� �"����Ň��PB��B���xD������!�r�Z��PN,�8������@z]�'����j;��e�'��`�I:�	���X�	���s�	6��BGf�ok"د'l#Id�y
��\���xv�pAj�h�lXlc	ƣ�I @�0����K׸�Z��派Q'�Q��dkΣ��)����9S�8ޝ_�����O�I,~a����0���.�Rf���A�������.�g���}����P�4�QX�������D�4%�訛&�"#�Cb���`��g �O�E����.�v����~LER'�����x9���)��������L�t��7AcR�Zf�u��;��sX��E�𚻝�̢��/(V�PN����/= �PE����hmB���!P�=W���>$� ���
D6��"P�=�=R�O��g��|�mI� ��� f4��� �nd�-˧�t%R-�l�'M�h��?L���\V\4�v�qO��Ց̍+��3r��y R��'�.+T��csD�����PƼ;�M�|���L����JSJ!�AXsH��V�͕�*T?�d���0�4����x>�J�g��~c�y;S�,���[^�_S�$X�)�%ٺcEY_^
�4-����
�� �P����"\���pL�I���杹_ayU�z{��H�\d/��*4R*(e�7�πT�R�;=�X�Q����w�����%!�)H��5��t�G�^����Уr�VݕL���2ro�F�`lt̰tvM,���A��T]���[^���#�J�ٚ��e�w-�?+��5~2)�`*��tT�R�L�յ�w�t�{I�j�T���	Z�.()�_1��+�!S�N��6+|d@�i
���-p��R����  u_�n�-h�xC�JV!�ӷB�� ��\ӼC
�)�h@Ɛ���\a{XH���Fq*�(�"�U�+!�Ұذ��l.�����%�ޟ�C�z���]��wZ����eU� X���I;�Yb�b�g)���GɊ_�~`O5����$��/wfy
�o��D�����Mx�CE�E�^��P礞f��Wޣf̱ߌ��<W��5Dځ`�ur�IU?K �g���'���dFh��!��4�yZ%���ϸAM��1�Խ�IbP�:�.��ӗ��N���F�T}�⻺;Q�L�b�l������.�(��0j"c��at�b[x���1�H)�A��0�/�(�1� �a"GȦ���L�cgo�Y��'xH@������������=r��Wzd� SiL��!]�4�gZ��
�>OO]�%8��^T�����Y������u	���|jʀ@��7j��g��n�r�M�1��VM���0֟�F����*�Z�C�ׅ`�?������Y%D\�͞�7�)���bs�b�G��t�9�;6~�h��ŋ��O0k��ܻ���w����C��Z�BvP��<!�u��/9!�E�G�V��RgaWp^�� g{����>���)���A%gh�:�;(��L ª�Qx�. G[��Pp0f��.X�qN�z?�^.Xur[f8Ƿ����!ߑ����X�i�eM!Re�v�G��ў�Jjc2ٮ�w%vFV[|�V�0�m9���]FehD��,bLt���i��7�l����}c?��z���?����2��k��!��Iq�j�1���ʷ�9��@@�s��B!�m����;�'���� q&��f^N��+�
����?���˷0�J�@�����g����-��(�ee^!{*��6M�,D'o��$}�9�H�k��&:�ҹ^�qwt�Έ���_3	��}������p<Js�Z��l��-���N���x���F�#TT�?�^P�N�&[*�����!�#�i�1	���	͂H��� �W�ʑq_s��&$?܎3�\сR��n���A�$�����F%@t����ժ�Ѡ�%�I�r;����Tψ'y^'YV�26����Z8��ME�?�YhO�_�{�Y]*��cס���x���G@�ڰ�e��P�P+��	;�V.��ld�g?�ïӅEj:���{ܹ��mRAUokcn���,��G����W�CA4~J$������k�(�Q�q��!�F������/l�����{�-�E�v(�����Q�h��=�Z`�+��dm��uVؖ���>n�v���N�C���-`�ԡ����hY�{�&*W���E�����
Uҳ6-�h�Ǯ ���R�Ƒ���.�������aZ4��g��kH|J
�  =��R@�}̠�֡Y5Ö�C�#�)R��!�@UCd�	fL;x��%.�<�jۄA�7��]���Ŝ(b�ۙ��M~k!���IZ�I�fK����pF݈*�(	��0u)�M��������)�:,+�-�X�.P��;�CJZ9�q�G�yG�)b��O��][�W��J�"v���w
���}����vY��'ܓW�Q�5�oZ���Yٷs9�Y���&Z(���E���@��K���y4���l�����|�+6*��3D�P��!�t���F>�z�qL+�eJܱ�QAj_�	�b�<�(n���= S����m�#�3� �ף&�=���do)Ԡs��$�הŊyݣ���W[���W�.��Z%��i���n���"���}�b�z�WY�>����)�Q�?j�vw10Q�V�6��l�k��-u��⟍�S+mmwm�ؖ�E�0f���4�4�,�G�o���$�J�L+��"���:���<X�!�h��&��5���5WucA��m��Dg%3#Z�P~�iZ�72����]*�{똽r��OJ�s�)VTѬB�c��ӿ"0ݗ>��ޱɽ���"�ʬ���ќ�[00^~����|9s)��Զ��Ab���n�]`���F�����Y3D�c����F:��������/�����Hs欼�n�>4���VG��6���o��@e�8^N�\매�^z�Ԕ�3��uϱ�f��N�.��3f����|2vESY<�@;eU�V.|*�㰗�5d ��L8dy�RHܥ���1��Kk�"�d��1]���7q`0r��,w�� �u
w9�qK�(Ő�v�X��CǤ���A0G�O���c�ʈ	�`�;�����ȳ�&Y�8�R|ѩ0TC�w (pؓ��Ib�ɡߞ��90���������j����Mφ�w�@��5�����q/��O���<?�3�����%K���}� // ��<60P����g���#y`Ŷ]_L0��#m�$��G�������T@?��a|�O��g�;�T�gz݆)���R�գ�UdA��՟�8�d\���\���np(#dƐ��/�'�xq�]�����v��3��~{�og��2�V_�dDd��->��g�ţS�L�wy�ܕ����n|;��}��*c53����[��b<Y!S`���o��f�a'j��cIu%�1�|�Y��d�܄rB�}kc�B+
׋�z��z�m"���t
馌ͷG8�)ㆡ`tr����s��I0�_�"�_���l�8�\a��n�P8��"d���I@�p�뇾Yz���r#�"�}�# ��p�^�=�H�fk�@�;�������!���Ĺ{$����P=�[orؖʠ���!^,�����	4u9�E�1;Ņ<d���P>�@8�v�L�����9U!C��=���i&d7P��I���1	��� i�W�6��E��L�fդ&��G�vP�I�7j�Kqc!vu��Zk7kK���j�R�)�J��n�Y��u��	�ib��JG�i��{��2�f=��ۏ�~����ZW��>���n!�R��KC���ϰ*f�3DW*��=�����1o'�u�-����}�Z>�����a�Ŝ2�Z+��e�I�=�,�tfD��Fp�]�n�l܇~�j?j���o|	�ϖ"�fI��y�P(���ϼC}�}��>�r�-'ʡ�$Ye��4�4,��H�0᷈o��(F��8��S�R�$������gQ	'��z/��ޠ�HM� ����}T���=���g
R��Go'�Q���I�1�rmm �w4���"��閬s	��Z�c����dg��#F�̼�Լ@����Pw&Nb-~�#:ˤL��S\1�����F��7��9����K�t]2B��L�����+q�(��	��A	���3��e�B%��4\�x?�������S�n��	�2�qU�D>���Ti�\�ϵ��z�'�B"�%.d��3�$��)�z5آ����1����Ŝ0�ka\v�W�Hw�?&�
���T�{<}����IZ�&oڈҕ��t;5g�B<
�'G�*>1���3�{|�����0l�D�\�.��9?�<��u���8�1&����HAw�;�ǒ��G��(7�"(b�=pS�W�W0���'uſ-�P�v��T6`F�2~���q��؎�D�����E�5���<��5%���콚]e0�3�@����K:���!F>D>�p8���K�s}�A�U[�=���t��}y��c�~16��Քo�"m �ȍ\t��1t���y�f<�*B�-��!�_��'�#v4��Ho��%ɖ��4��T�b����a��B]�r�̫q4���7�{���h�6�����h�nI�FdU��/!�3��j�xl����S�:&ń��7y�c8�3�*��[��u�%�U ���&�#�?QK�|�'~�5��Z�L�ӯ�W���{�q?�]�Ŭ�'u�{��S9�[vʮ]@Fc55X&T{��0�i5fl+��z�s�e}��\�V�X�߿�hU��ክ�z,
��*`D���.�O>b���?J����;ys>���S�^�f�q��[V�Y��`�	���Z<�N�\R��~2^���@1C�~,Ю���s���/v��k���c������PH���y]y�4N�&I �3dd�:� ����8��ܧ���ӈC'^k��en��c�����g�T�����i�ͳp�雱� )"�!����Y����;	փ���� c��{U�y�K���"�q6ܸZ L���\\�x�
�#!�I��j/�hR�Q�U�!�AMvK��6�'�>��ɸ;lx"�E�`�_\�Ҥ\�A�*�j���j�����`=�E��_�QЭ���E���{���G>6�V�.u�����"�Iv|zK-c⛣�"��b1	�S����0�e��_P���A�����/����:"���{�e�8�X�Q�{��]^�s٘�&�S��l�b.��{��|O_)���q���b��\��V+-vF�7(7Y�� $�-�7����w�@Kt���]ɻ�j��H��7��(�5�S��������?ZCd�_���4�2���bS��F����Nx�ݳ��9�c��&�)�k����Vo��RJ�)��Ő@��[��y�g&Ψ��Cu6�S.��W�o�p�₂�xts���Zq:�3�^qJh�����zb�� Hߴ �:e�2��4�%�V���p����D���<��rn&�d�2	�|~K:���i�>��BRe`.�χ�M�g{��x �ȷ@�|Ē����q�d5�~��,H{!�u�
������s���3�{����Eh@���/��VR���u��,�����A�qn!פk����$C-�)�U`��C	w��:E��R(9���!�����L�U/�����KL��GVF�c�+f)x	�߫���E������Hg3ل�(�#s{nx_s(G�	�Srz��ʸ�H^E��gH�5n���_()�BS��UQ�ް$Nc���Ȕ��Z���SƆ�7^��;��.|��Ƅ��6��,� ��)ѻE�]&eN�)D|$��]Rfܪ+����8o尧�ܹSG��|��Vq��L<A	�jjXc֯�u��Փ(0��\���8�qMr�zưT�z�S���"��cWQ%��OigI��A[������Wb�m�l�	���!?<s%�6���W3��e3�>L�v�["�d�Â��~�@��r�������O?V(lGaQ�N-�����|�!x��$W ���<�謧&�M�'0c����,�	��.�.5�[6�޼�
�s�����F���r�e~�k�F��z��ا~�`f���u�X�6��jNa���qR�=�� &�b�����8��e�ѝ	�����xd#���e%M%}PQIh�'̟�/����@76T$I�,�ٍ�6��]�᪴��~�̑��T3�^�g�	o��$g$�,R.%���Ł9����"ŖҬ��./cu6�P�{��^=k�%��#f�-�45L5��EX��0iCC|�f\�F���'�EĽl0�]M�f�A��m�7��K��>��u��5h����"wDN���T�q.�$������)�3�Ut�8e7�!�b!���E!羭nF]�Ȅ/B���T��Y�I//H�=xeAE�8�O�}�D���w�w9��c�qB�۱�pcR]˺eTbv
�"8i.�w���IsMK}M]�������iݒs�q�t/�@z�̂;?آ~6�]x?P?r?l[�£�/�Q�X�<�ٕ/�HH��d�\���,.�䴞Ƭ����a�����운J��|6�j��=^n�o��j���c�b�� ��>S��L`Q"�$HI�w������4�'�0��f�$ߠ���� �$=Q�qٚ�v���97O
ry�`ֲ��ʵQl�?�ZKU ��z� f�iU0H�ĥ�~G�R]���ܟ$�ڣn�_�&|{"b�v��m�����Q̫��s*�	󦈢�� �$hQ�|�L;�p��F�p�HY3	_�0=8P�UǑ��
Kk��:�U鼉��o.��4E1j?�i�eL<K��kvaڈ���b��W2�A����*k�qyz_Яuݲv�����;��<d���.>�;�����+���bH�����<��q�2$e��E	�\R�9j�v�9(m�G	���L��������s�ߩo#SIJ�"��h����N��/�n�L�%i*���-�o7Nا�jꐘ3I����Z�y�c����Ze���j&>!���m~��Ū�͈�m+/��!��Og��v�r<pӻ�Ix&��q�p-+JuF)$�Q���Ӛ|����D%)H8.����-�B�r����A�S'+�h�"X�>^^���1�Y�q,?��{ .4l�/�M�������-?oKsDLyS��r�=��D��WZ˪(�I	4{%��>�[��;;rD{►��)}#�:�{΃ K��%2\x~�q?��E?ȫ2^��r��y?n��&��9REH�8�
��$�f��'�e$OYm�j��&$���7}���\��
1���dk���+�"�ۋ���D0��"���؎��Pfc�le�eg�f�kC��Z˻�*�j�ܘ��
.�/��i#:�>c^ puPي��YEPw�(�&`�Q��3��5��b'�+Em'˟����LN T()�g��wѮ��#\���,C��R���W���Ջ����R��nCJ$�!�o�&��!��$�*���H��A���ܥ'�����1����k����n�-�5#a!�A(�$���������m� �v�b�x���p螒���(�y�^Z-�����Q�P����9��BS�$)A�F�v-˜1ҳ]+fw�bQ�5$]z0���b<T�|u�а{-�|c�礪�:�xq��:��g�'��8��0�B]
�|ab��c�������s�y|���-�u�H��|�`��6�\�h�)��o�.V^���g��B
F� �%,x���L?�)pZ۩yAK��΅�w ��A�*f�Ca�X�W^���g��﷒�V]���&9��AN!*w򎜲�R���e'�[^g���Z?�fa:�|�	��}[j�魀������� <�|�A�E�9E2��(�)<�����;�(d�h��z�jlu��K�	��&����-�i,�k�přr#�D�;�l��JܤO�������W��C�.��h^C��d_�����L�r��Z1��us�J�G�)�����/�$�����H� t9=� �9|�n�A�E�O�0ϛ��$�ܒ<|����vj��a��A���Mp���(�`��&����~��de���g��^� �M#�~���sw�����/��3�}̯m�8?2Z8��x����j�r&�#i?_c$I~	1&���_�?` ��:%?��9/_�Q,ߦ�xDrJ�j�? �0�h��E���Y�V��>׆�Xo��ѵ�����:����o{5tU�~�8�O$�lY��rmL/�Ĭ��hW� <����#���{b�<Q/Aԡ��IN�ۓ?,�8pDd���B���A΅�MO�q)/��w�����p`�f@�Q�?ᲁ2S`ݗO g]�ME]�U�����q�}ڂQ_�������ZJ}��-4����@�D��HA�G�-��]��M�U\7B��@�w��^�V�5S��qcU8[s�͗臟:�QܪKR3҆Rc ڪ{�²T}� I�3����^��)F5~��h�%6�N���{����1�JI�4�U�,�������9�_��FY��4m�j� LPoV�/��P��2׆��b�/�$���l�&Qt��_��(Yٮy6?�p�{�"���XCZ|I�+��{���Y���k���ݏs|��y;�3vv���?3�� Øc*t�����v���e�D�_�ݞ8����	�|������2�M�.�
�u����t'�/��1�4��͏�`N�a��ɋ��� r�F�S�pT7$w�%:@e��X���r������4^�Q3�L������xɬu�	H��)|E������&�!�y�3\�����;�0	��� {�zT��C<�U�-X*�M�!~���Y��4z��~_X�NJ(��Z�!5K��1��ėc8���yf�L���y4 �Q~ۑ
�~b��^xM#�'�ݢ��b2�:2�LT�����;议�A�N�n�#֛ N
oC�@�C����P�ݹ�D��|�P4�'�ȆS ���U^�>59-�G���
�{K�b������$�?PL�Z��jsia�|I]�v�0�%�V��,0��&_h:"����Q�B�*�S�m^����>0Ş�=�/g�H�%��@3b*�O�Ώ���8j`>2�}����̛�]��]���⏄eW����%�]�	����˧�R�9�!���>n��֚C�sOd@��pX0���ߴgC;7����H�����˵�����0PN���+v�G Fu���n�na޽6��j�� bb��������8t�_��Ř�8&���S�i���nB�r� B:28��`fv�mh������]5��Bǖ(����u�l�����H�.�(G��9����ͻ�nwo{�n���(0ݮ�u��M������Y�݉\+��[c����	�A�pBQn�!��nSKB�Q��|̏֓��f�wT��k@���=�U�Åى�"����>���&�A���=�u~�'=��I��!\J�\�Eu
�gQ�Xx�w� 6�:M"��QTD1�`)Zq��xG�Iٵ!�$w[Έ���}
���J�=4���W+'�h�¤�W-J�]��E�M"����v��!B�" 2����OX�)9���D���=�� ֱ�I�}Oo8=��o@^���Nk�D�*�w���$Ţܺ���\�4��w�y��+g�����$�����w��ڛT�K8��6���PoE��ϨUsKX/%m�&�Mc�!D*���F1x�	�'��ܬXj��@���Y���s�]׭� g���Ke>�@��	K#���X��3�?G� �s`Gn@��Os�A�����^
�Vb���G �[���A�?}VA�����T�yi�&[igO8e�azҐ[�/yTa1�/�k���W�BdR2r�V R��4U*�rc��Ǫ^�hM����Y~8ڰf7uz�Vq��*%u�ӌh:�8,1�F��4�g��ܻ��6=�0,��ǁN6�w����z�8������N*�a	�*�4?�н	K�],f�(�c1s[^+,ҁ�xiO����D�g��3
��w�l/��'��h":e,���(��)��)�@��u�U���F��q�p"��b4�+x��z��ޫdC�E���,�x��!��W�U|6����4!��;���	�nK�k�D���eĨQ)�z.�����؀��c;"���{��Ux@ֻN����N6^e�D�*�_��8��%G��5��	~��1/J:�_�1�N��0VH��D��Z,i����{{�ݛ���Op�Ԟ4�l�d�dr3�4&�H���E���)����7ᆑ]��xn�̧�H��b\R��.�I��[��B������Ş���J�}���@/Z�l')h+��Fc�Ҁc�x��#��W�#�y�{Nq��T/v�����!��y�50@C/����0D:.!!@J�|�H��մx�������p���B���H����ȑ\S��4q��v�PG֗��&̼�!f@.0�`�pz�絭2���HUw������cv{������*s���H�&ԈU�(ɧn�ө����Z��|� Q'D��6%���r�tb��B��X�]�y0�q�s�劳��u+�a6w�P���	���ׇ���<>�bI5��&JB��Q��>���(�T55��X�y\Bv�@�$Y8]L&�ﺃj�/]�˹R���ȍ}?�ei���O��@ �_��Oڀ6΋�����qŬ�:��n�r�������L6����<�ϡ���Ka�<�w�{7�Z+�`��������f�畕W.���&O��9P�s��	)hZ'.3ِK������U���Z��I  �Be�G�> >��r?�Z޼GSR��Ur�ܾ���£q����+ $�,8��X���R&����'\�sr���v`4�l����`c`}s���l��������@^E	R;��M���wxq���P˰~�0��kQ{H�A?��p>f�6�j|z#�h��vCf1x�JUq��p�]q?�]+v��Ds��4�y)������0����K���B�M�'�#����D�GJ\S)6�m�D�8U(���"���4.���t�ɒ�L���g�O׊�8��h�dO�v֋����^R�?�Kw����ڵ;g>��z	��F�s�Y�Q��l\��u�v=��`!0�:�i/�u�<�h̕X�����re�o�x��Y�;�˙��|�O���������I���\�Y�����,���uZg2���g�&�����xԂ�N��8Y��)˙�c��dmÆ���l���8�v�f8�����I����u�����Vlg��M�I�p1�{��m�щF����.�b$�Y�J�s�H����5@�7?��S�k{��Sm-��l̓�1�2YƥOi�@�}0yγ#!��# �@�����a��� ��Aл7��eΞ��?YS�ya>8��	������]���X@!�^%T��&<�� ��H
��:��b5�����H�-�G��SsZ-Nzu�4�G�4N�-,D�`��Ǔ�d��g�#N�ߤ���G^6;�1FSA;!yR�����"R��b�H�>����F��q�-�Jn��Цք����K��	���h�{�Z�J�%�s�c�]���f�O�n� �bčqb3MS<<���O���1�:�ѦYV4���d�Y���LTӌ�c�Y$Yn�0�
��q�����>���'����cs�*���x�B�V�Ek����`q��{����/	���f��"��n��;��Y�hQ�����+nJ�9����ꦆ,f�j��P���3���y\�;خ�r������Lu:���N4F�r�\v��4R����H�b9��a�d�m�ػ5��}.t��m��V�v�aV�h�Ew�l+��ĳ"�n�g�@�P��Œ�.A�rxL6@�~I�2��pD$�Z��4����̔~�K�d��u���;mv���1Lq����-���X)p0Lx z4��{��V߽1R�JZ,ff�a.���l�@p��Aw�r��!���h@�a��<	�ʾ�B�����t6�} �C�2���k"W�+�5�y��AM(�G���V������OJ��h��9��k<p^�nr�N��C 11�J(�1E(ADƼ%gf}�� W�I��9F;�pJ�oL�ު�����~W�COIb�!�t��9�S�8ڼ�H��t�o����xBO�h�"�#��۹	�k��R���/	&���Z�|d����U�/z2Ɯx�������jG,);���	Ě��_#p�QL.���~�����;����=���UIb��p��N��=���~W�������.�k��\�x^��i{]\. }�����ζ��l��JFO�� 
�YͶo/G�l꧟h��\�לp-� �y:$[Jz0Yoj���IH�[�u3���=}�S�1C*�<�z?��9f��	16ǰ�@(9>G�<��tUT`�Aw�[,b1�>�x�.��΀2] �R��l�G��l�={= �.f&)W,�yT���,魢�(�v<�}N�8}��%Tկg��q�o�]���*V.��}֫�,��-��U�y�8!�!(]�76z�c�]�(�HYW����fY�p�f�a:)ST�RiE�~����c~r��3��\h7F��d��!�9pU��p}�Z.=@��ʩap��s5��$]p�8�+"���z>..'�7����?��L��S�v���`��ͽ����o����S��=�0�d�/���hн ��z�����g�W_���^�3 ��dJ]��h�ɢ�O��"�6H�]�ґ�DUP��뺳.�3����N�.	�����͜ �Q�9v8��!�Q���nP�����d���1�Wo�������4ݼ�M�Փ�t�e�A&�粮��� Yޤ(`���Q�s��(���4�k�����yg@1�Q̯�w���$y�����\����\�}�k�Y�������5��ȷ?.�ӑ�3�����:~�Q�'��f4�]�q>Lq%��k	 �JMHk0����v�g�@��59�z��i(!�@�~�P.Ɍ�$�%����a?Db��8�q��O"�Z����y�L����G��f��˝jQ��=�V��>;v�ͩ���t��H��cS��O�TMɬ���]�1N���2ty��5P}_��AF> Y�fD�H1��D?�/��<]�NS_�k���y�iվW!aV"�3��ҍa�9�\"��jU��*��ݓ��۔������{u�+/�
��s��G���}�SΎL�H
�3F<����u-�Vn:֢�q3[e!�|��|�0r�U���a�;��U;��Au�4Qɨ�����a(e��`��鮭̋kж-�^7B55@@\�n�� "G��z��Ez%��LCCcF_�9vz�E��5ǔ��)�]�����m�$�v�m<�C���L�����]G�(j6�pQ���Ŋo��{�a����S��᭵��߾څ[js����I��@��`��_+]�J�]�N��9z��G�O��(��wB}��c-h�ڤ����xkQv0p�	Oi/����]J���'�F������ٝ��j2,�H �;1/&���X�!��}px�ע&J bAKpN���7���QN?�E/�ue��xb̋]O;M����iէk4�]O��
��q⦡a����X�*��܇��B�q���������A�>kt��ve�Ի��t)���;F�r�п�r�$'��L@}KD�V�W���"��Q�}!2��I-)��}�l�����wY#hT[�c��z
�Y{P�����J�!s�d�z�M��/Pe�4as2��1�����%k�#�ZU��s�����O#��n�/no���2-��ҷ���$��E蝩Lo���_R��gڅ5</��{֟���M鲉��|�(�a���L�fV�<��v����e��PY����l�[�ma�yj�,��Y 4>Q�AӕQ�Z�o�R�$\g;�#��L��{���)�g/G�3�s<�����Y���m�-b{q�{7�!*�;�eA�� Aa�)����*�)�6:He������^�ڭ�$'�D�)+"��2�g�Oc��02و���oadΕ� хy�&̮���U���� ����&��@�!+�U@x�k�O����,�2�-��/��*�M5C PJd-@	��7Z�B�OZwz�T2�3?a�(R�<*З���)���ܐ��Jta-	J��ҕZ7<\SJ\�C�Ъu��g�����������PJ���0��E%-���0�*�7o�� 6�>I�;q=��A��QMXw�.�ț�UnH�;g�l�DS�=�h�p�Gdod�;��N'���1�����uU�$0��:D
gF�K5�a�$�X7��B�4c�M|s6E��9,�������v�N�h֜qI��'���L2��,�E�q�g���>H���6L�K7�;P���Vd����6�y"<����%�0���3U�+�h_H͇H�{ �G8W���G��t��i�҂��e8PFg2�)M+��:Ж���{!�u^��i�'W=m'���J�0ZD�gH���К��rM��4�S�����,@1/X:����1M<���`7������,P,�-�M��(���;(ղ0J�z��$>C=8ys�/�s��C���:���S\g��Q�)�K��k�;�KHމ��Y���� �x܃��o1aQ������y~�WN)��`��i�-
��3����L+N��[js/Tj�V��!�dL��Bo L*��U���l�/>��&v�L
��`*��?��f����8�`���oZ᐀�d���N���L��q���|����h�FX�ݱ8����2��$��u�Hd�*���e��;�I0Qr�ch�y.KW�y���B�b�� B�qɫ�j���6�"�"V�y��뒾��6�}�I�F�k���"�"E� n�B珶)��-����!Kih�}	�-G�M>��ױ��O���2����jׁ��Uf��{��nw��n�u�^�Dm�3!*�(y�o�8��T�o��tA�s�@lb�"�1e��X�W�`��&	N���­�g]���S�3#��::�*e��T|���I��P�A:sl�:xȼH,�/�<O.�v��ߴeݷ���KK�Zu�'*j���f�Ek.Y�~:	��5ٶ,�N_�.	��.��"6�:�7i��<�R�1	����X@:��fz�(`3���z���R+�E{���)l5�vr��l�H�3���wT����t�!�m���+����_Omz?!$K%���RG�1�,��k*�?^S�Эf���!�	�|�B]�?R^� �:h���̒a�ȣ�u�w�k�AXb�<�~���Ф�aߛ5��>�eE�;׸V���c�W2�Y�X~��ɭ�Z4ǴJ��v1b���Y)�b�8X�/���)j
7D7�UA�A�UcK�����O�SX��S+:��!-�5����"�FG+E��H�����Ӡ�~j?`1%{�*F��^2�.�L�(����"G�`W�ph����S���l��@�V!��Ty�H�+xFl��zo���h
�7W�p��#��vL�����.�v�͙c��^�C� '��4�7�'�MK;�H�j3�~ (������|��Z%!��S���kX���Rh	
s�}�sA�Mk�] $�i���7y��@lG����Uo�J�x�9�z2���j��(C��6�I�Kt�����04�E=��	]OC��D�̇$Ht2�?KVV3 &������J��/R��>?�ffv
�H�v1�[m0�&G�D���>��鄎xG��'y�'�,��6��E:W^1B5A��hv�F��s�c����?.�į��D�;w��"IGl��"㚶�=��8�5�w��k��_mҚ��"�?��dSt2s�\�8�TF���esz��%�,R�3�[ܣ|�IU#Fٳ���!\��@���t�b3őkh�:P�t
0�/J?Y��zv�Ý�3�� ��k��pz:�������?9s�xg����S�U����Eh����B��Q�{��z����L�����N�nFNB��4�C�W���ϓ
ڲw�B�sk��~y���]�,r7g⠾;a���.�-��V�����=Y��/��/�Z`� %Z^��⡍��bA�˗�Xl��D��U��-Y��<1';1��a��)J�N���hΉ�7�FiR���ة&֎���P��CX5��8��ٟ�Bn-�����F_��P+���8��m �lH*�
\����R��H��!|LU�~�� ����Q}�BR�G?t@���Zpc�h�7�O���c�_�ul�4�V	� ��?t�Q�_�[�=�_�BP<ZR�ՇŸ]���-��Ӻ��$$�# M��O�Y߁��n�G���~��{����1\Y�"\�� @��nG����\E�zQ'�����#D�d��f���ҝ*h���Q;�N���9>�?��3��������-�t,h+�|�N��gO�#Teݽ�Q��L~\��q����1�:�����&��r։"ƧUh�����e8���?M�=�u
Z=��&�Rs�,�1&�:��]��M,	��cR�������O��c/�K�ҫ���,
�vɿ#���y�ВR���MB��	+y�ܩQ�ŀި��-}S3CWJ�)�5�90���T���ۻ���-��6C�0�qq����� ��e�8�b�Ӄm"v8&[QB�#.U�U�I��)9	?�&���d!�>Io�Ě|a� p�/�z��%�<eh�U����zi�-�V��C�� +?���5�C�4��(>^�IgǨ����P���|>�G���i�ؑN��1�.�\>i#��~�8��"�R�Z/���# p���b������"A?�$�������h�E
�܉�� ޮp�����AM����!df�}�j`����D�H�GU���
�������� ���̓4+�����T���o
�����y'��j7~���˷��s�Hd�I�)aJ'�� �Ɖq�!�9��n��c��b�4�9����7�"�P�=�D���� ��`���h�<Q^L��&�[�e2��`/��oz)�ŢN�PzVL�2���}p727�.�{�xd=,�3F��wF0м�`k���'(%b\HJ��Ң�̪<|4ڰ�"ҙ���qA�sH�W	�*=̈�������E��j���mt]�F.x1��;!�m���$��?�	��e����h%��]�Ğ>բsf	��U�?w���	c�e+&,?��)6����y���Զɬ2Q	�#&���P�鍠-\l��x��D�pB ��T��4Ђ�۲��	�BB�f���s1+E�@� �ƀc�J���c*�%O�K�'�K�䝪�����je�<y"�o3�Tr1����+F�Z'į�u�sY���W��0I�% z��n�"dj���PUs���T(����pgH3�wۑώ7���7=�PK#��ݶ����5i�ȧ����ף �����g���E�^l��}L�[��1��zsS/O��q)E0"`�\��;5�}(-�tѶ��dfӶ�!\�#�&!��4�fT��#�)"P{��4G��9p������jW�#�'��9�-�~�ᕉ��*:=����Cdd>v���wM��n��H�O�k��+�QG	�vx,��4�g(?�0,��r'��������|�9)��2n����f�t�i������߭,����ГB|�����p�J�-�m�״&)S6�l��@�0�ҳ�V��i%��@ס#^�==ǚJA�z�6��� <���.z�Q��YCln+.A�6� �K����)O1CT�T��.K�(��l<���p���]9�r:8��!8(a� ��4��F��Ϻǎ�xA�0L��ߟ@�|9�{�,��4������@.���dR۷�YDAy](eqUEw!��{˕�o�V�"�t��hR��mY6�1���������9��q=��;VN�Dl�%/WiT:�}Mh��u�]z=���rܯ��7-��`X3q3�m�W�/���!HWť�m=���~���M��?���p�7zӒ���i���De��+���9I�k��ZHFqJ������0XY�,�Ź�&��<s[����L?D��j_��*"I���M|�����Ou��.����Rs�����>���r�@7���n1�2#�$��*]\�����4����q�
4�|�1����'�m�R�u�-`z!#S�����tm�X�nI�@q���%r�!�9���Xv����i���,4N����l��;	Mf	�Q�s�]�AC~������aH�kZ٩u����'�q۱�m��e?�^%IL��LF~b݁w���҇\��j�!R��_Y7�.{�h�������/=�E����9���F�/�W��J���؂�IΤ�?G���
j3@��{>]�>74�l���(4:qν"������UC��)�C�}=슰u\%]_h�_n�w�P�G�!'���*���ƭ �:~̦z��BM<����������ԙ����eYe0Iǯ��n�#߬��;�^a�U~��_Z�RR�B��,R=�9�y�EB.���WI�]�Xgs��&��"x�E*C"?X� Cɫ���U�ܞ��H�4%�� QAS�$���}��3ۄ�Zt���y@7�	h��S��#�౰���*E,]q�,��Fg�k�(�<0.���	Q�_���C��(g�Hs��`�c���:��d�\����C|D7#B�Wdn�7�1C����k%�D��������O����y��!�:��9�ڽ\�p��{���dN��x�j-ׁ5���{�a�q�yJz�	��(�f�㠇[e�
�>.4M��� Y�:��ߚv����u�߇v�?�VʵGFV�6�KZ���[N0L��J�~t���X�K���($�N�:h%х�~_b��bD�l�t�.u������A�
]�=˶׎}���Q}�^J�ᄺ����d|2QR�x������?�$~�T���ܲ�;nz��C����u-@ke�SS�p�$�Z�,UnC�7�.e�
,�$�V��D/F�+��+ds�>��#��F��,)M��J��=Y��v�*B����u��&��� FT�%����j
Lb�^ ���4�1.��B��J���Q���XX�����t����è~�ryAH�9�ɯ�ľC�<�����4t�|g�U����?X����*����Z�;d���n�6C�( |d)@5/e�Ñ�]ZVu�T���W��:^7~�����4�h�a-,�W�TȒ0���4���TnA��CE���/������2�Rl��(S��-#�Ìw_�S^Z��G�!d=�O�����E��D�$��D�	���{��� $VcJ|`����� ���)���S)��i����EM��H��
wu�6�܅�^t�D�&4����R���5�93	}q�Mr8w�:�U;Ծ ����L��z���9��]�$���^�G������E�OX�`"C�!�� ��Tnȣ �]��V���L_�,����3|�	�o�.�0(d�Q_�&�G���Ѻ�R;�����KW����8���ʧi�"!- �,ϣG2ߝ<!#bKr-~5�)�Iq�4M��д�Qġ"P�w��7ْ̖��0��ٽz` q��CFM	�Ś�'M��I0�P`��/$�E~�tV�Q�c������^��0@�B�%�o�r'���P��6ٺ�����cl��#��l��^o�'m�d�Rc��H��2�JA�����9�@�ͶRR#~�;��g��i���1t�M~[1{��,�{+�l�Ɯ
�V�H�y���V���P�����ώj��ڄ�ey��ϼ)�5�t�)z�_7�/����c_��9Q�մ���-:��)���s�@�8|>�T�m&�)�]։����"G3�Ed���'���Hf;�����ٝ{D}�,٫�`8ӞN #Y;��x���k+�\��,!k1����b�s��8T��=��|w��T�U�W�>/��%�`
)�yA.9W�k�w;�,U״�)m6��F�
��u��zC�߲/b�@�LHS|��;ΘFr��n�H�����z��dT�bB����M�xf_��'��n6��%= i
Qfk���ND1� �8U mJ���N2�cKv��T&��$�y�@��0r��w]�2b���>�^�I������?�{����u�i��z�b��D�ͽ�|��5�����"�?����d}�K.TT�[A
c�_�`��vl��7E^�Ƽ������6��!����t�/U���\w�W:7M��y}��Нͻ:g�X,�Z0׾��/��B�a�1^�8Wy�������Z�1����w,��[=�+J.| �~���}+8:R-�h���:kj�+�M�_�Ќm��B���q����#�p�=Ǡ-���M�x`_���'`�<d���{�s�q�  #eROip�t���������nk�� ��r'8|�O��y;4����Kћ7�)�\��8=�^��Y�-�\�P��'^�u��D�A�����  �����d�^a�
j:D��E,9[^�����]�C��mV���M,���u1^dUH��_�<d@I�aܙNr��'qk�����|N�	��?$<(�'+��+>��]������'�గ5e�c�FK=R�/��ؘ0Q����K(�������G��k�q�C9��w��swl�����&�CKb��옔/oǹx�녡�x�(7���Fe�8��	�[�gH�(�=ey��ɢ�-89c�[��}�S9��h^9f���W��^�ky���|�ZT?[��>�M̪"�iYHJ]�A���9H�����K��7���>��"�*w�7?_dA%b��4�J���UuFK:X?�8����g��&��T�`-U�|0At���\$�_set�P�фV*.���vW}��l���C��M��u��g.�	��.���������(R�=@�Z� +�
�??�|ipc��8�@PB�Y�al��;�F"��g��xg"�ʽ�*-ΚGX�����$t�Ź�	�F��QG<�V�����Щp�BY��U�Fg`GG�p0Hfm���E��MT�~���I,�rb �!W�s�J"`��ߏ��%�a=�pJY�NܳJ��70�]�롟l��QcU+�E���.���2;�� K�T,�j��cBQ?Z�`SdGʞ�&�ȇ(mr|)����mz'�S���Eͽ��j���2%�I�<�E�^�#e�a���1a�R��22�i35��*��R� ������
��TiF��o�F�o�"}�^DƸ+�,��;C�Q���+�M��AV3��CƜ�i㕛
�l�����J�Yk$�c/�i��t!�u�$;AO'��������(#���xZ�k����_��tk���Q$-)D@1�{cz�ª����ذۼXnq8���Ȳ1C�ٚ����(R�X^��N
�i,5R}ȟ��sp�m��P���rFzJ������R�K�̟�E����S��_�B������K�.,�<` M&q�/�ŊG�Y]<�W /�5�)���L��hy�L:�^[�o�8Bؒ�=JSn�7���9�.��(���1�\%���
=�Ǧ	є`"�V��|�L�*X����ca8;�X�~0��x�,mҵ-�s�p��t5���n1j1�v=�%)}�5�Řm��u�Ǐr�jII[���db�M�s���֞ș�
��g��#�Z�v(�~�pү��,WyO��BbF?ƽ���n4��zY9�0���}0fU��C_��)�|��lq�]J�RgK	�Cy^�Njk��id���m�C���*�6N��u��Օ3�I�l׵�+�Q>�	���ŀi��YReN8�T��-������ݦ��!���e:Ah���VՇI�{�I�ooWݴ� &�kJ�cY~��ّ�����qh�b$���N5VG��W`K��������$��u��9�s�;,6������`�_J�"s $4�,Ŏ�P���鹫���\<D�\w��G��ϼ32�m~���U����X�u�G>0������B��Qpn�b���'��UĀE#�OCj�� 1�0�}��s���bK����`�iQ��Y�D"Y�M<���lf�+aN S�Rݝ�#����--�@6���$�v�%�~�1�f��IF�J]-���6��;��39���M�}�C��B�ӛ��)�϶J���G;w��ST�����h�4�]�Շ/EO�lj��Ѕd՛�N9�o4%�9��",0u�aX�S�ʰO��e�T�m�"^\z�t�A��#j��Ng�q��K��-Y���ʜ�<�X Rl��T,��iS�x�:�Q�J�c/!cm��ܩD��(���ܜ-uB2w��W�&�&�Uq���!7?$��eЛ0���)�r!�x𡬫h�ld(��t�b���4��]>=4�Iא���T��~Q y<'D �M�r��oti�����tI��V-ʉw�����?��8���!~����6U��VZs\���T��5,�k�(a�����5,���N>�����C�^ W*��aclFvI�q�A��ћ����]܋#��|tc5$3������m6c���Ҝ�nx>}<����(̹P�	��\�؝ɵ��t��D=���Vp$��"��\m�������F(o�_:�@��)��Y�P�
D5�.���0ԶU��IyKtgj��2<�)w�����g��j����Y��/�'d�)d<�2�|_
̲"��2�6c��Ҽ���V<?�6n�s�˝P�$��⪻��:�@H��m����B=����Skl�ϳ�y��d��9��c�l�����/ݯ£DD��gy���(3�X��A��zee�+��S$;����Iduڻ�j$���;�&�a���
z��Y"�%b�z4��q��J�G!o�|��Ii�+#��ѐ�ڧ�����R�'�\��b���(|/��:��6�a�R �Jd�O��,�o:eԳ���<v��z^Z��9��Bތ
�־UwA�N#�Mx<��m��f o�©є� �1��v:��������Mf�v�%J�Q�1���Y��P�481�.0�(o�ҵ�.J#�R�L��xb䕱�ۋ_���{��{@��q6�3�cR!���h4zo:���xQ�HR_v�؟�����ؗ죕HX��C�e2�/��e�R���A�� 2jc
�f�@�I�5D���f)�ޮ��;�g�OG�xm�h����Ƥ#S�u�4���B�l �!��SUA�"���OZI�Q�ۥ���MY�5}j��Ѫ'h���ffZB++�d��{�X�Ya$�jٶ:ɧ����,=����na)���:,�Y�8�u^P2���3��������(I���_�w�(��Y�}g{H���z�j���sg�\<m���j8ré`�-�eD�qRR�)�������Xb�0� �Ի�} >�W1�R�r{�3#/�l��F�ϋ���kϱ�����/:kWE�^{��`���t��^�\�&U�5�Q�V��5��T�n{�����5�!%�Y 15[V�!��3J�R�3��9�Wm���lg���%At?�{���A�G	��;� Q:��,'�"�UL�h���)y�JeTH]'��Dե���L _��P�Gm��DI�w]ݪf�h
>�F\�nE������%b�����2
)\�����E�ٻ��,�>i^Hc\��\=u�{�ʳ
J���y��m=�[��B�Gs%|��������OW���%
�q�d!2b�s�@��F9��_�z�
^g�w*�"/��Ok,[�V/Q �M�",��0�y��ّ��<�A���U�j���ٻ�X� q8����٦*�S0J��Ư�~x�|�է�� >��MM��d�Q�d�Wx���� ?�kːcY�NiN��|�:G�'�,�0�=���u��nI���:��@72����:0�1�N>��F��)+g�N�!�f�����������X���~�ԯ�����$)�] �w*t��406N�^��pe'1����� ��kgr2 ?.����PE�w�gء��z�L?�6�"M2�l�>b��\�}�:��[������2��V�a!/�z����o7x�0�����cR���7a���sИ ���9��OV�g�a�:�I�\�%;vVjz3fhf� �Ok�!!j�ʌN�c�tv���Z9W�$��l�Á,�9�XA����y���+�S��%����j�+��� ���`�q�Dߟ�]9,<Ԗ?�ܿ��Āe�,�&e��b�}l�n� A������T�m�����U۟d��H����J/��SS�ן��e)���=��$�q��:��8�ͮE	��[L/��
*�2_�������׍�<�¢�u�Ki��w��"���#�fr^X4!H��\���R�k79R8y9
P>��Y�1o/�
��:�%1��/X)�`ԨE��X�F�#���{-���=��R���~n��M����4: X�+�a2���2�a|���/��Z�^i�ST�m�N������3zK�����������K�شJ�6�8vX����_ituK�8���F@��e8�B�w��"˨���.���γ�R6s�ԭ�p�l%��:�p��GvRʱ����c<���g�w=c�Y�)o��"��Ey�h�j�H�1a���ڨ�+EM�5@���~����P[K���j�WX9��e���C�:��b��]��\�� x��������X�����{&m��$KW�|/���S@�|U��g?���%�a�A�?�Tc���;�e�n���#�.[鸀����W�ߙ"X�'v?]bz�~S\!�Yr��^E����^�#�{���#Q�ƕ���I��ށb��NVq9m=���j
�PG	������k���Q����D�N��͖��͡�c�=#���KaU`JP-�K�)��K��T�`S:`�;M�q���ܫ��9:�n����V��uu����g�0dp�˕��]�a���͆zͼ�c[W���r�E��A�H~�`�*.�рK)
�c���hDܶ���`���DhK�Jړɱ�����@�T���+1(���۵��X��[�d�eΦ�n̂q�<�]w�F!J*��]u�7`7����	h=u�R�YqG~����T�Ƃ�q�@�q�L��Wj��US���a����m~��8y��Qw���r�ff�v	m$��d�$�L�I�̟S:��餮hh�M6���J��g��C�o�o��X��xcxu(�Ÿ9���l�Jm
km�FN�7�t]"���Y��p$6B �ً�a��=���X�w}4�ߑ�gf4�!���FBQ09�`�-��q�a2��R��U�Nl��ҍҳtk&�@����0��$	��Z��r�����,0�ã�8p�Q�pή���KDZ�i�$QmS`�:6��0ǴUT�$���{Ξ��{I�L�~��ˈ�c�I3z��)x��*&PN��c�[-s��`�"���$S��w�=g�]o ��A~XU}5��t��2�3�2h@������V20��?�s�o[����s�Wpz�~0��pѩ���1��	�~x�|(��9���X:�z��OH+��Ӈe�<���L�K��������ؘ&Nur�(���+󵋼�X�3&����?'��J	����?=ϗ�/��4o=�+c�LW�D�� ۵��ӻ#-�mu�q�c�S�����&���+�f�	�����I�ݤ�0�-�!s�t���98*Ы��>��w�Zi�T׹�x@k�������V�c]�0Q=|yu9�l}��=Юa�Cvfo܀����B>��L]�>���f���P�-��D���@W�����uk�60)�N��,�l�
�Z>�$���t�e]�o���7�cb�0n�Zč�nV�p�iW��0�l>��Q��6N����È:ׯ�'�!Sxv);�Ԛ�X�D�U
����b@˘��8�Co
����E������F���W��͵�	�<�T�.P��<��q{���j[�d�2�x���
�q����v���K\�D<�C:������� ��t�	��մ�ܑ�́<}�l4ݐ{
�nep�>�����?(W�o�6*��U��aQ����^-�$K?�\��fA�^$S�y�d��̅�l��g�I�\�C$ݟ���&�F>�PATW�+=��6�����L�:����Rw���IAOG��^i��&DEt�'nt�u�t�M�&��) �;1"�B��Qk�č���8��<	|0���L\�S}U����ĻC���鋕2� ��2�a�\,,bd��8:�;rO첛<��b�ʊX���N�#��!� G���0��&Y'��G��5�j�Y�k����X��#��-�R��Z��zW�4�k�A��4,��[�'���GҌ�D"M��X����:keW}w��9?�Ƭ8�)��a?|.��������.�$�?�8����̈́���,Zں����5��xI?�'�[��PE�Z�惫��;36�M�(US�|�X@�/�u�q�ܟ�tU��:1�%�g��'�B�a�" 0]�{�� ���v�l��� �W���oDL�9�|2g׼E3(3�3�~!���˼h��?laYZ����ȡǜ���za�����e�&�"a��9��`8܅�0����-�CN��/�*+|>��jB󼢲���y�3%��b��0ì@��C��R�蜝����X}�=?1�ֳ��<����̈́�+�-�����*�8Y�G�KL���{�IR]��$�w]31A��\��O��*���Iu!p��V��I�g��3nC��X�cO2���-VJ=8�w�;Y�]�e����}�%z�����e�r�����y�}���nL��*���?y�&75U��ЫE��$2f��Q��w9Xy}�Gx5S�YA��0>Vc_�ěR=�Z�a����_�H�� q��)u��=?��q@�� ֊L�2�6����<�
�^��R�o�[Ζud��F�+�T7�.�ۆ�T^[s��7yq�-8�v���F_'�S{��
�"�"���ߍ.p��"(D'�k�#q�]�0b���wuhu@>��d�:ܹ'h�;K�Ix��G��6�gI�Rqz깓�HUe������&�_z���h��߃�b����)�qQ$T6N�=��&4����5�oʟ���&N���8��]Y_�ٕXb�Pg<g��G?�4}����!.#[����� �̴��k��Yw��6)�mp�3b.�D�5�Y�gڌ�/�=2�U�B0R�.X�pǃޮ���!)[��:=M@9)Z���R����?,b�@\=�Գ2r]�{����!jk�Q%�?�ڄ7U(�	�9 f���Tq��|ȶ������[��Q�q˿/�P_�>0"hR�.�����N����1�k$�yY7�6�>P�NA�����`�p�O-�{���d`2�	Ì�Uԩ6;y�E�zJ�.n2}�^{��[�˽��D �`�6�����q���LgA��>�HQ�ԙ��U����}z+[�^�Rg�å����q���c����VI��(Q�a�~.���"}-�:3����|�!#=EGG|���Sy�c6ߪ]���(7�W��I��#�݈�tR�������D�*#i�T�B��A�,�A)X�ޠ]�*g(�;�0Ϋ���;d�J�@`��t
S�OP��߽�7B�;˽O!�/�U��Β�w/�i<�� �䏍�J�������(=��^o��'�Gn�����I�-܄�'�%we(|V}�be�((�ɂ]E��+�m_S�o�*��F�h+�R��iݜ�
����|�ՔH�#��Ū�Rx���LϾ ��I> {m�h.fZF;��d���M� �},0m�GY<��_f^�-���ձ<>��"�$��
�x!�Ǯ�3���9��/�y*`G�*��^ϡ!s�қ3�xP��+E
��L���˂c{S?C�9�=v�ύ�r�r�P	�7��Ȁ��ae�����g�7��n�=u_b$�C�،�,ʺ��$���q�
�h�=���z�.ƿ
6:��.X�s�H�.la��F������~d�0�MA����*�����|�bTK�L'�$%�	S��s�ݞ����"��S��8#�����); Es�/�]B����]��h2���_W�k'�_.����
�b:EY�FM�o�\	-Q�=n9Z�q���A��b������w�����Z �n���D�Ε�%ru�׷�#�K�]�b�W��ؠ��l��S����9��+.������3�B�9���xTuK��5�p��`���eB3Y�7P|Į��/=�(�sxJ�.P,�
t�Am������'�����ۑd�������,@ڊ{n'�SJ���s�N��t-����� �%��&5d���& .��N��R�͍j�t8�$�<���mT�\z���]Eh��Kfp:qui��=��r�Ü�jz�Zj�8�*d03�H��4[���.��2 �w:ɐ�,�O|߂ﰣ�s�g����]������E��y�Z�ۼA��Iv�ol�ːq�T���ĸ���eC5�}�D[�h��n�v:E|f�N�i���p�A�	*��MD�-�4Dk�fh����\���*E+$�|�n
Y.�;PG��Z$�Ⱦ�����2�s~b
`�Jz�s�*dh�$��`��O��P��#<��,��uW޸����k؀
�/�:���?y��� g,�tϲ�m�5�ũ�T���ݿnlXj��c��`��|R�����X_gP�ck���F��Kr�	ΥX������5���y�;�<s>�	Ԛ۽ ��$_3��?ڐN.�/)��$MKR�;��Y�B�$����	:7.[P�I{O��D�����f�!����쁑ub��5A�w9�W��"���H�D�c���Y�ٷ){d*ۏk�w�_��V��heK��ң��P�Axl��Ӌ[�?�r�<��߀`��⯻[��m���.������Q�=1�LE`9a찃�E_���o3g�&�kSg�������lB��P�zX2�Y������KJ��d*��ےѾC��è5��@���/LK}a8�m��G��a$B�]q�p���m�rb ���{��!�b��:5CA����@��v�= b�(��T���:&����n�[�"�e��af�k>pp�t_�Z U�BÐ�%A��A�@>�1_L�]�oU� >4ZoҶs"�ٟ�'e�>m��'T��ZI�G��Q^���o�kǱy�3[�2��FFy��!O���J���'�v�ﲖ�I~�A2�s�/�O��jy`����ZyФ�U�Թ���2{���m�����w�}����Yd��G�oQ۟�ˆ���s��S��6i����%��� 8[-���(�TISyq�;Ҍ�F�*��;7�5�c����O�C�3��滤��O��u�!7����Up��"!�T���ܯv�o��A1L��=����V��a'�*4ʒ�Efޣ��R�����,x�IG���dH��j������sŶ5������[��x�7��'�^@}���s��'���u�vl�xf}j��l[������8��r���5Z݆����D���#"߰��V��%ɪ�������M[]m8x�'E�
f&/E�y	L.��}ʗ�</�4AOQ�惔4����B��Ƌ�q�]�_6���j[ɥ�D� g[�>\��0�� x�B{I���}��o04��^�t�Y �$����8�V�</H�T�s��Ţp��]�m~������+2���BH���_l���/�����Hu�.7�*����۳ME@d:[���x��v,�g>����p���c��,/aD�V�TCٲ�㟬�H#G���2b?"�5$Ƀf`��������4�LV����ިK���Q��}�*�i�����3إ�@p����Q<�����7�R���?�>z���@��?���H�X�E���H�8ɢ�wM���ڑ+�!��� #y/��ӻ�c�W�1��w��D���R�
vv��6`c��Kb4�`�s :�_��~*�"H��ǂ�[+�^�'��Hȉ�r|"��\�U�O�s����	L4�c�ϯ��ox�5��s�4��&�I]�j���:&f�H%��a��Ѻ�Л��=��q�2\��h����Hf���`�lO�6�U��������RE՚^G�f��5�����1O�v@����	'���|+h���Oy��G�c�]��R��px<u@*'dX���/퉶���ZV�N�@.u�u��H�k
��1ˊ����h��"��c�q�ׇ�<��@G�Mu0��8��Au��纋^��懳G���w7���Ԛҙ��D0EƘB�[M�D�Aߺ����G�� ��P�j�M�9���:�����m�x��\����x3T&�˷���-�*��%�����/����'�X�_�>l	mf����~\�'�*���A��Ig�	(�3Y�TAS�0Y�
�-�j�/`SLC��c\m"U�M@Eq�7�>_��褎�◯Q2��a��~�˷(0����}D(���d)w�9��t�������%�Ӊ���q_�)��rqCW�*>�����MQ���GY��wԼY��rG�ܽ�iX��
Q0�b��A�W�5�����!��'��������`�ZrH�,ăk�4���.�֒1��p3��^!�J��\�e*��7�_^˸�Gř��x>C:(*�nZ!��2�������(l������򙼄�!�%�|��r����U�P���h����[t��հ�L�JkF�,���1唆���ֈDFL{��"z k �J.d���8OL`��UGp���H�둚X�3�+Vr�)t �R$����!������W��Lr4h��L�l����0�v��Zo-����j��s�}���!�3���6u����֮+}��G�iS¹��}����"�(xt���zE����_���ע��!�Bk?�ڴ�M��e� �]�8)�/�VW����<����\9נ}a��ǡe���̱�-u���	nڟ�*'�W�ܢ��(��W����L8V�t�r�X���௝��>�2<(�����UߊR�.������� e��;�k.Y���A(}�������n��C��A�'�~}Āֻͦс�0�4w�9[��{�l��&��)��	��St���;6Iw�R�$���J�2Y��E��jJ�&ח�Ag��mF-��Sk[�R)��^S�:p��_Pl;59~��k�)��LP|�ezS�7�)��_b]m��OSX��"��zL!�K-[g�i�����/Z/���{3�h�t�J|�Я6��F&�[���y=킞-�fީ�<;�v�O<���K�-�x}8��2i�M���Je�Ng���{R�r��[3���T�0r9Xó��D]�6I�Wu4���ᕲ�z/z=��+�+́,������d�[B;�ΤN��P~�	�>Ix���y�Ҳ�}N*�|�֬��ӡ` 2�� y��+�6b씯�vR��7g;�wh�K��1�&�2���I������MR����: >��Y�e�zp���i����%�QK!�[�g�%S"
��ԃI�P���n6�Zh�Q�oL�������\:������ѪQ����>��:�\p��UXz8�7��> �����)�ٟ����$�έb��&2���Og�!et9|ba�|�;�'���������
��A`�mjuSI�^
���A쑭��������y�K�>2�Ĩ�L4�4ݣ��L{���N��1���~.J�];�#sN��g>�����P��1�G����~��FqA	I��?LCK��
Y��Xi����9�=��H��ɀ���3�
�Q�1%�c�T�=�)�`�����Û����b�}$��M۷��P���m�%ܗ�YY�6�G��ـQ��6ˑ����������|��\P��f;S,�4�"�� �86瞂�0,eLW�l+a)"v��N��"`N��s�n#)����[W��p�z )�T�6wSʃ_�g���jGT��7�U#Ɗۥ;2���A¶����>(�7!�l��(�E ��Y�#�-��a� �i>o�Dg��6��cg�R#o���(�A9.�
 h뱑1pK��t�6*^jN�E���1|Zw��cOz'�ɲ[��E)5V�[��
P�E4��p8~�g�4�f�C�Fi���� w�%S�!���K���w��?@���7��dnl�Huۍf�����U%���3zuwr?'�tT�c�ؘ��Äⷑk��<����{[8�__U�)��ӀG8�	ú�>Y�z�������Bak.sۭ�)D'��&��/z���$����jZ�%�[�� ~<D��,Ñ�K�9���^|���UڞO2&�i,u�;s|��c'��I��<-�lXJU+��}&M��b�U�D]���R[G�+��tu�ݼ1T
��^�0���-��;��U�S��SG��}S�ٟN��Q���_���;�}���b�\��vĜ~"\�i�S�EO$�{I)�/�U���>��[�Í"�� �|G�BA�XW�}H�ycۓ9�RgR~�+T�-1?�P�bcIc�`j�_�m`r�uX�0�ֆ;oC��/޵����Qgvt��AH#P���������9��kYDj�v�b��`��X93���Z�1�!Q:,�	�0�h���6٧]�W��T<
��Fp�2C<"D�F�J����E��7	�Ϳ��_eO�|���9�������["����h�]H�HJ�'Rt��@~u� d�"
��5�o����������e��I�:5M"ş$y4����(;�ݍt��w�ʊ�2{�$�X�V��mͯZ�x`�r̵���gA�4'�1�mV�I�Nw�U��5,�V������{IH�炽�Q.��<8���)S�P�t�O�������n�y51�����׊e7��{�-ޏ�����K�Yu&+�z6�^�K�Hͯ��_Q�w=�*��nf�O�>j��Z7�d����C'�%KV�\���*^��R+�̸�{�7�y�L�Ž�p*|�S�uh$�Wv���h�V�ȥ:�w�gc~���s���|m3�� �u�%{���lQΡ\<+y�TB����6���3R���7L�c�V�Zb������P��qjp�0�30
���IS�1�>�y�n���5�mjs����0(��<�Y��}��*��;c ��k���z�<j����|�K[@�g1�ō��_�3ډ�٩\�.qN��A�nbUG��AN�2��[qE��F�u�!\c���|ϛv?:�{�i��~V�(@�� �~f�	�/:P��l%�"zh>�u�ڠb����qb�(�/����}�@�Q�q�{k���7dB�:�O���k=�w��d)9��39	z}��)���\j�Դ�V�ӿ�͚ps�Цw�|v%?������(B�Q����ᕲ�E`-ٓ�`.g!�8/Ӭe��!ka愫|���Sg��uM eva��LËx�K�2E�t��k��m�����X�'׋�Zʖ��1�b�0}�/pv�A����{�K\�!҅�e���=���ا�2����)ߴ�M_f���(���4��P���9H��!��-t�c?���Α�������4r��1�N����`���P~����3�|>��+��	���c�����@̜�e�W�~gq�o �]/*y
��,�Ö�����US�;���v�q��&<�Єu��/�u:4�S��1H�ӹ5ttE�C�W>~��d7��wإo�=�)�7H�&�#�">����8?��}���x����4���}KAU0������l{� LƳͳ�y���۠�!د[J�\k��="��V�FJ�8�EcT(R�o�g�@$EV�D3�G�L������|y(�Cx%g���Ƒ5�ǭ�n״��ON��:.���l����[�;.>1\N=k}��.��a.�j� ���`�w�|z Y&'�l��ܚ>.�	;`�NQ��=v�Ě��u0h��~��*k�mW2,&�9 ��0IE�n#��+#��t���B�	[�X	1`�hv�ne�_���������y�{d�p�ѿD� =+&UIq��Ԭ�MW�:&�A���Z��u���������Z�8��`�:^廾�.����e�y8x��Ʃ��������"���/�ߞu�l8���Ӟ���ZB��#��o��/v���ʱ��)��x�4rϠ(k8v
@�0�3;o�(��ѷD������]�iۀx�6�ā$���)��8�{�]t�FW%���ʫ.��\���QRj��b��:�E�o��k�j�h�<�����D���X��W�;���@5^�����V�W���������b���]��m`���^��0��dւ3�['<�Z���|�U!kf��5��վ��Y�ѮZ�_�h�`��C ����L� �&��`��h��V�i�g�~�|��-�Y$�=�y��;T�q�Cgm��?����VwE�s�IX�?O�����buRh*"gt�˗���^x��QJ��:�L���C��dcs�r���f'X��Y�PXh��҂"#����G����<�5:�P���V�"w�hޘD�r�0t�o@�XN���l�*:]�i��f2Mv�N\�� `8�۷x�i�#3g�mdj�������ٻ�z�a�q�B�����BO⍠��8�h<c���0�_��{\��O4)yt�1��묅UMS �3]l��T/�'F�ë~e#;���a�Ӵ";�-�:b������a3?�SV�~	pe���
�_���N_fu�v��]�T����K���+T��haz�<��|jnq�B®��z_����Mؚ�E��1�
"���:�h�Z��wi|}ۊVçû�2�׺tӓy��V����p�Z�.66	`��+�i�S��C}�O�ɂ��kVM%�sȧ������;a"�����ަ�����Oq5qA�����7�8T��D"�
��(�C u9�t�7O$�1���G�!5�%A
��I�Ɏ1�p�,f`\N�>�mn�Y>$w��l��s��8LavP0�3���L�EcX�e\5�H'�ɛ�yG�\ ���۴-��x��Sr�C�;N�[�h}k=n]f-e�H(y/a���N����ޝ}�V ;�a⪼c�)	�W �b&������U��"��UK ���y���=A��aEkvYC%ZT��h,��}�R�1i��A8�;�}�ƕ�Z�W);k��]ԇ����9��$X҆n������4����7�a#�������NK��Ic�	���Y�~ܻjږұ���}���#Qtj2�G@���I6SqDc�� �^RP�nnx���(�������p���f�S5T{������2HX��r����`����t �\*�����X)DA������8Z���>%�?t"^>e��q���/ʡ��l�Q-3PY���}6Ri�%RP��Iq�L�NW����"���܎͜G��{���K�T���A\��*.���A�L�G�]�#8��q<8��ʴڂ�Կ�LCӪ��L��-&�� g� ���ib�̀��i0o5K	5�!0 Q��L&)"�蟷��b��#��4�e%)铵�i�F������s�
�f0�N�=�0�o<���!����b[���4V�������v�ʱ_a���ֲD5����N���J�mM�*;˻�g�m�F����_�2h�5~�Toa��=Ɔ#P8��y��x>~���3P�����k,LA&���~5 ��h��rJ��[�f�QyxG�v�pG�c�8�,e��ɹ�Lp.�S/h[m<�3��j�h*~��b�p�N���.�AL:��܊ބ��C�VW$��J�7�.���Z:������0�K�b��K̎x��z;
VK;2��mض�ÊSIUl��'-�_ U�	q��Mp�8Pw%s�W���ݘ��H���ט��3J/d��j$�����Ru2���D�3�y�[[�:Y-�/@g2���X���Z��f�nm����+�JJ�́�o����0]�X�����3��K����m1H!�Z���t�A"��H�N�C#�`�&�2��8����N��ƞ�-^��T����FP���O{o��"~���<2��Eԙԧ\�Hc/��0L����.�q�,d:΢B>�6�qe:�Ո�b���T��  G��$K���z�p�*F4l��=)�ڇ*-��k�� ���b�.�[k5��鋙���aY<�	C���%mD�M��]�Z!�Ӌ�5���NF�/��-��/Z�d9˺��+��ӤX!�$=*��c%�ew51e�?��4|��ȣ�]�a�K7Ѩ�IL��^�$�
*��O�:N��1�싷��f�IT�4צ�39�=�Yŵo��T89�0nG�BpH��h��zY6���^������->}�4��Aɀ�o�u���ʏK����|=��������v5с����1\�R_��1s����|aB8�gJ��*�§�V�a�å��A���yk���0���k�h#�:9�ݨ�}BO�MߞE��q�z�(@Ÿ�T�l����c���9z����ˣ���Uh*�+�&ȸh@�;�iʨ�Z�L�D6?������|��U��{��I�����{ I�C�5�	�qo���h�.�m|����D4Od$|���1���u�����#�X���=�p)�U�0�"��gԟ.�s4�u*D39S�Sg�8����j��{�)���,���@�T֬S!�IPo#�S�ǍYcį$LEpI7m_��%������Kn�c��޴o	X|��ZCp���܀<�2��`ܴ���J��}d�15)Q�>�����^�ob�\��Td��mw�D%�dH�V��3�a��>���겻���c*���!ا������EY�O����HzT�\�k�J|���F��J3��E. q�,-3���iŢ[����1��"���ª�>�Y���r�8�	�m�P�ͤ�+�+z���;[��~V�����.0�o�~����ҺO���`����ߦ�
�[50��x���Rbr�Q͝��k�v2��;r�K
$Ǌ��4l=�z�m(����3�M����r�R��z���y�p�f�Q�)h0�������&�?����V���n���d7�ي��X
�yG�!7���}���Z�w����I��^����T"��F+
��oꁡez���B�3�c�"5�������[�Ȩ�!Tz�A��R�7I����h�S�w� �
�����kĨ�G�YX6T8�$��'E�+-���vb̄�L���F������Y��Q�x�,��f��i�P��8б��_�I�f�S]��Μ����l���_�c�_�H^���DU�a,	��p;P7:��݉��7���vX>F��9{�˸���p��қc��$����tN��o�?��ICw}�'Ot�޹�5X�rd_5�u���@t�]I��5����S�|��~?��#"F�ߌ��`��l�^�T����%����-a=��j������4n�I�o��V��ވ�K��6�"/(/~�m��L�+�CJ���\]�N�a�8�{9ͭ�o\~:�����ͷnh9Qq�\�5��5e�_%�x�/����X/����J�#{r0��)c�`��qE�����.�h1ol����H��S?\>��>`jtZ��*f�	K(�e��%�ꘖ��
�Rw��4K�}�0/5��v^�I���@�����:��6j��ML���1��]�;ٲD�\�^%��L��W��S���@$��b8�'0�S��\�7���ԴlMw�U�EC������d��(����,�[r^(�/�Sۛ�ğ��p�7&��N�A���b���(��u��Z�H8�ݚ���IЖPfu���	��4!���o�/�v;z\῰�"��'t�)� S�R�	D9�Zц9q_����M��~�S��������yBS ��:ZbDoX} ����nZ���ȮA+W��Iꐾ���e���|���$�,�����曭{%��橉�T� �����) ͍$C��S�mr%�~��~\(;���S�z���M	~������%�)�V�d�#�w����y�^��d&h9�)YN�UL!4�w� 2�ם&t�Ǵǚ�50��N=eY���#�@��f�OF#�Yt��<�+�?v�uɜl/K�C���%\��(ߓ�꒿\����1ë�����ӝD4��oW�}U�%�OՄ��
3���L�`hAa�����������|�%Ϧ��;�ǲ�WQv3ڷ�2KS���#�I� �B�ћ�J|�:	_�#��\�QQ��l5ML,��'�����MܸI$_)�^B������)Ɲ�� �aO!�A]V�7���]׹d����]�n��{Y$���/g��/@ӫ(�S��b�����F��Fĵ�'�\��&Y�.3����R;@rdb���:�>j���s�u5q�}�'g&<���S�J����WRk�f�m\�
�o�
����
�A�����M�uӁ\v�	�p� [��Y�6�ŝ�n��;r���VA8S�h�zO+yx�3� �.��#l���E̾���_u):����4�-�����p`@��Po�Α�l�W�6�6?�z;]ӹ��sv;
����M�x��ÂY�(-���e�%_�K�#%؛[S��D�<�X9uBO~kkH�q,��i����mc����f���,���aTd�9^J삺U>N
'^i&� ��o���uhm��<b�l�^#���ѧ�d{ld�1_U̋p�s��y��I8�,^H��μX�ڱM7;/MF�t;�H��q���Z���Q�K�ZY�̢�&��O\�Z�N�����~/�.va���y�#e7	��i��ǅ��c-��N��..}0t93��1��<<��<���?�]w,�r��X��#m/���!�Cc&�C��x�Ҹ+�QLE��;�����p�ôc=�i�pR��/�_±�c�k­±�ެ<��8�>�����&zTȵK|D�Z��ڵ':����h@<�SX*3R�j�f1��������z�b��Yyc�x�	C��&B���jP=6�'$��Jiy�f�0(�7��6Tz0���F/`�P{��Z�&'�`Sp��4\l5��m�4E
���.ɳ�C�S�n��rنk[D�J�[�7��x�9�a���<���5-��r=ʊu��uB�HUrr��M~�GB��}��9>�4J�-�kQA ��NI#��$p�$OR�Y��d/ޚk@���d�g*{1�������ɵ�T�lnO��T���v�i}̰׾,d+�֎ �E�O�:nӦ4�6}��3D ���6c�w[t[�Ȁ�'XІ�j�;n�B0c<��9��ET��m;��E��&��a֡�wFՠ�p�%�ٝ���y@H|ۇ�+�@s#A���K�s��2:�u�te%u[�R�)w��o���{*�Vt�:�"��9�)���������� u�3�VҮ�f��kA�fx��؂�W.������5����*`Q���@)\���9w��s���z�uH���v�S�;r|��\�������c�i4�����lS��BE��>"���?lz�(��N�K�8ʶ���ڍp���UJ�T���M�Y|v�����=J�Sx]��@�:���u�n��4h_�ecC�9mp�$��
���$ΰ�ii������P��!��T�$,�qNF�q^�in<���X[z�U�_�fki��A�O��?�kiIF�fƺ��������ڠQ��>8����?v��M�E������H�A--�U1t�3�6�"���@������^�h���x8��'�L�ķX�+"�t���9�M�`�ɓh�p�8 �"���Z�ni� ��hՕm�L1E�`�� ��"$����cl���Hw�w���7��$�7�,o6��q�KV+A��F��p��W�+�r*f����T&�t��Y�%"J���-փ����h��Np�d4ya�!ɍ�p� F"�H�[4z��A�0��ߣ>���$ljY���	�����9�*X��i���>6}�.������W��0	Lʶ�׀ds����I4@da��h������ZC�8W��7tGx���_�u�+�G���6�o������.d�j�4��DgY�-ԡn!k�%�H�錌��?��$?��R�ͬ����4$�k�2�i&@_5Y
R�TɊrA.4�9VtD�����x��6w�oG(�ZPj��+x������,B�0�˼NiT�A�{(��?8˰v�)]'�Un�f�l�&��	�\��Wh�=�T�6v��èk�xq��Swg �]�	���P��Q���op�URL{��S�ه� v7
B���P��C����;U���t�x���|Kx-H����6bX�N� `_p����CB�	H�"�o�,��z�|���b|�g�@����{��iaI<�l"��{�l$ٺ%�Q=8�w�� ?\$�A�N�\!�i�I>�3��\���,�o�;y��i�_`���-��3q73R�7#�h;oM2T0�P,��"�M��L������9�uB�;��6�ՓP���騶��O�h���HlP����(>�7f#om�U���RwG�iŋ�ya:�ڂ3E�g���2C�U5O��e�S}��[�ǝ����T�ˁ�S������C>h$�'�^%_A��?�	k{�ZA��it��u���>��,�5�XOV��d�<��͖
ڡ�f�ҁ�>�����C<�ݮ]���0�24���]��%N���/ yJvQ�Hg���.]⣁-��K�f��MZ��6"�J�9�ga��3�f���2��=�M�i���fR�ݦ�N�S|eZ_�c+�h���}k?b����׶����<�o	X��~� ��������fw�� B�B岛=O�{��1�n��CL_պs���*�A�M�0��
0zk���=^,�(��xU�b����I�"�t�S3�* �A#r1j%/?j���\Pd�[�3D�\�쳿���(7\��j֯��΢X������vՂ+�`�u(,`�bK�Z���,Ufa5��'q�mеG�a[a�·��IH��e��5Db�r������T��B�[1&�*eWe癜D��t��M�T�q^ ͭI�@���dĳa�h����F���0(E^^@M:sJu� ��x���˱)��e���>��]����H^�E��s0�m|�e�X�L]m���3s3�1�E�\��y'Q!~�����V_fA�"�G�_9f�hջY]�Mt?��uꔗn�������~�<�!4�>�B]��Mc��u���Y^)��sY:u��+˗�<�����v�P=�>�}�l(dAy��pt�vbc/����y�c���A�HY�$�*z��W�l�t��,b�T������HPV�h�Km��4ĴQ���[�]�]	FI�-�M[�������E���s�q谰(Ӓ	Ō?�u�ҁYWnb��z}��o�7��1Ny�MDa
�L�� z�X�r��n�X{!�&���`�x��%d�x��0	�V�#�'�:��fd���R&�L���� �t1CM�%�Q��E
a��M�%>H`ˠ6�ۏW� 0|�M�}2�k�k
�翠Wi��0B_�����Z���a"N?,�|�R�%5t��KWc�g0v�!��d���rL#}w�\t�2�|��	f���,gg��gj���5�/W�XH�>>	�c���02�-�D^ �|������$I5v#��'�'eX �+.vee� �YqZ�b 0���������.�����Indyv�mi�&_��Ov��d!(k�u[��)��fۙʗ��cш�"��ӎ���{�W`��F��<[8�}��d� ����f����ķ\�s��y��gA����}M~x�?�S�-a�ұ�(�����.���d셐��F�NUZ6�g��w�y~��0����c�E����c�	�?g��GЩn{-�&^���{���L���*�N��?�� OD�z��mm���g�wA���Hg�( Q�CfQ%N��>I����ԤE�5p��a��6�xh���;��U`j�x�C���;�!FC\��rQ�_yA�-,�$��v�#.��?~p��ܮ����]1�1C�$~spu\�1��a|�z�\(匲����D����U,��3��T�mR��n�F.urE�"V.���cؒhtӆ�|�w%/����~W�^�r�.)��m���3^FO�\o�eщdiȥV[����L"���ъ+��glm���ꇐ��tv�'gT��4d.����J�xF�״�n�ٲ?�dE+��Y6�#k+�`�K�V0� 7Z��	���=��$��';E�%��7_ݴ���P��3-�e�!v�����*�J �*5�|�o[�����Ә�-��N!/�#����k�ᵫ'�)�Z��ܰ�J>�А��ʅi�.�;r5���N ���;�:�vE`~+g�?o�܃�Mp��A�uT(�>�?�ء��d�=��*�����/��� �#����Ѱ5��x+�P|���H�A�R�Y5�m$f,�Kx���]������&Q�i�㩠�[��� Օk ��k*����{yvH��H�lOe�?�^���@��T�]�<&X�tq	47s�3ʦ!��0�.�چ�ψ�Tx��9ML�����[R�v���J�'~.�8RcXv����c�o�S�E��م���m�ٜ^&�U�ꥒ`�@6o��Ok����c�#D�S����vOϺg�ς7EZ�t��p�:�Z��\�&�3b����z|mP=3C���
4z�eM��<�zL�����)T4*,b��!0����1�l79��wLө~gP	�Jɮ�$��bC%jeĦ(���z����.PX8������U��3��ɍ�ta0���%��Q����ĭ�3,��J�λ!i��5c�O[7k�W��;��Ȁr�C�~~�?��G�P�ȥvŒ��8%xM�F�U]T�-�H�+�������Ќ����8NC�E:su���Wm�B�
t<���~&Ѵ�����@�m��-�TG��@!~��!̬*?z uH:���fא����=��^�yS����ҷ_juAe�S�Xvy�E�e^�$̪e��/9\i�x[�t�׹�0�'�VBf^��u��-�ǒ�"��!�ߟq�<����j���V��|� VW�PaOp.�S�����uI3�%�Ia���˲�����X���OT3Z��<S&K�_!�B�g���3��$9��9^�K��>�\��Q�x����Ѕ��"��;\)zo6����*<p��<�10Bk���Y��^r�}삤`�����^�3ˋ��)S&��K~�6��~ȡQ_N�}�6F~��җĩ�Vֳ��yA�G�-�b�<����1�sO��m<��j����f��T_�ݸF4LeG����:�g��|��	0��b|2���,��������O�c��=���F(���j�W�wg���X���'�>�&2�47�n|DѬ;��#tÅ���h�@��&��
�KzY7�������^t;M|E�<`��Ԕ� ��6�a�|g5ܘW���sz�}4YyT���RŸU1'�W��6>q��l�]���h8^�ys=���9
�b&̙�����,SqhHۊJ򋴬9�./�	Q��[�wX���Q�<%���/��X������|�g&-�h<����<f��(�&G�O�p;���װ ��4b�h(��G+���D?		Un��
��\��6 MJ�3O��E�Ñ���Y�=��C*m���&U9�Y:�i*Ikp��(φ;lW)
��V��w�����K2Y����H~ە�edk�Y�:`�\��?�����_:OY8�q���z�M�́��托kM&�ŷi��D�ic�r����xϨ/;�-�%|G�S㻄�˰Ū7_)S�YV���F����J���1����v5={�9�,�FeR�!k��l�����Ȃe�ɬ�e|��4y�B^�����[��kZ�9�#��\�鏙d���i4u�v)ÿ��zt�I!a9��K�M��i�Ă)�&dDF�`�ͲBE�^&�T��O�G����q�|C���_��D�������:��/l����#��0*�蓝/N�JaJS�uү���6o�{�ͥ�p%ʶ��|�0?HAv��,pz�of�� ��f��0��%����Bˊ9,�^���$R��Ś�"�°��O��~
+�1j��Xiv��]�V���aL��LZ�9�N�2����݅��^F6;]0'�E�J��K�v�A�6I�4M�_KltB�S�3RR�^[��[έ�\����8�X�'����.�c�wJvu��Im�2�G/'��J�R8�v�Gx��A�}'�f��,F_�m�5낐$V^nnN�9�rN=���P&���R�R��48��\%�N�1"[Op�ⰼ[�*Qu�o�}'���sA�z�&�����8�~�S�=�>�k�*P���¾�����w(5������e2e(��>x�b���U'����z`�Qq&ut��?�
6�'&�0,��hc�b}�~��[�RULf��O�&8bO{y�dW�X�������#�Vl��(�+��j���f�ȗ�zJ�d��*�%�Ga0^�rZ��}L�*l��7��/�	��v�,�j�}���o(V)�,��sߵ���n�osn�ʊ���~����_Jږ���C�z�#��^֔�{v��D��2�������-	e�fjn>?�͔��5k���Kڠ�g�y����ܼ��C�u�s���8\;.I�ax8 ���d]��ǯ�.�ˏG��6y���HZH�9 2���M��5L��M4"�*==�e�C�H�J��m%kk��ξ���U��a����_-�kC��R�u��K�s�s7~����g��J�i��zP���$�.��Gԧ;��V�2.����׻�3��joi��;�ѫ�c��^?P�Ac�: �p� ��c��aM�� !�̇���Xqc��b�먆���|j�7k^o�5*��(����D��R�)CdI�6S�7kO�2y6,�+8��$�[�J�/偿`0��0�ק���������yx�Y�-��"������X6��=�Z�������V�g7a;��D-wAe�8�c��DD-�8y9?*��|�z��lD��V{c�S?����D�>��@m_H�tj��n�YP['��~"�I꩑X'�T�r^�?]r�
�����}��ܟ#.T<O�IJ8�R&T|�f,n�߉�c
�ś�SO׋�zk&��Ls!�T��gD8vG�oSbn���D��quO��L�O�V+f�]��DJ����z��e= F:�W��j��~�E; �c:r�������:�IR���جu���xE�u���ș�F\��9��].�;\��\@PI�q
����q�v�(�RH)���XΑI�\�Q!)��ծ���!�$��	�!H����y�����u��.�b1Җ����9�9�ϩ,��Ҹ�JSס���9H�=}�4���U^���W��}��[dF3M��O�V�y��K�����G~4�{�GHi�x�$��⎳vQ�H�}�L:��@s�hŕL�/��4P�>��\g�H����\�i�B��20�����=�3�{=�׀	�p:ꊭ�F�b�
:<�r�(�zI߭nfṪ�_ɉ�ƥ�!�QF��+�1����J�8��R���9��R�7$��+�7f{S�֧T�}�-6`��W���RF/ˋk�'^>���/h_񲜍�(X�b�.�3��U�� ��JiG��?�G">���SZ�G����<A��6�q,�"8�����-�p`�T�4N#=F��e�ݧҷ�1y��Q�_�:8Z�UT�NXDj�GMy��y�	3��(vː�1����/@��BL�y�!L����h�����*���{��δ�="�����/����Ze*zY���I�C��lv�^P:�&����2�L�mDnc�=ծre����%��As�������&��8h��-��D�0��S�V��O� �Zv�TDĊT���w�Q� �)�5X2�!
��l��쎬tp�~X��g���u��)hK�^q:<�b��A� �ە<��57�?d^q���E��`*k���E��R��MM!�ݑt+��W��K	�	1&r���4R��#f�����o���qX �x��"�i�n�x���*�W�.��Tt4�Iom}���B� Ѡװ�Ҽ��͚�a���� �5��j�O��O���n��6DY���XBL2vN�-�qȽRr�e��9�A�_���v�H�ᚈT�^<�@���3b��k�鞢��T�f��Iر"e�8�
�"�b�����{�}����H:��̒!2w���r�&�������[��̓��&�@V2h����A��CL�><���ۺ�5�Q�������N0�˅PU|��(�!$�g�Q�7��!�ov�т9��/�Z�.<nڙ7N�{�^��r��6@:
�0����.]M̎�:OK��P<���X{ +\�%�����|V5������pUy�!S`�ZpFǣ��\�$�bh�����D�`�$���V���;��.Ѡ�:m��N,)�gJ�;���c�R��M��Qc0�lD"#��pe5.�@�Tv����L���B���M�E�0�]�D8�rs�M&���c�s�������03շ���D������-�WuK���t�-j#�\�v�+���X3��Vm#�������x�c0Δ���ݮ��!C�t?��m�����Q��l���P>u�T���>u���j�n���6On
:<@ 4fs�}q9Ķ���A}��c�p�ۣ>ټB�!�FY��N�oXa��k[]Ch�m5���p�؟� �p'@4�����?<d�xlul�S���@M�Ϥ_�6s9����}����;/��	O2�����I7\��п鴋ZhG�cWQxD�%���p�W�7�P�p���2⣂�t07�1���J�G����p������<k[a[�o	�0!�'�"z|�xa����H�a��u9��)ߣ���7{��7_
�Z�"�O^�$��w��⹍��+�����z��p(����8f��5:��*��w��i�4O�v��X��ae�c9����RJ �j핅���K�w�o���N�N%C��2�c2쩲[��g|��z3����1}�ā����t�&J�?!i�6��?n m��x0e�6݇���<�*�t��A��|?�% �|8�{(���E`E>5'ת�q��P�d*3�W�k��KHr�U|�D �
0癹}u"��7�Q|J
#��=��9�~ ��I��}�6W�k�H��r����A�����x3��\f{��dm,�ZU�1y,F_V~�A�&�ڰ�/���g��;7��<�%S�Q!�j�;�`�zʈ;����Õ~�{��6/������[�*�<%͑b��S��ףj������F*�=��TOP��K0��?���	�xE:�x����7Z�4����������i�H���e;�Z땖;�K����\��qP��3Z�D�*��]����Sk�fG����Ie�K�痈�In�s�&��?���h��5VhX]K�=
WB�چ�g��?�<U"�V�L��6n �Їa�y� �/�sW���5y9�`��J:6'I&��l�q�ڴ�� ��, dd���3'��Nx�B��!p+�Dm�ܯ1��0�E���ϩ`�~ڼ-�kXZ�?� �	Q�^̯��� 법�ZFJ=.�<�/�&Ǎ�Zw"��9Q�tt(���t��5IK�R(S/�ge��&ڍ�Do����(��[�4��� ۸�c(��ov@0��w����t�뾦�HY����qa��}53!\W����2�n>�T���Kn�bJ�bk��X�9�77��g�̰�"�c{�h�(�2;=.�D~�-A��%Y@ZrTw)K�B����.��D$ )���޳�Ĉ�oi��0�.�Q,��x��)�e4w��/O����u۵]t7�R6��W�žj�GG`J�ט��K=CZ��H�UxF �'_�j���F�^1:��*��g���֜�%�,�����Ճ,&"�8����.Jo�`�Bt��L�RG1p2י;��Eu!e�����9���D�ī�nG��luy]Z�l�P�F��YYT���(/U˲1���TH*�P��h����v��s����]�0a�����a%���K�ׅ�ZǬ�ٔ�v���'�u�E��G���?��^qy��&�)��H���y=�%��+�YpP��NzB�BX�gL���p��;Z��Q��=br����NLʧ8���v�;��@��LFk�ЛZ3��M�bݳF�i�K�c�;J>>�(Y'�C�/�^��õ.y�mm��G�[�'T�Q9��/?�M�c��`b.�|2��M,L�h��!2��9/V&��W2ۗ�j@�KHp�4�Ϊ�� A�B1l}�a���z�5�.\)����q�|��.e�Vd3�����@�3�I�7��Ho�S��7"�GW5}��?	 ���oXU�<�՝T1Za:^��ZKc���(=�L�#��jO�)�m�ΐ� �W�nO2�6�K�ԅk}�aŜ�s�m�c�H.�R7i��6�*~���w�� ��;WK�e�^%�?Jg�ь�\��V�~q;�<�@�~o��K����0ޚ0V+	�^7@�"�����}T�����{J��
d��49 Z�5�{��Z�I���ZxlV��
��R�,(O�bo	�j��c,�)k��#���N�۫x�
�>�ܧ�7how�8Y��z/��6�1�'�Y��\a-ʯ8b�-7����6爬��ȷ�f����ttʢTV�=.�Ύ��2�* ��p2Y}���>�JA�R˃��ݣ��*��=�L�
��,HE܌Z���޳�=O�XFƂ�lP���}�}�5�e�l�F���P�9�j0�e].-�����yk�-�ͼ�v����5�|��?7T���9e��v
�|2�hg ���s��S��K˳��e�OrK�w�z'�
9��i���_K2��m��"�tkϐ#��T��~3)�N��x'�:�~(��(m�Q�6��IǗܟ�Fzۣ����Lc ���-����@&yx�RK̯�Kh{!�:�C�i���;����+�#h��²�H]�,q҃]׳������O��179�P�����R����iX${CQ�پ����@7���{�Ժf�n&l��l�N�]���Nb��?��s=1'�������̸����$')Ul�HI$*� -�K���� ����ω�I�(�f=��%�M�^e8'�h��%㩣�m>;G�l!L�r��^U���~��.l���Q:�s�LpE5��1��z]6��"���:�l(�#|�=K��rO��&���C�~�x�_$MN
��[���$��*G�gP��Z 0��]��"۟#gݿ�l��5�I��
�R��K(a���UDf�5����}}���)���gG-�lcKOji�D�f�h)���4����+;gGE~8�,���ßc}hJY~�$�Ri�B��Б�|�5��7��8��W-���#W-n��ͮ�'3�;����SF�?�}�2�pQ�x+mZ��LiRImivk�����Zu��E"��'7��|�a�_2e���4�[V�7A\)�/�Z����c`��֚r)I�v����pY�M�8|��	+�������E�2�X�B��E��j�>���=�w���>�t�̱�8�+�)UW㶆��I�G��ە����¨���3T���UHhO�i?�ڂ�	g��1w�� �w���f����H�B pٯB�v���\��}�wXa�����d�O�R?���rU+��U�wLb���E��\�M1�ʥ�
��jHF+ؼ�m�dpe�7\����vXc�Y���1����M��Y7�ٙ��w��ӛԓ�d�8�aJ�[�%LO|6[U;/�ܣ-P�в&����E��
A�=���z��;�!8ꧼbٯ	�x�i����x%�&�Vh�}R0��C���!m�U�Bav���ݍ�����O��$F�����C&5����'C?B���w��n�J��@��<�.�{�3h����L�tD�Qaa,�5v|�j|�j�����0���Ne��O��(� ����eTx$n錾��Ӳزn7D�-4�-���z�^r fW��G���a:������}mq� ��ԥ�E���O�T�^�53q
�^t�q��Q!�_���ֆ���_%�8]n9w���ٖQPn/�H*Z��'��Ů\��{������������=���P�mZߑ}��j?���[��*<����_�E�o�$�rD4R��y-�~��!T�*<���|_��	���9�:$�Ne�l�v����	�ǽ� �Uw <�@�ZX��<��
t�	���I�V蚩��ln�K\Y�E�>/c�L��a�ڱdaP����V��{�`��<�,����	�˜�M%R�"(�k~�-3��-��I.MCRޢ�0�\6*���|`bfJ��k������+�Ѓ�����-�nM��T���'�nw�jt ����A��Z*�^���HI����{�5[2��gTMYz���*���" �S��D��"��z�JB-�R]��A���7qgh���]R������C�'��,D�1��D��q.(yZe�'���R�-�����c���٭��ZCOXݖ-�4�@��Br�yc+B����6�h>;���M1^� �c�E@�2/і��pXL��!2�t�Q&��/��<^��#l"�u7�Y׼�fkA�p���N=����� K����,���1v�K��Β:�*fNJ��|���0N�^�#v�n�|�B��|�,1Zݽ��V�]���B9�o���4^B�u��+��� ���Ŧ�9��7�	�}F�t|�MLE�Ћ�������v�-U��NQ�k�J�EU�#�@T_l�{h��%�Gm����M�)j�-��M�cP�����?vϴs5�p��h-&��'�<A}��.�3�	��W�{jY)�l�L]坞}Kj��.k�MJQd�,A�am���ӛ: ��{���Z�`�0��J���8��AL��g}�z�C�0�O�n٬�e��Y�?�O��o��*9�4/o�J*殜ļ�dK|�V�;���ˏd+� ,���yw�Yo���u&/ɮ�Ye��v��� �]�O/b]p�fKSo�U��|HO"�nS0Vi��Q���)��1ȸ�I�(�Xz�n�W�vN�-�A�T�h:�g`�N݁Q�5#�{�:a,*��}T��CK/�d�<%*���Gf�ڈ��S|�*���J��p����o~8H�=z�7�r�S�b��ς]�ٕ�fP��Cfk��N+1M�^.�K�	��^1ݼ$�����ri�^�>��j��<��h^�#���QY��>8��/:1�������`,�̃���t�tz���q�qP��x�o�ڛ��ص�67�آϧȝ�������C'�<� |�Pf\��21>�.e4�|���9-�΢��D�ߟ1KK��L����@��SO�k����Bq��Ē�Ļg�G��Wn��O��S��/hOo�R&&�	UA�	�o�Os��I
H��hP���any�Yt����ϱ�W���UL�v�>δ�z�P$�n֢��qȂ�)4��S�t���o���@A�@z�K���M5_~�Q4�z�s`O[������6���U�s�bbDU��(�"�RC���ߨ+��KT3�@R�zV@0��B�UH�g��1s�K��y�V[0�v����0����Ao�_������q�LLp�p�-'�@1��#�R��(���Jk�X�o��=�[��K��÷�j��j/�6*�� �R�pح��\a�� �@�")z�c������Нv^0s馓'�aw���X.������g���i��{,W,x�����Pj�{34��`��5�����
����E�=Z����
	��Ǿ��[N�\)Vm�ǍG�0��x3W�-���UD�qѓCxFX�<N���r�N�)W9jº󡱙1�.Z�,\�3��:��~&�lZX���`��������l8Rj&H�H�1�{�f��_x���j��!(X^�?���!?�A{d�w�F�%�(��]�L�9(��F��9�W����<3իo�����x�ˑ6y�kA&��¦f\*���!�*;�ޣ/��ˠ�5	�v�Iog�\��ι5����Ү��|@^"!����i&�*Tx�~�j��'��,�O��e�[]��,W��G�P�"
?�" �f��kڄ(�K>�E��!�o5:x��:�_D��Î�w�9��kNg�sݝ5���9w�k&I���9�q���С�9f� ���D[�6YXZ���Ll,��y�/a|6^�*�3'A�P�
���Y��#@�?���!Z3����!�_����>Wlށz�!6Q���6��Ȉ��`���]�i���k?�E(E襺��X�Yݎ{O,�)Y��s*�J0뙌J��o�X�:���43(,߸*�:�J}��>����P�{C��|L��oÑӪ�I+�O�֛��U,�OE�{R��>��
��`�����w�k���$a��(���ɬ����~$�'3ś8�l��u��^ͦx���_��
B�d/t�ѧ��	W�>W�@F����u[���9C7@��̢���ˇ�ذ:s1~(a�+L��(�(��%�j ����"�>����#��iEwy5�YkO�%���w6�{Z^Ηܗ�T|/N,-[J���}��Ij�� N�f�$	�A��|�̅k"Z"/���	�2(&s����&#�)*G Ei!���L����hT�rε��n;45f�K_/��c�kþ*}�g4�[dS���-t�&�,-��C*��nh�L��A�R�<�~�4)�\�>���+&����C��#��l�xp�.p���}9�Z�z��>9ei�G"ޙ��O�	d�r�A󋒍yU��P���&,�~NbL��n��!�|���)���G�7��b�u6MJ��jQZ� KűI��n��e2ߝJ��s�G�\qs��#�4��s��+c���	�'��%��5��@M
�U��L�� �A\�o�O�It�L�^�ԧ��1��X���4w����ѭ�g:�M9�a���}���yp����6���c [�B�FX��uMP�NoD[�n9���,�{j����tvL��s�+��J|,Q"ϑ�`t�2�J~|���ފ���8Ŕ���R�<��i`��wa�쪱.����h�H���c�Fȣ�u&���[w�*�V��j"X�c�ߘ5Z������MgĖK�eʖ�m�(�Ӑ�6吀�Wt�4=C_�[�s�l
�#�>� mψ��]J�μ��IZ�ΰ	�)���"��'\�qdNL/t�	�����:�n�s������U�~傾+�2C�TCPwT}%����I⢤�/Gї��0o��y/�gf��O6 �uP�+(�s���4��q1cj9M:�*+��H�)flE�8k$bh���4��Q�O.D���p�;'5� o0�y^p�Aa�@{����B��3�:/%���V��9�p�y$����6q��=(��G�lm�Y:��ʗQb�x�3��R�'�cQ>H���ѣPnn�sp23pGO���t�#6?�F��}��Bי�A��S� ��o��y�y�ۉ�FTi��{|a��)Ƶ���*����9Xaz�@����*�Bj��A�}��ۘqHb��Z�q�'c$�����=A������[���9�.GŇ��܅�h�U�9�$2�F��k��m�چ�+���H�Ft���M��6X:�JO7�
��W.��U�ryd�|�s�{��;ff�"!)�$]��cY�������,1�S�0T�*�!��(ʬz�`��m������I4��>y9ߑ��#�����=��Z������f-�t�'ü�_ R��B:�E��6S�&�s�E���ff��oXf��&��_���#�h�6Z0b0����E;����S�0���c�`736�!ΓǙjO�I�	���gK���
F�?�,&v(6~(�~��X��(��Y�R��!b���[�8���Rq������<���EE\.bߒ�0x�����x�|�*�a�p17Hm+��$�n{`���ˈ��_C��0K���j)��@ҿ\<P��b��,��JI�$[����"�������\F�+ݢ�~?�n��X�@eV) }Izn��Iؕ*�	�^�:��[N�w�5�|�^3[&^Ԃ�,�*�iJ��]������O+�.��:�ﺋ�O�@��\�[�Wd�$�v{�^_�}���aL'������Aiu�a�c �Vة��H���w��.�����fCƇ��y����uN�����p�Ya�Vw���@ K"&��	����Q�H4G�@?��<���&緔�|Y����v.�8� ���Q̃Ŭ~��������CN���PeUU����@'���tDK}â�M/ڐ�dw)'�_�U^G� C�J،҆f"�Q�Z����!&�M,�;�i����q��#��΢���A<����Q��vqC����W)y���� �5��b5�԰�V�k�����2� �K����������ԟ�&dSFE��/l-��d�ڶ43>I�_"�\j��4y<lL��n_��Y��9C��{̌�1�������*ȯ��lA$��T�x>v�}�>�`T� y�Y�e����@ɫnD������	�G`���\PA�1�ۃRun����8���0�! ޛ�Ƕ~L����@��9�T�`�2��Q�o�<��<����'�z����Z��/�S�x���[��k��q�!t���9�yN�"�HL� E~�W�s�� �7.	��,���'�DD���8�ެ�jdC�����I�i���
�[2K����>�v�~%�T�mK?��'�@��q6��*!Z�)H��Jl��.jx�C�g~TYA�����^�L I����z#�ĭ�6��+WuS�xBt��M��3�5ӀѰ L����.��t�J��q]Ny�.
i���T��͉��`sW�P�e���"+)S�1
��h���Uk�����ۑ��ہ���g�&�%�h WjU԰�\�dGޡx�ҴCž0�w�{*Hr�ͬ7�!���鰈,���/�W�Q,#$#�-���䅼V.���c~��e$�q� ����yb*Q�� ���?��&��z��Վ_.�ﯻ�K�p��ۛS��3�`�﹑�E�įpx�G�YM��e�m�}܀Me�������ע�y���.΋56�v��	7Y��ր����^Ҿ_.�j��[HV���
����ҷ��_:���BJ>[A2;�{��o+|A��e���T�#��~(X<�N�7i�'�7b��y׵���b�"8��O��7�Yg�F$w�ėwtV�,~�	Ү��M�(g�ީ�|�d˾�m�*��;���Ty 0�\���13N�H �A���Ox����-{,��{	�=Z^!v�ߨ�f
*�%�;�F��'�N��X���I���Noژ��E�����6g����Pi�ø|�"㪚\�&�'�tŲ�5~�|[Ǟ��|Y����Ē�3�s������o���;����� rc�V��3}���J���#��qXt��_����Jej�|��bfԈ�rj��ԄE�}<o�psq��!��9p�*�"c����*��3����Κ�o�X���ʝ�E��'M-俲.x��p�8�� �}@��4����2ط�}�:%Q�� e �-����F��q�ݯ&0�Y���G���M��8�hR���-���?�7���OE���k�.^�+w?=_���5�t%�#MO&���-5�m^����_�@o�����������j7�z��eK���.33�ݬ�M�-�x4<��@�3HMc��"Tz��7#��aʾ�8���g�����<m<�M=�ϻ�Z�ߡ�	E�b��ݫ��n�-�����^�=(Xd���p��(�3{�W���B��������H�N�{�JV� ��.���*��jkb=m3����t�~�xH��[��Aky�&�L��b������	_g�ی	��m&��I{�����������)P.�̑7�ѹu�<��ރ7�ɜ�A?�/,�u�t���l�`S���oj:l����%�Y�:N�3Z
���s`Nv�0�֔��=մ�):�d�)�}>�Qe\�4�^�z`,����!!��l�����T�3"e�k�ת����B�&�����n�)6����y��_h�/�4HAZ���\]�
��NK�b��-��1��p8tb�&�#�cwTn<9� x��a�Q>��&ע�Ȉc|D�꫅:��)��c�7��(i�k1��W�ԍ����wXۻ&���(N��X�7,�~{x��}u�b�M'S� ���I��g�-P�z�_�@���[6���x���kh�{��:�Xo�Ĩ&{/FV���D�-y_,ݏ��aM3�&���ߋ�zCwļS�#��|�91ϐۢF�WG���K�V�/KL�l/�}N��!ؓ��D�X��j?J��� �L*��	%.��xP�1(�k8���6�O���\SJt���F�Z�ʖ\̐��K�I�y�_\����
�UQh����!(��afx�H��zLi�.L�04�MzI.��NS�7򠖥Z����ɥ$Ϥ6���(�0���]�O*��lf֓���h�ϱ����y,�w���ēm��Y�⸲S[̭�����/������'{��0��K�ѣ��]�GIT[�;�ض�N.p;xY�9���k���Ȟ������9o��虄w�hV��l������,��l��Z�3v.��h�����t��В XDm}^�v�%�`�ie�*Y�(����J�b�Th��� ���\u��E�'y��iu�-J�k���FZт9W��ͳ"�xo�A㫦Qb�۩�nZ{MyGe�ĥ��F��ٻ����>�A��C
F*R�{����
UL����������WB�_h�(�2���ׯ�����shmn�@"Բ�'����7>\m��ˏC>$L}��|��:��]�8��'H&�gΨ���Y��4�Gތ�J]��g����;�8ܔV֗m�|I
:W@��������k�(ROM�G�)��+�)�n7�	-�y��%�M��}?{^d�A����'`��ԏ�J͝*��s�*�#�(���e�2�������=�C�1nH��D%[Wb�`8G�nn���_�6U���T���뒍Nh�qZ��b�M�,��~?�Xs(#�)��B�Eh������V�������Ga=%rm&ۃ'���ژU^�h�E3��d�[�
!z�L�~2(k)� �D�Y����~�I�$R7q�L����A�Ʈ����B�#B���/�D����CJ�UZ�4W+�\��f�̿��WR[\��u��}ێ���H>bs��D��XmV��e�}�:� Ϝ��Z�@̼���jd�=���|B��:9���$&�Z�W:]�V������Q�	a��i��+~n�� �S�Ly��+��}���|�T�5�-�xh4�Wo�����!яV�8Nw��$��LVM�]��Ϝz��7R%$Ix��
�*� ��l��d(����d����44��V]d�7�䠶y>ᚃ�"˄�|��̍Cf�g��^��*;|�)�<�p<�⥖���f�4��{��s)�~ ���Z�;�t��m١�ep�5�n�YX���2�����/1����?�f'�5�m���+-�屌~&d�.�ʲ~�(Q2��d3f6u���T��1ۮ�-�aѽ`�W��
"	^��`�||���� .�@_P��S]����;��4Ђ_��J�82 M�)���1N��$=� {��)������&F���T�{\T$����x�Sv�4���  ������ZYSb����7�0P[�`T	9T�~6/����H7 ���m6eð�>�����6��k[&�6�"��iz1��TO�܁�� Ps�=�#N&2�U�c+0���>F��u�����[*f5'\��w��yv|b��=f�@=s��"M�z���%͊9~K��#׎�k`7����'+�i�z�
�ؙ���(�~eM1��#�k�I���[���H����,%=uҔ��v�G�,/�����N�/8�Z��l��t:1�p�����9��Z|�����!l݁�TD�o� �\�>Fq��a �7&�L�N��o�|�����X
H!yBF�n� hkk�e2����u��rN�.�Y�"yC?�EI���zw�`F�wy�����8�?�'*�ʁSS��Y¾e��tr��^�
ed!�*+�h�X�93�g��q-?��. ,TAæ�������t��I�m*����B�p
ȕ��5r��լ[=h�#�js�Z߲�8��6�|�࿣��������H�����)���iS�/฾E�L-��_��g2�U�im��An'§�#bu1�w�x����v��Z�d���:�1>pco����~�{nK�v��4{��߀�0O�%���m*���u�f��l4~�i1�k��g�|��Bunb��W��_�޻��F3��9�����Y���	þ�����:曳_�v>F��T"霧~=q���413��C=�Kr��w���N�`�2�J��Ӓ�R1)��^������Ju��AH�K��ǲ&�,���ʹ��(S�H�3R�ٚ�'T�
��Č<!��F�K�ε�XV=���u���_/������"��	������}��`}o�{������9��DGb�<Q�͐�m�^(�if�N8�sc[��u���ށ�v�IP?xTjB~hښ���!R��@$N+$���w��nՁ�!��T������b�$$�.7��?�
o-SO=ffT���p�ue�|{&�=���@�_�?P7�b�,�v��Y\T�s�QT[�>�"�/�s��xB~>����E�؄���_�h��,#J�Os��x��gw�`��*�p����B4�p����NDZ��wۈ�^�DƔ+*�lG_iS:��E%;�[~j�4�|[����o��D)����y1�:��G`���s'ۄ�ܔ����·N#KҌ��
�|��ojE�G<�A�3}`f诵&N��6's���g��n�J�̇V�ț��j�;��u˙�0�_�+Pp����~g&|3�8P��m�S���ݏW���X�7s�j�A��S[��t�R�U���`m���{��YLp�%��zR���r0�?�2oW���z-�/i��j��cJ|nt��-��-���Qj%�aN�$���1I��F+����	����\��4��FEJ��hp{���?s�V�3�3���Lp�V����zᔀ���M���'9��~�@π� v���J�:�lN���-a�Ө��%(��Σɖg��˸ui�r��YJ z��t_ZD�I%|�� �!��Tuh�-�Z�J,:[���~OiP�\�9����ǉǹǤ��P�TЫ09�i���vLڢ��*5�����{�E��QA�(�`T-����!�w9��yJ(ЫY��yᇵnG,�r[�݋�������Y��K5Do�"j5o�49��M�tqB��{>Q�kK�`"[)܈��BJm0�;7%^p��B�� ���4�=�����]|ۢ�AM��I(�
c&�p�:A�������n1'?����ں�	�Q�p�M��-y8�uR�.��
e(�����Q���&ܙ���M�z��~��f'<{.���,�ݶa�{DZ��#Ⱦ�j/��{���n4�äx,/ͼ3S�\,S�	iBɰ�Y�E��0֫z��EUv��/�V�Ś�9�hvѡ�_���
���M�U��S�4�N]WU=b���1���iʭ4P���v5���3,+ŃN��vL;���^��G��tg�6И�����HD�Ƕ�0�	w"Hf�"���b�\�#��Dm��,�jߖ��0����3�yW>��" �d�T)�43�]�_6�S� }]� ��#����^8:�[$"�c�w�{�X�V�e(W�|�O�s�9\� 
a��GfT�R�Ήʆ�/4��ʁ����"p��;��IV��؀E+l��C�Fx�d�K��Z�����q~�+�������e�zO]'���x�'����R�v�������h�Öf���ё�Bib��m�d��W뵙��cC2��#��M���ѕ������%�F��d	�Cnol",`wЌN�vRkuu�~��<9�/,����l*�'݋*��*߱EF�V���������O> G�H&ZR�U��oX*t�����\�h��i�@�
��P���e\�2(��i����U^�Z��n=9�]f����R~dʊ�Y��Φ~�W�&Ӳ���u0 h�rab���cS�E�lPK*�-#L ���Ju���]S�.����w�(=RlZ24��m�I|y@���OP�z���5ՓI��)Tה�;q!��٭��hķ�<��#S�qiČ�m�����8c����XA~A˭�F]��~�묦n�-���pH	Hw{�V��3S6+>����ngRžMNH��d�`�?��V|���7n���P�4y{��EXtM��2q?�<��b���+<�!d2��E�*`���� �����w�,!')���.��¾���k�(����5Ե�Z��'��ئ�h�2Q�'��&(G�SQ������x�U���L�d��o�X�������Ę��R���[���[�)H��ד�-�p:\q���i�Q�X�1	��j�_8�d�|���z��l�0!\lk�p�Nm{�Mm���vς�)u��u��&$aX4��Ї��	�_�	;,�b���I�C��Rf	��I���-CE}B�~8X���D�L�(�Ř��ELfjn�E��r\� 1����D������S��Y�L��'�,=)�JˤZ��S>ݍ#�͐�m���/OJd��|J�X �����D,�:�]i~���WC��=*1��Z��{���pDH�a��X�-�]�
��J�?l�Wcs���1XVٕnl� >����K�߳fӇ��{�5�UX?Jb%RbsQ�Y�8b��,����r@!;=�].x#�r4����r[�8~ @��ԗ烯_�|(�w����~ �o�4�+nuk9��@����U3]�	n0�F�!��8(:���^�\�6�s��^f�|�my���K��B��� N��ٞ���#]SD�{*��rC��1�r,�� ע�x�S��qz��-�����z�^�i���0�{N�o&M���#6xiͩ�Z�R��sWH�̢�y�(��>���*4A0rd��\�(#*B��K���2G�1������ؑv�	��xXE({ҧ�M��Zُ0�`��ι���S�<K>v����V�?:�8D! ���:�E�U��w��wƀ��k�T&�kuM]��y=i�ѢZi}�=�6g�0���$-
�M����Y>b��/tl���ӄ�]���
��b�a�
HB�>n�yơ�M܂��L�RX���2Z'��C��Q؎8�2i�-��w���J�j�μ��=E7ld>Ml%Od��tl��(8���LVC�#���3wZML�Bw��c�B܌�n�3.EVa��M��9��8��_���n��jzɕ=����(ʶ�b��	��}2t`�h����0g֑���)ܫ6�ݔZ/��9TY@e��+kZ�t�*B�V��zREYFO2��5H��b�<L�'� �r��k�T�b�GI���g��[���zG�Ep`�O$r�v�+j�~��1��y�\QL��/��_�G}ц�*�T�����N#�����U��J^���'m�J�Q����
�&6Hx��(�;fWE6��A�\�|/����䧓ۭN� 3��dw���;�S����V�+��˼O �e��s[�N����8n&��8Hͻ���@h̔��,)T
�T�7r����V\���4z/v��>��?_W�y���E�tx;A�a��7�N�Und��uf��ho��Y�LQ@��&���!��Ɩ�'!�>���u�����ę�)�����j�/G�1:���I**���"FN�9��tU�T)8� 5�mNb��QR�Ӽ�fF���_��O���@kR�j$�)���Ή�8���}�~�C5�����F<G���oN�Y8���o�M7BH�p�ۤ�Wv�{iܔ����1������T$t�<.�aú^7��ȕP~���:�ʫ�^6a���ͼT�Ε�fE��eʵE'E�%�,ZN�@N�-���μ���@\T$̖g���ތ�CTz�B�zA��w�n�0��ah�iw�V|M� _��︊�����:������j��l��|i0w]Z!$h
����\��4��,�l���נ��/]H��M��U  �Nq 0���9��{�b�<�l\d����၏�U Xs�`B�M�U�� �7(n����� 1�j�N�b��% � �����:dg��_�n��P���F���q�݇�8��;ʪV�|F���Y�++�+:���X��^�*=�ȔP~n�i�}G�l�(��tF1oԯ�Pp"���������HJ�E�`5y{�ڗ^�%܇ԝz�Df�C4$������c?�@�3�d��O'��X6z����Z���K�~rŽ��L�pWʤ]��N�(mQ���s|���	�ڔ��/	f����@Fi\r�-���ƈ:�Ybi֪�1v7�'%:8�9��T)��D���]β�!�+tK:С�Nh�8H����p�X��E_R="y+�.�ͼ���|G�ݗ<{�uS�xjI(G{XT�n;:��W��B���@�$�?�L�g�!����)�{P��M�?��c�3��k��Iy�!�_C�6~8�la�Q�##Ń���wv|dU�)��X��_QU�F��{�Va/�ivǾЅ�&e��Q�r`�8N�50�ߓ�?��g"�?�~o�%Mkd]E���-��9/�q��/��������\r�y��w�g���ޤ%�"�Hz���|�o����� ��v�̿��,ָ;�(�mW"�屮�*%g��ŀ鄈����*KR���,�y+�w
��lV�*>���i��9��+0�6������m��M�sN2���{34�׍u�������u��#�tP�aqђ��p�vލ��ِ>��3mh��/�Е�\Ju^�C�`	����I臙k�����&	��9����㲨C#r#�gP4N
h�o�n��p����~���bg-�F�ƫ��K��L�^�<��Uʫ��o�Z8("X'���Ul�[&W'���P������voH�q�e���71Wuݾ��LH;�-����w�}����W���8��!f�ܘ����m�A럃r�>��ԝ܈�;���znC	����w��1��͙�vġlQ	����@�e�=R?��ڒ�>)���j�6q�Q�;�q�K� �J���ߴ|�l�RT�ŁQ�H\l�.&�\�8@���>vX��25C�Ӭu<m���]ƍ�xŗ!��l]��\oI�&�Q�e��£�z��<��_F���/d=C��c*������:Ũ�f���Ȇ䍑�/*0��=r�}CU�
��i"�P}��9߯�i� hG�4�*P��rsֻT�i� �nLR�8\���IQT��uZ4 �u�)���0X���BJ��	�|�̢�՗q�����w
���W#nOT#��W��UZ�ذ�X�]fܗ����t�@_׳G"���8A�I"�^M:��d(��:M�-�Y����-���
so�{���=�@�
J蒤RzL���	�(:���q�Ų�����U#�z�� �H�����o���٭����� �>��uO����ߊ�y<w^�6�����P\��R'�D*A�S�7��������;�<�wuA�ҍ��	��|9-{�7츓�(<Aw�X}��M�����?O���q�%�72L:�V��(/�i�h*��Ք�CY>zu���V��{���"��'_(r>:
�׌�3bt�S1C�<�yEy�7�M.DUu���=�ڀI�t^� � �e;Aϓ %i�����~L2/�4�-��h��zt}x��	2ST�+]��>h��� ɥ�S���J�/�Ʃ����+��.{h �h��h�' ��{Owq�V��o�5 N~{�XDTH������!-]hFg+q�5��<窵�AY�h_%�=VB�#e1��4\R�w��p� ����i�%�(�~��1�Ӳ����`�9�&��
.w�HY��I���؟K���t�f���ccsҲ������V��OMhPQ�K쾢���>ox��;?C5-E뇿P�E%"���j�]E>{��`�wm�7�Ȝ��5
Ah��{��z/� E��	"�4	�6��J���2�v��o��Np�칰�����Z�A�;���b�t�v"�Wa ϜynݳIB�T��7��Q������ӀF��m���V�`���^��[A�U&jSB�+�	P��Ǝ!Y'uZ ��-^U�>�3���a3oD �=�o�^t��͌>�n��vU�
���QH2�a,���ǆP=�d/�D�eCA��n^��_b�s�`��-���q�FE��I0��{�;/�x�&����(�Y����i+©�L**")+:P�V�����a�-ل������Cr�#��+��-"���r�B$�>���E���pי(�2D�C�r�p�����+O}M�:jp�:��6�v�bD@opYyN��9�Z���R�Y� ���j��I&)�T�4	}9YC����M�G�ް�BbM���� b�".��
�vt�Q���C5 �L�]�U�]�&�&�ʺl�{7��5���&V���fH�mw�)��D��j�\�V�,���e3�
d���/���	���L zX��#q�Xm|r�P�K�M<�B	t��{�\I�a=���}�����#�@L �*2)vJz�7�/&��s��y�̹�!!3�}B�I�.S!�Y��r1�Fq%�4`�����{!}��'�.-�l��_�������1���|��z���Q�W
�h���X;&�#�~���ה��?ݓ3�.[!�!�ŀ�����p@� ��}��%�,*�e�̏���><�)h޲-Ϛ�b�������2nm��4��S���b��b0��2��a�C�Z���f	 �~�2��d&�%9��*;�cy`��N룠bʜ�Б<�Z������\����������JC�G��R`Wq"��h �/"a�J�5�
v�!��^��l�bE��p����˪\����EY��V~��o�/��0��b�rW�� _d8����p�H#��*1C���܂
����,d��>�ѷ0�����Ρ�S_E��"��NY��[�d��}O����B!��>���!b^�w	ܦ�w
È��$83F����O"�8���#�A��d���HkE��N�����f�I��;c�y��&nIT$��,����ҸP�nz���+��TU���Pk	���~*�;졗�.OڧV�N������.I磰aSd��f�	+9l��τ`K/V?��,��	=n�Ik�{�\��7n�A��b����~p�T����!��Z]��D@y�b)*LF���Ֆ����r�A��1�]�*�8��;�{i��>m�ǌ6t�ǎ�v(JE��}�������M�d��k[ �u� �O��w����g=��I"Y�.~9��,S�e^׽�N�m�1D�P��y�{Ӵ����s�R+(�g��D�, g��ь�?Y4��m�ܥS�B���9=\YG�(G��V�4vr���I�Z�ډ�z&�YJ�[��5RT=-�l����H��G���_�@�ٛj]�1*^��%-g��\��_�R<�i��7i�0�����˱Ëf%݂POp��S�j�d�H�P0镬��V��wH�/�>�y\�'u�}S����>e�5K������2q�F7�m��[g�M}^_�׬���2��toFkOZ���sܢ�:��|�C�����t%�׉�'�!�'��W3����ƞy�eb��%�!2�P�.�4�i�o�㰤M,��A��Ҥ�0����m�Ռ���8�b5�k8��I{�U�h���=of��ej?6����<��
�M��S���+E:`~�e/�f=j�Y{��8U�'����x��� �T)^Q�M�3Cmhx���
ؖq��S\ �����73�	������M�_����P���tAr��Z��+�cs�i_�7��?�ܫ�䝏F,�����.[��TB��c��d��ʭu�Ҹ0գ"�|)PM�c���!Y6���}�1�r0������%YZ�"�"���	g�K�}+��>8�>У
���߅����y���'�Pѿ�	Ds������&��-��������na�/��?./�����<��lW9����	'Č��qμt%�.n�s0�R��A��/Gz�����*���Սg��D1e�$c�F#������}&Yu@���� 0���v/̆o���`�g��Mt���p�N}���[Yl�j:�`ɞTwk�P�H[0��h�ĤȊF�X'��A�2w�ި!ұ��߃zI�5ᢥht�2��o�s��f���C�<�y�m����H�z�w���s����'P�7���7��",*���E��`��@1؃����2NJ�*'�,z"2�	���(��h�4d=(�]�38�._��d5`q��)G5ɩ ���e�IA�б,�c�Pm*�(�.��3���L���0��d�?�r��9�����o�a�!l��T�K'�<� =�>µ������>��!Nl�n������q���7ir�0���9U��ś�s)�E�q��n�_pd$����'Vk&a
�?��kFj���j��T�'�e�-����-߯��X��Ͻ��첳����$B�J< �ϻG�-'��uo e�_�+`����_�� �8 ���2�Ea�A�s�Dw��u�)`� =�bD��.��ώ�=��T��S�С��(bm8��T�WNVc#��EyVVq4�V�踹lO��J?]R�?ߠ��_wY�)Օ�T��9��{7@�|{Q*��qj.06hc��O��&�����pzO���z�򨩵R��62%�������a{l�|�B�fT�9E_Y��d��^-R���n�c����E��C5Eށ���eb�h>m�3�W���觇��\uk��%�.�	<&�����R��N�p�L�T6䧇���5�p~g=?���<��N����_y�b�_?8ݪ�:z�~u����^�Ӫ��.��%�>�Y��U�]��HUʖ�T��k���;P���9~g!"��e�*�UR�:�FV���p7���:ts:q!2"@;k&ܼ�����n��n:��ȿC�+LB�.& <�X/��ݎ������r#�`-֜���l���z�d��v��N&��]����RK��h�A����O�7��Kh����������Є���Ņ.<ɛ����Bt�jL�&Y�u�`�E��:!�0��㟔h �=*��ݔ��%Q,��\|��s�/�:���8U��X��hah&��u�)����"��V<���l+ښ��7d�)��KUp�� d�
�q��D�_S������N������h0�t�k�z��+BѬ����0>٧��e�A|z�ڇ%-�r�@��ƒꡧ��7e�X�\A�=D�:��MW�{��{��1l]�:qL���dH��B�����!���@��̡N_nf0�pT��@0Π
��M�վ�	3�XoھF���x�;P;�V���.ߨy�7_ىr ?|Z�'2��h跁c�K�i�Qٌ���c(	��`�Z���_�B~oH�M��wN�T��T��O�#;�S��Y��z�ߋw�A�3r��jo"���������ͱk��9�����w5B\����iG���1V����?=��HAѳz�$�!�C#闊�������i�Y����ʛ�Y`8�����͈`<��i4���;�G�7Y����`��!�De�RȞ%����[OE��O�������!�Ie�s�k��� ҄���$	D��1ϟ$;�T��LF[:T�����!}3� ��es�F�0�T$��������1��E����F�K��}N5q6)������F,��1���}9����ɰ';��w�f���]	8P0���!2�a���0&����
9�L`�H�쬗�	����眅��wmG;Љ��Q_"���g&_>�W�O���q��:�Eb��ŉ�����lU�CU���n���l_4רE���w�����Sz�j�0�ޤ�{��;H�5a�E�2����q#Ĩ��*
$�-Ȳ���:B�>�����ҏ��*�×~���qV:�S�^勭����i3ot&0q����Uɷ>�F��C��&;�s�D�-�q���9�=P��G�E�tp��ث�.�P�����@�Ϥ<���7��p�Z���h�?ݗĄX��d�1m�Z�ʶ$�Su��s����-E�վ�i��G �5z\�eM-,~
x	ӄ�m	kI�]%�l�ȍ�=v���{�ݢPFn�NQNv���xH�%S���>$��(,]�&/قD
���p�t`���F)ߪ��`�G�NB�r�w�}�78���y��w���CoP(Q�%�<�C�4_�_m�v@�� �#*]C������u�sDݚ�o~��_/$�����0I��[�������N0,��'������J�ݰJ�r�~65!�
В�a]��U��#_���Up�~j	��HW<��:�}ޕ}]5�=ԵO�
o��.O�XIK;�?BV�����ЋT��G�.�~�k���v���|R�&��W�SB�j"-�Y�.6�)�և�4=g���fC�Zwo*� 3喸.����6�@�p���0���1����=���%�ؔГ�9IN�XF{ r�a��h�T��+v	o����Y{T,��$�%a+;"�h�w����x��ãv�m�ŒH3g��'����Iq@��%Er�ǝ']5$B�W����%:~�K�H*�%�`.!�?c�,��_��o��B#���Ǳ5s���щ�'�LqޣW��"�f�{��n2��=P������q�Ԧ�b������UO��R.ӗ���S�P���$$.�e���1S�4T�T\�$��ĒP<�+[4r�8<��5p�NEz"�����3颢����@�:������ώ"G����u���#�E�~��L[�"G������in!\�-���2��*g�951�r�i�
yA���<h�A��/mF3f�hh	q��@jR\˙�g��9����F��1���3�y��?cr�u~>�".x�E���#�9d��Ӧ*i>ܶ���0�@�2�$�t-���]?vL!Ǖ�Ð�S&��#���,]l�Mґ����Ly�pg�a;L��%G��w^뢩x���o���W���xԎ*�nA�A�^{�����Vj�lg��K<�a��O	��_���tNݜtE�a�Š�&���;RuC�8,���{#�ۨl���Н�Ne;�G�n\��s��Z�R5[�
# ����4�	�`x,����*�@�<�����1;�1��94�x��{�Ɉ���р!�0��7����h���/�>���Ex�-�����z�?e�]�	�@���2�S��%�4�<������?æ�ޅ��ħ�ff/�2�]�W���س�����5r{�C���In�TsH�_�iAk�����dp�� Bϵ�v�k�C�4��z�h�kWP����e��e~�.e,�L%����'��޺�w���9&��p0��b�y�_�$q�_+�m�6t�v�N��P�� ��� ���<�ܫ=��I�;*#����������y�H��R����"\�y�w;���d���0����.X����n�����=�x����f�fC� 4B-�ӀWh�ʶ)�*�p�lML`�orse���X܃�vkS�%�82�g���qѩ�o=m��ם����:��`f<������ט�wg��G�:����c����Ii�DA��q��:�b<'��7O�f�mA�ֽ���x[$JYkf�g����I����\�h/��Q&
'�ᝪ��r�埨�� '�v��M{>���-�1g�ɠȭN�l7e�C)��Σ��7�(ڔ��G����o�Z2ޠ^-1���RC��:Ba!��Imڴ��-4�Y�	]�\��:c�4���e1)Z��Z%�B+�����^��=EpH[QLV���r��K�:��8�&F����}rd:���M�v�J���<ՋX9��s��ۺh�F7~�\P�?y���)�}�L��0���W��6ç'��,���A�߅t�k �G�0�tA�8���9V o�N�g������C�1��J*����W�K��e]���6}L�I�G�ɏT;cZr�NT���-T]�O*Qf���6T��M/�y�pOU�fO,�rM{�ӕ��wt�)�A���i���~�7��OM�F���_���*�l��K r�oheb
6W�H#�5��i� �5V�A��.njіdWmJUy��B�..6�����7��ӿ�]�����9m}�)u�m��<ό��q�W�X
���N�$�?�����z'��a��
(t���ل@tqS[_[d��$�^1Q�2�#���3��cJZ%�^=]X����WR.��L���YQ�Ng�bw��mm�`WV,/���~�%䢓6J�����Z�
�D���}�@���9��Al�O�2A�\����xk���L�6P �_h�x���	�rM����-�R�:��?���Жϓ�UR%��*�i�.e�uI˖���DM��T�O��Щk������v6�D�=ó7h,�t�1Ѡ�\��KC����鋫)��:��a�����oQէ��6��:!Ƣ d��}x�xҧ�ŵ\�CNљW�2�_��;���J�ҹ{�����x[�e��I�P&��Z� �}:�Y)4�xT�A�\(N�Q��㾔�{�g��q�ާ���%s��].HL��3��P�����	�r-��e�Pw{��^րZ�u�z*[���u<�Qo]v�%�c���f@��O	��!��$�^$��$ũ٫�|z�[	��%������⡙�Z�-�번Kkݕ��vV�6���TZ�pWB=	1����&���C�d�����{���� �5kP���!���96tV���p��	�L�oxn�[�ǝ3��� ;�����١L��z�g�+oD����2D��#�����mgV'\֮t4�����e�Qs����ؼ�8!�Q�8���+ը-��+T�ʾ-�@Nϸ[�.�սl����o�|-c�\"�a+*$�+>~�$CL�_c�X�����k"�O���cB�[:A�I:�N�.����2l�w��s����&N
p薍���T:�o��k�D��̤�X������N�W�G�p�bq�z���e�)���<��~�YrE���p��ց���Z�`
]#� ro��_�5�Cߩ7q�G�2��7B�� c~�0w�����Ǎv0R/P�����lu��`���_��1b�Q=ͺN�\�{��2c��V�ˮF�Woؐ�o�P�������uݑqn]=��� ۤ�V���`�1�e�|OD5��|����n}$h��� ��h�eb������"s&V0�$�%�R�Ė�3�ǢNk�`Y���y�oYf��U���6����5�΂�L���Q��3d����_t���Z�[G�`�:�K(���(�@���N�m^�.�!sO�/o�)�To�$��������I��w�3�m�r-c8���C�b���P��g�I�뎽�q<}��j�ˈ)�P�E������X���� k��u�$�VS�Di�S� �V�W�+�6�i��B�(x�ٛ��Nς��U���0�C�0�i+����<���x�+�$�)_���/
		x�P�F$[���<j5�}s.�6َ8B��0LY,�?�j��Y��?m�:|�mۋL&}�%ڂ��V�\�D�e�{VJ�O�C�nNLh��,O�",�K�Yz1v��Ku3�4 ��3kJ�r���H ���ZU�+���90�����L���Bm7�c�d �U5�ڗ�H��H6��@���3��I%�3�Um���\�˝�A��3����r�3B�5a�4I𼓎]B$hw��b6)~�D��/��^�<k�=Ҕ*dir�j��y��<3U�R���㾸�Q�f,����ٍ(�>7�� <ږZځ�>Ґ�6�A���u�n╇��Ӗmꁝv �H�$��X����eM#���̟`�S��鸳�˟��c�M��x��o�h쓬U&��I-=�ɜ�>�,e�r~*�~�$��������3U���T$��rJ��$k������!�t�c�I�LCi�L�EO�)�$����?{� ̾�PI��c@ƫ����$Iפ~����Qy,�P��뗤3��m{o�"6�����Y5//�k[�~�h7)�i���?[��,�O��	U>搿>UI�{NG��>=�ݒ,	�Xe�C�zY�s����{�Gh�)��.ej�}�.P`�4�P�y: V�3��H�$�-dv6��+�2�/I�T3:hܕD���}���5�hS璏��x�{L�L�p�.k+y�D[a�y;��2\C�����K[��$&sy���%����������Ow��lv+q�WM�T܌�X�7���v�qt]�Վ`����_��$ᆮ=�*�AV�3�_��>~�j1�@��dt6e-�6��2`Ov~����o�y[�li�\]�'�
V���c�N[�ȒCl�;$��s�HF;n��@I��Xsz�������ۓ���̈^�]�w�ӃI�P��z��]�0��@��
v��_��KuJ)3-��c@��\�ȏK�n�$G����m
4��/���Qc4(�>�������ʀD{��S8��iKz�pd_�vo�Gb��s�(o9��bsm%ǳY8aR ��Rn��E�GT����!��k��!*��
[Ii<;峲�2�Oi=L��:4��EQ�q��'�Ac���[*�>+
@�ʽ�B|�X�Z<�����`���.K�fxj��P,XŁ2S�Ô�)��/q��1�KH̺�ˎ�)�Q�^Vn��ł��d��\��,�3��Za��P�oſ=셓?^#�A�֏td����Z�1���B��4��$Xv�cvәd<W�$H�T�ԥ���kpPF�Q��!�;U���܎���l̇�p�]�O����������oF�!78Q,��G�k]@A0{e�! ��oNe��(���X����a�t=��w��S.F�)����3�%��F��y|L��<�b(����T�����M�پ2�{�L�r[n(���|�C�!D�%:YO�<�./�x�dq�#�G1�*~�:���u�h},��E���t�T}�|�q��
u�Cc��G�qG�^;nӬ���aX�EV���1�~��_\��:&��[��-R�ζX]��cY��Ƌ���`�o�@��D��i-7�8oz��Sv8����1`�]>����qr�R�M��%���8�t��3|cM�Äq�¿9��(�b-?�Y�p��5�!�-�v�������?yT��4�D�b1ӫ�1$�¿2!�M����X-d���iv��M�b�-��C�K�[l$aie1��7����6w��&���Y)-��������B�RG`7����#ў�ޕL������Io"��5�*h3W��\U�ʟ�9�Y�Ũ�|�p!&j���������S���K�H>�<^v��Uq��@��h��BA���}]��-T8�Bx\ч��S�R`��}�u�b���F,h�D� I�����E��xVe����M�'t{��=�0l(J�E�"1_�)��}*ߠ.!��w�rkP~tU�3^"^�j[.v��FI$���Eѿ�b�\�S:E��NRVj̇�i��4�P*|������|�NR�wZ�^��~T�2wx�+m�����bŜ�=R݉Q�7DH�4�\��]�������J��Z�w4����V��{����nO����˪���"�docX�Z%�l�@cJD��-D$	���m�1�՚�w%�e��1WUS�l?��"e�X�؛I\����ށi��������9��o� �6�@32=��m&�5Ԫ��b��ɠIs~d�a��zY+Iygl� ���:��������d}���WL7o2��U�{��zq��c>�>t�s�r�=��rÐ4UV�Ц"ɗ!6
\��|(t`'ۚ�����g�	��<�\��U]���Q�!�47����j�#��z�hZ�s{s���X���%9�'ð�wG�I���BK|<�8�U� ��-+��ƣա�T<<u�gԂ���3J��
2˂��fp�'U�|�'�O�3��87Ǒ�/ݾ#�K�;��v&c�q |�����@������n��ԕ�E��@��!(�i#@`B?[iF1�d���(�n��L�(h�ܴ���XR^5�ݸ_Ƕc���%�X"���4ML��P���6�"A&�d�l��oQ����q��L��^s��1���	�֭���Rm�Oނ�)��ǥ��o�֋���^���4#Yit+ -V��r4�HD��(wQ��z3#��r�km!}9iW3K�/�#�[�J�Ҵ�eve������<¨$��q�56d5FG"9�5\YJ%�S���hr��w���q�k��z�d��U{�\bž��2~��ٓQ�r��6�x~��al��������C-�N�Ι�v)=��>vB�)�Q-f��q�iQ_�βK��y���	�K!� sW,�13������
��c���*QM���Mǒ�Rl��l�n��@��qV7�������@wf!ڋ�2��6���#��
�w���]S���+�of�
f���@���m5�����fx~��3qO��!�=��B��
,���zp��:{���,��!
k������5���N��J�\	6̏�#��6E�thE'�לzp�aG�D 5�^N�8�!A��Z�l�&V@��
D)y�!�T�	���*�7$�K�匋t����=o��+�^�zr��b�j�,GZ�P&>�����=v)V�'�]�@��>���~�-����ՉrxPL[G�@���J�����R�溲L1�?�Q��f6�f2���	���������8�q�d�ȹ�M51 t~jX����r߆�x�E=x�+�y��ݓ��o��W�f	
�NںG�L�ݝ�������|��g��w��qj��l������{�4<�v=���x�J��:,����|�O���ަ��vM�H�,8X��&#9a�ʩI`7J35�#2@&�`��c��ܤK����Q��0�{K �7
��((
c7���g�-���@O���r�����)td�]�a���_�xFH4Pp�D�9�qo�J�0����W�R5ȸo����&�<54e����p�4M<������"G|@r�"���a�kr��-���tg2���?�<1�#�����D��*����,��0尥�3;��Tz��ո���V�{u*Bgu�ZA%�@�v����c
��6�.��/���m7��LD�%��h\��j����0=|o��٣G����*����"�F��e�p��r�5�%�C	�5t0�>�{J����^����������o�h�6�˓���8"��ui��5��b�RXw�eK����]��i��S?w��I��{tX�h}-OqPɗ.9��{�s2��w�	w0��<���%�~vXR���4��R�"�ܙW��[z���U~?��w�K0*��1j��VY�ZpIkV�eם}{B�^�{ �k��r}�R���8�R��V�i7����v�:�:)��������x�G����in&��eA�K6ѝd��t��63
d��Hi��CS��wuu<�-��C4��@�a�/�B��6Z�bRJ��s���b7��b��RD�!��%��x�B�&�.��a��$�i��9������?�~�����jBԺ���Ku�;8��`T�t��o�%:���r�|E���ڎ&3B�t�Q|�$u��E�F����,/!�W���j�����E=�Ә	;
���(l��%�" :��8��L#֙��+s5;�ç%�����b��-s.d�W3���]�ӿt/��d�-��]f�)����H��͡媛��� )�T j���ݯ�,��-����t0}�ީ+�_��]���)Սt��Rp�F�k����q��RW�"����{��y蝲���v�r�#G��ڟu#�JC�?�ג��Aޭ��Uy�2=O#s��G�Y)8�:���u��m���ݎ����#׈Z�3���G�(�X�E�
�	U"}�)5�]�B��%i	ՙ?�n ����h(��9f|q:�D�P���a�"�;Y�:>�Epk�ǃ�)R0|���L��^�$�(HB U�{-�SD��sƨi3/:�Oh�ϜX7&jY�bVܑ!l8Oj#D[�������o7��2��[	aCQ�->��Y��B�ufA[�^�q������%�VÏ�6��pՌ�p��3�����|XR��T�E�P�y����"
���v]cfi�;?��>H�M:U3��􀕀�NE�+M4�����œ��7.$�ȕvX�26���d{Ͼ�������_�"[�sq�(ò�jy�&. 벶-��8�qׁ;���%Ub�4������ �0��_���9�ɸ�	>�T
mߊ]��'O�GA����A�S{��-l���$��4/��_��Pjt���R[E��ܓ&fN�Tz��$�vtԝ� k�Z�)Z���F�X��uϩ`���|�Kz����Eu}&Bj���3;�Ԧ����D1��{wt�l���̨.�y�y���5<�0F&>i������P�N��.MlFWM���^e��oi��p�Ejza����ұ\ǐh~
ߕ1�gꡧe����+�c��@�!�(��8>��7,��fɣ�sЫy�A^�2~HG�%��A�\E��b�51�ֽQ�5�z���/nߵ�<!i7<��r7Nh�yk��&��{T}m�g��Z���y��j��\ʃVM��/��z*^��_q�$�A�ԟb���Ey��P�|��!R\�hr�W������vN!��T�Q�'A�%,h�$�[���@��;�b����|�nIo�U���YO�.a<7M�橝1J�����7��4��,Б�l�{#Fv/<��K6���rd����;�C�R�%�J�)�_o#,{���%����C���˜ x�DC����[T@Qۧ:�Ƌʦ�z�����%���\�[����[ݱ�l��;��
�;~�ϻ[̯#P�I�#b�$w�����va�����6���쭈a��J�J�`�2�U�|�G��:ھt�	Ǉ�L�đ�"��r-�|!���(f3hL)�����7��v׶-��<��t�gJ�I?��ه���Ӧ��}	��w�$Z�w՛�1���*\2n�ޣ�,j������oY`��7?�g'���i����]~Z�j�BC��Y�%A���S��*ky���w\�M�9S���W�1������/��P��"z�^~(�7~��Q)q�����[�T�;����9�e��]eWv��|��� �T����M�b\Bۧ��ia��L
�o�f$득��ˡH�6FIH;��k�iRCH��]�w� �lQ��=�VqU������M��g09��fDtТ�F�wWF�uڥ�\��5,,P�Iq��ذ�Ͷ�a��3�j5�MƂ����U2XQ�4�ǝ�����c��kٿ����6������h���S�1��	��ɰ���b6i<B8>�@?r�)��	o�p`m0&�L�cV�u�I}��S���pߗ�`�ro�x����f��d����I=~�t���&\���n�ɽ�xE�*�	@�oG���.5���J����C�h?���<׀����y�fg.���;�Mх`Cv���\��tP0dg|��6�"5f׼��!�����g��B��%p9�I����j�
���X �p�kIT���Nϸ�+l��N _�Dr��3E��'� �@�n�&i{*Z��å��c�k���J6��y�|r
���¶�$�t���"�d��S�5x`�j�G>�gs���؞�M��y�t�kC�I���j�Β��\l~z��Jt�j=�a�
��}1�%����m��	zlZ�P��P3�v[�b�bq?�'�"̄hWm���D4�]����.}}9y|tS���
��-H��0�n=����Y6����TM�x��
i�"e�'�*u
���U�~ 9�D��W�_�b���V�ӗ���-�b�kp��D&vA���-�d�U�\+sk��K��	�����].�i��>9�d�1
��n�JW��wZ/���k:�	���٢r�	��=?;���)�M��O����/�i�~e�NS�a*���s(JSr���x���cby��Sڨ���^K�Mq?�g�	�!���d��R���k����x9� ��*jU���L���^�]��Pb)����?`�W^�0Ϫ}���z�wu)\^���]���v>j�o�s����yj�%�!ț2�]��ő�M�c��{�똼E3{j�A���3Ɂ�d�b��c�$�Q99�:�w�c��<����H��x�˵����-q��?���4 #����G4��0��f�O��ˏ�D���@�ME�F�$����au�aA�?<�
�]}��������p��_;2%�ō�Iy��*� O􏺬i�� G�0�����+~$}���:�.�V�/����k8q�p�-��X�6���¤�wD?��\���_"W�es m]��$�:�)tW��!ϙ���N-0���Qb�_�YY�/|���Մ���OwV�x���b��a�s�J��8KW��,�LN����to��`Hү,L>����6A3��k�$��l�F໡V��U���F�3�V�W�yO5�� 洀o�� �Lh�C|To�u
'Q�تU}<8����?qi#rs>�w���?��P���uީL�f_O����X?���H�#)凅���;��aR�y�+f��^%��r�z^((~��V��~�6��ڦR��R�@��S)��F�i@\�=`(o<I�
��w���x����ot��N�.2,�l��U�6����zC k@��c�"϶[�Z,Bh*���q��T �N��Z�OD��vɒ��{��"����=(P�K��Gh�l��\'`j�H ;�4�2�%�JwSMg��p�wv6k���!h?ޛ[6�;aAw��X,���(�j����)-���	p0.�n���q�.�2̆�"��F�҃���n@r���w=c�`�n^�'��fo�A�g�ZbR/�og8~�uj�������aV�)�mS�r��<u� �hi���_�H�U�1n�n\�[�{��EqVy��FNR��>��:�p�Y�^��n�~ڠ����_�� �$�(�lڦ�#��ｮ���#���{��֤�LӇ��(r�jf�K���^\�z��ڣ�0oBhz �!�ɘ�3��-aGP��qǼbaT�\��1�!�V#;�xˀ��k�G�+jF����Q�ɾ��M6�_�^iQ#��5^2�w�$a�#�r��E���y��9���Z����\ż14������׌���5h�I�fX�1q��?�N)
]�攴������TC�Y�ieBU�C�5ϥ�D{��> KO$vI5�!YT�5E}�C���wtc�����^��ó��HT#�\i�L�3Rt�� }���S�����qԁ0�1�`�Ջ�XL#�c>�\3�0K�_[�7ˁ�����"I'��*.�B�ޢO�6ȯLN��-��]��-�=~���?��r�M�z$�.�tZ�.��g5Ԁ�Y`�����x�ňJ���y������C`�v����l
�l�	;�)u	�[>:@�L
5U��&#��
_	僎�lm#A�v{4*�?-]1��xr�e���#��E�W�Ϡ�ȴ��X�[����x�w+ԇNxBLa�3Oa�i�X���$�{�}?�	- ������J�ig[��#epdU��ʪ�eAֆ��-P�9ޯ�	��q-�����<�����b�A��������ti�]DXq`W�O��C}E��O��)�Rή\�I�L܍�R�ƾj����A�3%w�q�@�|�q졙��	w��� z�R��� ��s��o��p�Ղ�Un�lL�Q3�A�Z\��Ҏ��m�� ژI��D/�P�v�2��X��6���P�s�-�/V%_���� ����9�k��#)6g¨Y�k�t�����Ǫ_p-����~E[� �H:����:����c�#���H�h2[%'GÉw=�!߃�c�:�k*��mUd��5_ɭ��Z��N��G�?d-?‵d��s��)K�Lޫs΋�Y��C������O��� ��c�������b7汄��NxO$-�.�i�
���k��>���코�9��A�j�N���1:pa���N�Hۂ֥�v�ʆ���K����ܭ��^_�F���_v�Y'�wԿFe��Uj	�1����;z��i��S��Y_��RpŽ����9�EX�͢�S��`���N�=M�ԉ[d��,@a��	X� Z��`0�7��(���-å). ��P���`���{�*���������1���]�U��hI�!e��JO�_*��S����� �wG�9EV��|���Q^��H�Bfߎ�!x�6�����7Ήs(F����-�R�Y��Y	\G��~ܐ�p�u�N�#����Ʋ`�2O�=�ݜ^Ɗ_�����&}�d�����W�^pg2%ǧ�(�"��r����?��W�`������֦����'!
�E�s�f�-HH8�Y���K����c�#��0���}�|�(A��~OuL���q���I85p�6Q�	w��v�a䥰�{븺�T�|E�&��ΫISl�h�>�F�ء싄�y�X��D ]�_��.�.�D�8N �o��2!�5 A�-���.�ȸqi^H����=�UI�:qyH+���C�Ig]��,�\�)}�i/��n���2gm��.C���$�Xg:��o�HwMn��2w��bg���c���:}j�����/�_�-�j���0;E��{DJ��h��ô��ʀҼ��0xF������)UqFM�.
ސ��g�� r��?���}{aX��(0`�7]`%�B��D��\�G�2�,O�%�����wv�l^��t�����4��pX�Wm���f�:�3�� ���8?2y�����i%Ԃ.e��.j�����(�0���kƇ"� %�o�/�=*	���b�A��'��!���U8�Ulk�������^�E��~��z ����F�e-<�ICpV���-��둡�𶄈�pu4��?��]��L[��,~��n9�4�ul@��z�xtD:6!K�
݉��]�;�[���@=z�(>I=K*��0��˒~�����cl��P��n��u��Ѓ�����T�fi5��=�8�3^Z>S�Z�k�ϒ�H�ݱ�B??"�?'X���뼵�ߖ�'$��5i��ȣs���	�>��2Y$���_�x�O�>8"5E��T��}hm�^�7M���Yp`��m�
��|���@ג����)�K�6|��\�T�	V���g���y p���]xr���D5�#9�>�5v�O�1�6��Q�@9rrIc��f�����ox��]>��$���>	�5W#��l+yL^��:*�?B��E0�=�
���	�3+����B.9��9n�O�}��;�#Ѓ->��g��[m�Vs���X�]����T,��z�_@{
�}��DBt/l�S��[�$�b��
�!1��a�p�K���%��d)�ѩLl��S(��f^{2*"��
 s�$ֶ�a"a�-ų�`@�I u����x�j���o�%P;��ṿC�
��܆����2��� df77��9�UL�]��v*D��&D�_h��� ):5/��2��h��!���,
���������elG�p_i�L�[:��Q����a��=r�1{%�O�Ծ"�����E���ǽ��8��?w֟W�P���������I'�n2jU�Ϳ!S���ZHe�H��q_E�1ME��Z�3#g����1��LE�zo%"n�d��Ә�fBj�3�~�.��3�EEa8���y}��b���D*oaä/<��X;?LRX����M$)
D-�s�~������~':���O��<�f�bKJ����t���~�w�ҠEf�|T/����	�Xl�R��q���sT�w���a�������\-hT�\n���!1|;��5:�n�J-~v�k�pҁsJ��0އua4��b����H�O}�&���j�F1�[��AR��X��/>���⬓������s	��S?"j\^�%�'s~� A6��H^�C��9��>�}#���S�Ü!EBv�0�~�ٺJ��̕v�u�/�a�G��]/��@I������H�7�Rm]���*���{�u��s�Е�<FS#��hZ8XB�W�8��#���b{��N��і��UL+ݕ`޻�i&�1jV!���`���!=�B,R�A��I&�`p�hze�o����� ��TTZ-��Qݬ(y7)v��J7Ђ�,�ΣK���,�NV����Y������i��֡/nQ0͢����ĲYI"�J�.^I
�4�[I.c��T-�9�V�fCxd�=�U�L��;����M3�N�^K���5���Ua/�`HXs/�����-
��W��%N���)����!�wv6#L�q'���&jq��>�
�bRDa���?����_W!��rT�<E�<��� ���!�'�g��:0��u0�
��*P+�d�7ԗ�����z��R�).x����LH5�i�~ߺ�)�>�\w;AW'Ӿ:�н�3z���Pдw�,����S��p*�h,�~���R���?LB7:��i�q��k�����]s�T]�@P{g��]ͨH����KD�7"G�|D�NՔSn37K�?@�=`
��^���6���'v�V��_5��j���򣱪����,���@�-�
�$�U܈]�8Bd��ѥ�S��-�q[����"t�X�]Em&u��opԵ��`��?m�OcWk;�]����]�Q��ŷw�w���r-#"���w������	�뿌Ϋ�I��ã�S}84�fM�iy�S�؋���=tü��P �}��=0|��)��?��c��A��8���}�7n�r��Ή���.���,*�Dg�
��%�"o�������K�~|HA��s�>q�J��p<�&�F&�+H�e�܍��ܣ��'/.�#� �����ȯ�W���'�� �T#4��3}��P�?���ͷQ'48�*�;�����Y��pԚ
�rH��+�>�~t���#*���$e�xj<��u�d�.����^����4�*7����lv4�+��Q>�OL4����r���r4���^�oXJ�÷d�yDC]����U��o��!���]֦M��
g�����68�T:'�p����ؠ��k�&�jA�4yl�KC9������ڜ���k�S\z'�4oWFWËւkc0M�ب`�z����U��6r�}��Lw��	�%"�$=X��o6~-m��X�q��r���Zu�tP#Ӥ8���p3����ã����ӞY@���j�6�	�v+tFgY�_m�� �ɱ:^�H�?�e=�Z\�����3�4�����jƠoS���M(��Nw��B��3=�3� �8E;�3L[�G��F�;��!xM�)�w�_ԩRQ_A���~�m3S��`����R}"����Pj�,�� �:��\�����;Ր�+��TwXyz��j�@�h�tM��O��ͺ���M��xf�nQ2ћ�s<�$l��aK�5+�=�3�&&5x@� (4�j��$��[: l�ioL'�>���4�����6�����Sg��K����$���"�	9��O� !�ՈгP�&�>M�]�����G�\7��N.D�ث�f���#b`�K�%�&�(��v/\;g�	�&n�0<SZ��y=�_���3NjǾ�R�P�+nU;Awsk$B�����7*��(�Ld	G���c�ǲ��DtM��H{S4����%N���XF�tP�o��)�{j���5��DD�6h��*�%;�����ՙ��1'd��m�.W������q�e��y
��D.g������F������G�E����l I��m	��3' �S�w���N�YT�פ�-H���B�Z�@_�hԶk�j�R�˝�X:Z(=�IK{���ˈ�j�`����(�@"��&��:�e�e�i*��Ѻ� u~��)����3'����0k��+r�̛�6ط7�uUKz��oXri�-8 v�����ߍE��<��b������m���^�)�@n���4<�=r�ȍ�0��1��6{��}���=�S7�yģ�P}C�+��a�
���Ǹ�^�rJZ�d��\Q,zǭ3�j �JmJ	{�x����.��g.}\ÚhZ�'zs*h�������QE�m�N�t����G�/i�0�K܃ڰ�� <��ţ	x�]���G�L�!�Ŕ��_|��M�L���l.�Z����%㼔�&�h��	&P�LI�f���R�а��Q�i<��Q^��~���a��7?QtOX^��)S�C��^�Ok��.�A�:������{�i�E��K�fń��muP�qj�)����8!��n��mr67��_h�?��t�{q��.h3�;
b���-]��0�g��&�R=�K|���.����wt�¹�1`�,�/�_.lTi� 	��wk��)ҋ�����3������j�s��cc�.R-�)C�ev�ݢ�sP�SU
(��}�?��4�drD;�m@N�B�S�����t?A��t?�|�<$����G�9(�e'׵�>��� S
�:c�0���vu�C�xVω:�8}}k�zk�$��욄Otd�>�����6��U:+��L��Z��ߚ;H�2�-��ۢ���*���'�֮k��:��`��N��S$J��X{~r�Ƥ�����8IܻH.��F~ :e�\�T.`J��o��^���<Ya�~����^�2�<?�e5��U���T���'y+�=ET�EEy.���ؽ[c��X�y�짍)y"k�}��B \��`E��K�;�˃~�#�MO���U�t)�_�H�dG	���-3[ZUѮ�P��"�+ɒmٰ�<�6�(���]ێ+
`��X �]�u����}t�og�,ϑ��z\�vg,bP"[ �t��u��8z����j1�6�+�m"��jC�L1�0��I
�n*rM��$�eT���ޛ�$�Q�r��
+}��M�z���R�p�����&FrX��s4��i�Zjy������'F؅,��P��M.�ȥ
>��Jh��3h2���g&2�F���|+^��4�K��+a&�%+��UI�"*_�h�]�6���bK�FblU�]V$��l��!��N{�w���M������88���PA�7N�Sx�g�5�iWvt'�����˅0�V��u�2U�Q�t��E��.x�{=;��j?~0<Z�j��nwy�د=\V�nS6h�-�X����6��r+����ʻ�G�0�E=���2w$F@��cU;���[��Z~T��b��Uɸƴ^]��8��#`���
c�Y��M���q�1�6�²>�/3�L��f�зDmI��'��i����shnS=��|�=�M���s��e������F�������Q�~�J:Dp���5��ؓ��?T�`5���(cL�h8�x9yREVޣH���ƥ}��l�����!XdP�,T�V|�g?�K� E��mKR[�klX�3��A	�Y�+NG�6=r���.J�e6����+-b����:�Lu��
*+�ioY
C]�!'��� �$��h������ V��S�� Vٮ���ύxUr7n j'��L��Gs����&t7%|M>��>`�{^�������1'�w�dw8�֟"L���Q(3:�|�ZO]�qM�L%}Zx���,��CN}[,$�"����*!��ٵ9Ќ������"��:�$�
���r��q����������VB]��X�����㟟���7��iW�Y؟5��U����+��w��Y*"B�m`Srj�����C_������٦\!�6�Bg_9 �78��5�k���g�8��6���m�W�-���*Kܵ䥃��-�����������M>���_@>��6W�9��L����]�xhl�ԭ���	[���F�0������O���D��>�"�_�f
�i���R:���{b������6�����-a)�%����IKp��9{d��spY�J̸�G��ws��f]�K���"k�^�e�|��?�J�� ��S��.oP��5�Qg���$A�1��g6�Q�ؑn�ySK�'5��S��z"bi��RB�&�����?��w����R��e!�ԕd_m,�?�(�����ʸ^�;�&��R�-"Aя���s�paz2�Lu�ğ�z^�U2'?�@��OِL��U��t���I�)�i�?E@����Y�C0Ju��d��q U����:`�vY��/p�?�=�?	D �^.�����._#ؒ���[`؆�H�i�B�M��.,�Q��q�&`|�� ����wZ��bE)�lqEQ}�q�[��#��V��,��������K��[=_��fsb�dB�3[T����o��Y��(�gr��Oڽ(!���^U�4�a-�����j���Y;�1k��_E���dD��m\,�_A��4�T����G(�8�0i{� ��-� o/�����p���Z2��i��b.z�"1������	6��"��>Y�r)�e�Ӂ �-����Lȼc|:N���f�����Ua���G)���z���T��]H����5d%]����
ljT���Y�Tp�8�5ɵ0�XQaO��q�G�-��͠�K�k�P�~��sZ&'(�< �$��k�r㠰�[�`��
�]���P7��!r.L��%�O�H�����xs{�	�E[�v �����p��CU�.��y���yL׺�Y|���͋q����g�1΄
E��)��fj2�xY�U�=3�B�-C@Wb �{C)�rx����m�e3����N,�5ي�������{��}D�N.�>)��x�[�_�h�aZ�\���A�q�i!I��Y1�K�}O�K�D�������bkU��2}8���@�	�e�PJ?:�m"�bK��.�Y+�\mZ1��v*2S��6�ӀC�m�+XG>���Z�&T�jE��
���xh�da@��U(��C�	Ԛ���%��,Cw���'���vSt� !w� �W��c��M1D�H�ʍM\4[��H�Hp]f,���ٕ�i�啻᙭lu�4�6��.E{������ZU� ����*u���L�R�j�H-�{L��z4�X����!�]9&���m�ӫ�4�r���7̤��.��k��8�B+qEkwD��O>T��L��02��5��h���>~�E�h�����+�{���=��ɴ��+��2#�0��/����)l����d���m���fs��M ��"� ����ˇ��6���áCn^5���\w�9M\����b��xph@�k�s�@2aSZ��6�&t���pu�[�nm#cֺ@{��-F�8ψ@��o�F��9ʺ#=��	B�vҕ���.�����|JG�o֭Hy�� 
aŽ,빕��.�b�v����<>�w�[�y?O�}+pd_< �Sa����&�ܵ�A���n7�,hZi��+ͼ@�[��~oR�jt��P	��<Ha�
�ہf����w����j���ѳI�E\H��"Zc�7��^�ȳq�Z��	H6�(�J�/EEއ���
$sЯ75f�������ܣ��|]szxu���k���Z�)v����5�����e�vlx�0�7��D��Y��@!>S����,_$���������z,�K�ј��_!Q#����B��i�t��cQ���XL������؆��A���m���0`������6-��ݰ��E�Mƺ�3�W����[����`hh~���\S4�ZbCx���_Oj
��Y�<Y���=b*�N����;"o��wq�'v/6&'oz���w����j��Dv�������T��P��O�߈����]�A�5޾唵�o��� �>�[7���4���N	D%��&����?��ZN2���G�_�n͠ޫ����3���/˯#!VcX0����h��	j�.��aJqO��M�.���ѝ���8&���N�rq�C�p�ܚj�U�vӫ5��X^���@8�U�G �g���hB� �@?��+41[C�a�^�U�y��^�R7Qs��	SX�U�����g�e�:���#�������U�k1�6 ��#mpU��r(;�|o�˵��5Tl�P{Ɩ>������ ku7f��{tE�;/�uϵd0{��9��D=,L�VY��C�Wq�=(/�к��}���g�s=wVp��8�ɫ�;�%5{�Y,KQo��uuy-}��ҿ����[K��9��I�_��F��gDy{��pG�i+ŝ�,�FGB,h�7Ŗ �� �i��7|�!�0VC�-:�F�uڰcRf�qZ���acJ��$~���l��Sb�Jϟ�UН�i����G���X�X�>�f{�>F�`�j"[[{��;,;t-'7n��K��j��.�@���ֳ�0�*-��1��=,��X�n��J�K苐�_�DB�V�n.V���y�E�5���"�z0�%A&X@x�-�\1߀�i�ㅔ0�
c+k5�7<'���w?6_>Il�Z�Z��DlѺ6I|a\^9@S��5&�,[u�c�b�c�@�� ybSj��*�S�F�����¼�꜋��[ٓY-����L��?#f���s�sB�=��F,c�:����^*B4�V��[�e��3�NI1�h�R$�T^Pq�% |o[�����n.��܂2�&���䓗^qd9�뤔K{/A��b�-\>�3�B ���Q�x�#T�g�߱���֏o�D�]��:$*	Y��p�ڙ`7d�U���)�+cH�;o�#!
��[�FFi��z	�w�1	1�c�����#6�7ж�}��^fzVl���G�%���Z��@�鸒X���vq�HtB�XJ>]d��V�,h�ډ:�p�h�u�+�%�60�cba���^6R撥��%>u=+NQ �|Qq���%�v��R�%�,�yJR��bK$R�=��"ɿ��%���u"�-��b�փ�8:�����yD���j�D��*r�K�f��AM����M���բ�h~�.Vz�z��� �P������=��V|�~���ލ&�U>S�'�Z>o.��\�s�O�W>D\P=ZN�^8�ܟ���L�}a�ȡ
L̶��:z���I�3kИ4M��\�my��MӇ�P���'��^�)
�����g~��ۈͦ�xG��x��km�݂@h��d�y��cƠ�[Uq8z�L�`.�r6;9��d�h��lngqBp��a��;�7n�rS��j2��Qc���_r
����Q�.�����a�7�+��mͿbɤ�z��b�%���TnV9+����e�`L� ?�Fk��*YH[�x��۷N�nQ5�I�58���JP�ER�`�Mb��F����c!�>�h�$�"�;l���·��Z1�u#8SW�"Sf���6y����I3��ɀ����nʨ���L[M=|�!��v�������xh��:��'���J�'K�8+�x��]N���y�p0?�i3!��{�=�-��K|�k����/�n�͉�#G��\�+z�|��u��D�o�������9�`�:\q��<ohC��	H/5�L��@�T��0�c����h���K7���Gk""���:41X��4-w�K�>*13b3��}�i���z<������0�8T����IG滢P�E�fm��r�=[P���ɜ-k�5�����-��O�d���M���c�2��,���hd��f;g��\��w�R�-�tdQ��|�
5q+!Ԛ�J���j�;#i�%�Bvhe��P��r(^�}O&A.�h�5�ب�`9���+{��������L+Ԯ�@��|D!��a�eYM�; �L ����\�?�~-������SQ���v2-ۯ��h��5j�Y(���|I[`��t��>���]���H���]��_i���e-73����T
<D����\C,�QPJ���� E;g�.殗��,Y���w�cH��2y�n�?��BͿ ���íN� n�L�9O��̳��y+G;�Y��kHE������=m"םf I�N��}.퉍��5�%ճ�f��A�	�n�i��	 �L��b/_n��
U+w�6�'��/;3-�$��?�ob����?��|i(oCed?�7� F�	]��y���b��[��%h���keX�Z���L���y��� �ϔ���U&����|mwe�~-��nL�}*���y�Kk.��^�a��f�*���E7�X8���aQ�,�o ��vӂ8\���Q6 �{���������Jp��Lw�Y�3��1�ėd�h�`�l-/&��t�R���[QG�r���]������xh�~X��	m���y�v�_�ᘺ3�B�U����e���v; �'����F�����g7"�	��L딸�Ѡ�2�ˠi˼a)���?=��;r6JGG�g�	\P�)\iRK�LU"κ��#Ѩ�L��H�R���W0E}����G����%���&B��������!/-{����������o��bOs�m*��b<��/�18��>Jn�����?Yr4x�($e�r|>�����0!�k����
���rX�w��v�lj�;c���N�[F��;Ù�+�.] S���x'���Qb�p:����"_�&`��s�MF��q�gT�2��m?e�Z��Xq�8�Nz�a�����1ѯ{`_������_7;������Q	
m�I�F	�M�.���j� ��u�����ؚ����o�8���܉C�!�u�o	�h�>��|Mv�NZ�eG�0fFY�F� �FA���u����}g�=�B�(-%��њ�ȸ�It����|��P�&�%<_��'l�+P��� VuW���Lr%���,x*�&�`��P�"�6����E�weg?�+��Z�3I�i���o�^*�9����IW#�o���\�k�N �k��F��WD�GfB�aB�R7�QM�J���,Cz�j�'�]��3߳���B��K2��VH�~���+�j��jzH,��i_���iD���N }5c�rF�㕫���i���q��"�c�ق1���w
;�g@M>�s��TXbr�s��~o��<�;��tEHz�x��T4H���]99�A��ʅabg`-���#�c���C4Gp%�ف�/v&L/`7��m jNkN�7�+2N_g��e'k������yZ����tc`��Y���j�`��FOHFߩP��u�J}�!�pX��[�Ag�X�+���������.�Z��C�:F���D�葚"�i����	��7!`���H(��
��Ѕ��l�F���0)�b�+	@�j��nw��d�AG�g�� ��A�~�Cd�s����
�k&Ш�#9i��Űٿ?�2$������*�e��;g')�72��sm���ԕQ���:޲�9�:T���!��3�9�_����@_k5�5&D�Y��+�[;A&�*�ɐ��p�Q�v�G	b��%?�0�%
S_�:��98����h��/yqʉ=�K�յt&9Ә�ˆ�iH�ڀ���1�4-��beSF�·�
xsf�eYs{�nѺZ*��Zd������Ӧ�!�Ց�ߤ�a���4�T PIC!i��.Ջ�l��<���Zq<��4�Iy1D`u��1���1�\:���g[g��������V_Ew`���G�]�S�پD
Gv;Zj3��<��r�6s�(�mc�tHR:�C����B	�T,`���1�&�}����!�I&R��%�����FX�,�ə�m�o��$�)�6���E�(�`Q@�17���2�">KE+S-�~�t?U��J��S��e�N�X���}4�C�Z��g\l���뇏�,�������Yƈ6���ɵ��;�M�oN��6xUڏh=��@ai)]V�YUm /��jz��lsg�S� ���(8���\]?��&HQ"�n�3;i�)]�\����҄�6�s���� �u9v9K"G�V^�XEN)`K�� |]�?�@�PJ��R�Ď�R����-7�������Wn��gzPE����s&�y�?�>�R��_�C?8-/a w.��q�<��X1g���.w���4����=&�l���˸s�\�jk��^v?�z�M�U�l����{O0��ō<��}����G(����uKZ���B|�����)g�����Ϯ�ZV�~ٞ�g��Fw��^M�q&��l��u��B�2�9��L��C�r��=�/������(��R�LO���%�k���׏zڻ94�٬��'-��c;+�#� S(�n`��л��)���B�/�I.��]	��A��FdQ�zT`ҸWO���^I&�y��M�p��5��jl�|����6l�ϊ1�U`�J�k�L��AC'}����Ln� ������LCy�c �~�I�}>>_vV��[Z��__̹��5�
�w�Y�k�Թ����ǩ:�*́�{�z�dt�-K����i�%%mͲ_����S|Y=۾R��H�e�\�ʳ���6@��
r����Z��l�
c�*V�O7QrFn��ռdR�T ��j��9�.���3�_F�V�X���=k�J�\YvfǙ�z�t'�v��Q�	䝯�0��O)Dί~�_�i�KޒO���+�^�����:�AUx,�� QC�V"C���Z��]�X.���6TS��@+�o��Т�`B��ΰ���I��x4�"�鲶��N�{����x��(H�)4~Ǹ�(�5A^�E?y�gJYB
����R��pτr >q-m�MFs�7��T��yT"\U���p��O��]_���3�~�1FU��	��+���Vױ���๋u��as�C�i�Z���]u�'�����"D�f����{B�Sp8��''C�X��<d3�HR# l�����&ˬ���tm��`�,~�����b�O�\��V`[��0g(7<����9�OD��-��&��"��3Tţu�}̉U��WKA��F�X�x�rBp]����g2 6�~Fs:5f�Y�F/��љ�z2��x�燧b�JϽ�4�Wt4���K����gݵ�7z{P�U@3�{l�)L�LO�L������� ���q+�Lu�����EҲR�x���<P� ��1��N
�f���*�|�<��7�)�����N}���]pT������4��*\��X�ZǐJ�? 
���cg�.� �7�B�Ҝ�,�(OϪ������e��_6������3�7!������ǰ��f�-�ڙxӄ�,q���@-���k�]+��QE��s�-�"ެ���9/��g^�Ã���9�Z��V
١	��'��������=���%��@MY��j�6.Vr���t�u{��5�������\��/��Ȋ ��3"�nnka�⃶�^>�ͮڗ�� j�����аlep(��q�vx�	�u�� ������������8�xZ<��UjL$Y�_��O�Ӳ�,�"���
Oɔ*��<��.��,[ r����E0�� O�ʒ�������ZXZ���N���H���M�`<�C�^��&���b�>w鈲��SI�"���n!��'Ɋ��O >R	x�J�ѩ�S��qѳ�
��q�o�[r�ƅr�0y��bޑ�9,�ȪQ�=uUa��D��Q����s�Bs�f����Όz������ f���TJ��_��T��F�u�/X��[��B�5��#ګ�}�N�?�{�뛹䌍���<o�<�NGQ��
}��MUT��X]�ဦ?i@���<4�����Uu�+E|�`�kHY�<f�vK�[_OCq�u�@q��
�9B<����u�K�~7N>)�]�Yݵf�~��D@�~�g>|0@l�A���m~Jo��d�%.��y�3Q^I����Md�%cb���q�7��3��<�:��=�������I3����<"�[�K�.���ֱ�H�?�MY 2��Qu��<����m�d�[.����-lsR=�k>�ɓ���.�p�gĭ�$qa��7�(��h]R��n�Ny�ƶH/�[�,�1�j.D��=��FM�%���a�@�RoN�6�����0�+�df]�57�p5��=e�iΛx*���c5l7��[�8��z�O�5��ִ���j���y|��	-c':�lG�b���n��4� C��dy[FV�aYhտݱ���G���.��L�\�R!�c�e1��fod�3 Sy���E�oP.qd�p*���#�g�Q�`�T�����,ѝ	0������b:�Q_;)��S�s�3ϦS~�uTߵ�� �XB���c#3��g��1�6�;�)������yYj<PhA	�[!Ťh��l����*���PȐ^X��ؔ�R�����w���}��Y�Hc��4ʣ�!
��aD�-Ӯ�G&����RP�5f��$▘Qj��)�{�O!>�𴋄3��(}(�ϔO�˛��4�+jQ��܋f�

�V'��t���U��+j�n��2��\?�.f&g��W�� ���/�F���ǽ2�U��M9���#�"�ALq;�g��b/�b|rd��G��b�����F]E��8�h��Yt���c'���B��l�� J��Ɋ\4A#�Wl�k�3��شI!��C�A��&�Y���M=���0ȫ	�[�1�sn��� �<gP���h0������"hѠ��,�1ހ��$1*�Z��wf|�c���52����`�h�e� �7�����T���!�1F\�-�]�m�S����$B�X���Q�]Y=L�* ���&�n_����6.�Ww�Jb-]�U�\�<�{k�ͳ�?�/V�ဎ��G��e�����J�x��ׇBeF���K�w�ĝBV�B��̷��F�lFW����3���-ɮY�f�d��;�
���Y�uǹ�(�_7�=D�l̊��2�{�T̨;��Xp��Q��K��Cm%P���y�Q���f[N8�{G���[�AZ;���7�z,`�A�&H'�l�n¥�ʏ{��Az���.j��	Y�{�4d�G]Qbr�d���̹͗��I���K_L��z�4W�|v���M��[�2U���q�E8W�Қ4/@"���3��R����ؠЏjLkf6��9�&�������A�VQ@/�?[K�Ļ���%/�佘��f+HL|�d�E��ޯ�i���
��[�t?�"3����d� D#��_ׅ������n4��-���1�%���E�P#M��D���f�5�wR+�����Oc��$�:RZj��
�M�8iw���O?�@)'3� ��p�08�96��Wj=�ˮ۟қ ��.`ȫ�{J�Q�a�V&ϖ$У�}w{�zuw�j���ĬUe�e���s 3�M"fe~�Eo-�uaZLU� :�0�}����T�v��Cg��ӑF�:�"��@1���ܻ(4��b���E��7�"��M�{��[�R��ptc�����[^{�4���x!\�ŉBpa׮ӱa�9�,���5�j�b�B���%R=՞J{�#�:�R�j@2���Ӷǈ_�%s�?��+{��j� �@��6�\su��T^W�֊U��5�����ǜok�k=&�,T��+- ט�oKSm���O�B:+�|��X>�F����+�[���ݨ7����L�Y��.�>.g� |�����#rn	���b�I
�#ߣǭm[=H�}���p���7Q�y�s�^�^��C�ʬ{��mt�þk3�n�֮�5kl��W�[�Μ�2~��� �W�6��j K&(���""��?�;��#�s����gS4}���?��/�8s2+�~ߗUѦ��A]y����~��s��й?��K#dpᚙ�Z�:�I��nJ'vc����Ck�z��qH���������&N�2V[���w�}�Q�f��~���o�#����Z�(%��'�).!����¼��EvOAư�0��f������]���ִA{J�����$�TZ֌U�ugI�<����W.��}$,r���S���E��NU���w�� W�ѫ**hf�k; 8e���92�,���t��c��w[�.����"�%�}��]A��c�9��]��(O��ƿۜ�JQ̝����`W�'�\�^�ߧ�S�Mp���#o���OV�\�j�̣N�{�lQ�M.3����/<�l���F��d���i�X��u�v�-��&�����v�J��Yx"I�cnb�2tw�W��H�#t���is��=��[p�g�`g�YխOUv(�NH�K�9���R�|D�߰*��Ʃ{�*��=|IOP4
�Yw�C����m�e�� �x$)���~�S���,C���=w)n�TK��o~Vh8��4����%�e��d�����m�ߢW��U8G��y��3T��<���∻ч:)� ��,e���Z�Z�U/�#?"��\�5=��o��]�U�I$A�N�S����@2��H	N'O�tt�޽"ʝ�XD�^M�-4Y�J	H��ʣ��ǜy��wy�P��*���s.�ƩkV���0/j�$R^[����5њ.�7I�]�W��rM�����y�1�@|��y�ތP4ً���}�J� ���W�о4W'�����ʌ�J�ף�@���4��2艸f��Ќ�K�O"�G�%fS���0n�ƚO���1D]Ф��ʨ�k�K[�����t���=�o�٥�"m�򜀖�=��B���8��p��Z^�:�{��.;䣟-.���G�����ƭ��2Ćd���k�6�g+Y�V�_z("�s�+I�O1��u�D=��R�\Ӂ_*� �7C�pӗ�@�۔ֽ6]բ��=�̙��	�����F�O��.7.r�܊R�Gc/Z��n�e�'Om
N6Q��({$Sh5��F"�<�#*M��4��d�'�A]P�����h��8

��ք0�W�K[Plzf�.�ڙK��FrW�Aw6O�<��V����X�R�c��G���M=J)ֵ�Y�����j�H�>��U�����IT���4������+�����)�ݣ��gM�Q\�>Ax�U�7�i�^\ک�+��������2�+��Cͭ/'K|IJH��}���|��(ͭ; �M[�𯙎���%F����M
�L��(�l$i��Vz�~{�˙�i��M�nn����=�F�>�����dS���]���ߕ�J�p��9�J#'v���>)���i��u6cH���>����!�^y��i���-G���2���g=��m@,h�ֶ���!�;3�-!��f�Oq��W��J%-�')��c������[|��b����bG�F=
N�� ����w�Y��Ɣ\�f�j�[$9u� _\��?�5i*��{!i�l�fuܕQ�~lTz诲�U�9��>w����y�]�Llѻ�њ�0,��&.��5qa!t�[H���`nf�[�՗�IpX�u�	r��B�0��iM�B�{KA�FG�:M+hΨ ��ŷ<'*���z�@��NWOFhc���{�������V�2/W�`��D��2���Ũ~t�a^ѷ��w�2 �����?4�����bb�h�������;*�@nP�����Y���!؃���ӂA�b[�mb��k`�QpEn�s�:�^��tP1�l�ͳ�F̆�ѽ��"3l>���`y�I�)a��v~���s�ƺ�f��h�g���@�N�FV.Iڔ��o��X=3���SR��R?�L�*���G��#��5n<������^�?���e	E�����J��eA ��k�?����g������Pmwo��TXć3�J���NozoUk�́��
�$Ko`��K�}���H���J��$�-5���Lh(4_�Ah}�i�i�����?��:��m� �l��H%g	���=���ѭ"�	Xb��p�yћM�R~ӥV:�iaӠ�F���9��|e?�P�:�d���a����_f�yP�9Á=B|��t�k�ߤ�v���WbD;�s��n�'�H� �3�U��M������W���T?I�A��̎�5�Y�v�k�
��V��
��U�_�J��N4n �q)I��V�nEΉ∰�hó�S4I*��l��G�%��Ed�;��n�y�-A�HmJW�pg[�5�.��Nn_��,�����"����P�9�孱|y��^�-e���FO�t��^��it�+�!"XZ���a��Y�cN��%�i������k<#6���ȕ>��=�U��4Y�$�+�I�O�ܼ?\�)���*D;��c�����Ga��}:��l��1����>�e(IOĩ !+���U"�sxm���9R KL8�lڇ���z�:��jm�>>�V�6�+�O���g��~D]���ژ�`��ň��|$�9�+ГuU��*e�H������M��<��f�4�0(���i�٠�����>��{>(}��	�r���ge�M+i����j�*��6�r9����i^�w�mB�06z�SYUD;�g���]�3�՛�QÊ����@I1��M'˄.eeV@��b������בE�,ȿ����%��h���.��l�F��}����{K������!��@Q�O�b�d��W��e.z�*�һ	�}�\?t9�t�߱��K���AkxG�(~줡��~�Z[@���E��]�T.[3FM���3R��ݬ�fb-8��p&����zX�?�{��`×��B�[�����7��zXD@8�S��av*�U�m�J�����|_j;.<G�s�܆��s��-?޿�خdѡ�(�
�?��f��Lo�s�Ke��i�n�o�/ƭ��2���^�!2�&�ڢ�/1�uL0���?��X�E�G F�}���b�	XZ����j����Ź�p�[L�cf��)�&��-�p�rZ'��]!��vv���	bW��Dnw3�K�nH��3�&~��ʟ��P�k@�Z���Z��uR0o-��U��I����
]k��>dV.��^�rwWŕ�T���Nq�6Q
=��[�և�k��Tp˺\E���X������1�F����I�=�y{�q�#�|{�=갪%O�2��W����Tn����CEbs69%�c=I�A�eٙ�R�� ���p�H��:.q��r|��r����x�*�R�x���'����#��oU��Ɲ��%c�`/�dX�NƇ��UYh�u@]i�a߲X��=_���pӵiL'R�#����p,��,�dz��P�)�����Q�F���)]0

/!^j��Y։�@}�V��؎DS��h�4�MRtb�G�u�#>/�9,>�̚��v{PV��>j��+t�[��yS�?Z��r�(�e��m��3Gt0(AC���X���
�l/��ݙCP-�.�:���PR�h�A�_i	 ��/U�k=��(#-�/�y��g���-����Z:ȁ'��F�\1<{ i���wlO�ܰ>�ݎ�U�p��#n�͇�~ 	Yԭ,nߔo����m�Ø�9�)���p���:Ş��i��۟�U���
��l	F���Z|^n c�-!lf5�o�Ζ��[������}��6@�Jg�x�~��F�k����	����P������ۏ�fd,��TFv?@]#�����!e�1č8��3���~@Hr}pT7ft>�\���R�?,�ⵣ�1�B�ݛ����s=.3��U��i�)����m-Q��3"X4T�}�����:�������G?|�x�����$}��qr�W{�-�("�l	�aV��D$�eP�-��K,U��3��&.��piL�aZ�
�AF�e��>��qj������p��c�$�?��n�J�),� y�%�=�����ʒ���Q�2٫=0�L��_�ly�T�o�sao��6��.�$�J�%~��f�ܴ�� k_�7���Ȏ���XdM�ud<�E���8~=w�9$ֈ\r�^	�8�nYjv~�F��5R������	p�N�󓾓b��q�i��x!��7�\`����F"�e�����D�?�Az���k%S	m�j�����[� xA}ܔ�'jLj�=�%����`�dZh�s��47h2�Ycm����-E1-�)Q �o�U�	P	�\�$⴩"��O����̍�����Mg���}[�eZO���n����L������ry)/�.�ԝ`�����RG�n��[M����&0�$�T	�ﻮ�j��k�.����\r�47�_��0���=��կ�^��^;�G������ViO�[��ؔĘ�k�Y�*v$V������9���?`bX�D�,�������LK�dn~@7,Ѳ-��ztc�$A��!���0��:�S[͌��@���n��a��?��XM���:Mu,N�Ӭ향��i�5#*����U���K���;$���"�������!B�7�[�@�ǥٿ����om�Gg����u~R�5L��Z����BN0$�f� _LAJ�N�m�!�7UA����U޽))r{u��X���gT��������I�#Vb�{�8�LQiq�C����&8���Q�M�El�N�5���R
��W%n����r��^R�c�~٫�<��6u$��]�������2�����\�tY�~����^iO_�84�q�Բ�mW���ikh�B�9����R��+N�'f�Դ��1חp[m�kh�{c��l�0B$s ���'x����Yy��l(������M�+5��4�MMA��m��_(�¦QY��-��e I_��:+a�r�d���3G���:r�U �5Թ]/0H9Kk:�7^�nbc�����Q@7�HH��AN��2�m`f�Z}�LZr�y305;:�Y3e��Th)~qW^���%y��g���֤7J������#$��=�i;z�-C�{go�Z���E=H�Zdf�u=;���[j"���e�K�bt���.�N�~�o����V�b�7�QO�[.B�5�]�dm���ǃ+���
�i�$
����q�I�Eӝ�(���l'c\Q�F�RC`Pi�	��ZV�+Q��0ύ����Ժ��Q���If��*�����`^��r�@c+��:qR�E@�S�٫�%����<��$4(S�`㾪h�r��W�������.Y�y��]���rZ���Uf��J�1�5$�l��g�pT� ����&+H�$��r�x!�D��%-���=�ϊ48�����o��i3"-(��u:��o?�J�c�t*�uj�F�L��0� O��� E�����ԐN�A��
T�3!�1�Hך�֠���W�25��jE����v����HJ�mt)s��s�=�Ig:;0�!���k��e�L"���B_a��w`;�s�ےT�I(�S��V��e/?g��B� C:�=܊˓��J���)N�1t��`�7IRpz�
���ty����d%i�������wԄQ6�XT��U��d�JL�¼�xڂ��ͷ6��87����ݫ&X�UZJ���Kԉg ��oﮉ <5N)�lQ~��Ͻ�R?�\9�c>�KH3[6���v�~��+�޸7#J�+q\�Z�2��7�2��O��7��D�F��G�;��L!�2� �\8���xV�ˀ�~��SC�9�tQ|�hn�!Q
�D���p+�YޜB=S��}S���0��9��VY���B����\�<a�}��#�K�c��j@�Kˬ(�y�eO���O�q���{#lQ`[��H�zX3ѯ�ؓ�Б��?zð��&��T�L�s��ȇ[ޕ����$b+5N?gc�?�mE�M���J��"O�<4=t����Y�Yc�����&���捙���ހM�A,>ӣ<��%���+�]�PdR�˭�}��[��>�B��S�jܒ}�r9��gUS��6�л[$��o��	�~���l�_��r>�(���q��v�	����lSE>�����-y���<p�$3�"���i�~V��bb����"!�K(vn������s���h��"�->���Y,Z�ED�Y%6�+m:�^���r�yS>~��h��O��ɥ�r�?��6�������q�d���4e���¥ �����t�����T�eK .���U{M7�l{�lY񏀏�W��76��nq�%���*}D?o���Z�Y@��.�9�, Vb�fR�|�zC���2�C�p����4�k+�x����Z�s�v�:���(f%��D�&����Z�w�TdU$���pjQ��	�ԃv�=Jw�N��~��G7!�@ym�Km~�޿��N~Jq���މH-�X�R�4����eڮ�h���i�UMc���5$��K0��2Y1U|����!G��j���| >7�RR�[�����>O�G����9�Ȑ��4F*
��T�Q���$ɏ6J^�r?E�'���rqt2N|�@jj�¢\eL�n`a2�*��#�Q;7�XS)��{���;��$Sf�۫o�I�_�N]D�Z�嬧���ڗfNCQ&��P��[ONtڪ�?��+-)^�����ݓ�H�{ )]2.V�9���뜢h=Z����53��{�0rP<k�3�o�-��P������M��[6���QeY�����tQ�5bĹ([6�Rn�B�U�!J>	x����
�P���!�6�{m�1czф����@��LiG�*�R�`-6�=������#���npY��]D�e�@�AF�$ц�3B�-�w/�����C� d���|�3Y��~<oϻN;�@ko@fW�N=�R �;�x�5�̽��+D4�d�7�k0���L����Y����?�#~�.m؏��>�# f�k��qwj���-���G���ŋ,�ې*�ɧ�"w�.!$A��S��)�(��N��p�d�������$O6έ��눙aiuw0��D�1E��
6�xx���m9���	$'����1BO�C����e�T`�'࡙�0G(FP��wM�	f��Z� ����ܕ��Gdh0�$��� ��Ĳ�\���n�d�`G�2ֹ��-�i��H��o����qr7�y:�w{ ���N��+I�i� �]��,�N�W���\-+������N�>{�K�a`M��s�>���l�j@ہ(��M�����I�V�,R��P�2=��"�R0�8ȭ����R���;���Py����rƌ��X4�1�2�8���(NO�R�DAۻ���;���g��EKV�P;����#��L��S�E곌�x�ύ��?nv��U.���L'��ůc���hr*�S�O6��[LF��C0����%Ctu�[�/PA{7��{55���:f^ݎ�K��h�4��O}�;�&вɃu(��6S
("�B��D�O�]�r��F�"1�?[vTU�bP0Ft��� �P�M��A=�l�v�ѸxM�t�+½D#1����"fb�2����SS�	X)�G�ъ-ZL<��p4�*-�A&eܢ�e�N�vD��w^w��y��Q��BP#�^xޛ7�R@�e�e�<���L)t��iB���xZ\�AO�O����b-0��N`ڠʍ��#�Mi�Ņ���`��9��yF����T<d�^��Zsm<�/��^#�k9���d<�Z+����j.�n�p�SӸ�}D�/��o��ۦ�羣�Λ�W�k�Gw
��y�8������ڹ�V��7��=CJm��.l�|"5�[|�e����כ[�*,J1���"�-"��rP*qY^:�,g G���[��!g7�b2ml�yG{hT�����B=��Q~tq���ڳ���%%#�7�5_�#��9jd@�jt�R_�0��d�`{���.>������. ���rD��H�9e.-���c$,T�O��	���E�C��*qc�{Gr2��I ��B�ܙh=-�Q�A1�@'�
5�#��j㓉B02������(��vأ��d�c�k<��Y`|�O�^s�긋�ta����Y<��Pj�/�� dJ}���<ֲ���z�W�y�U��N������;m{͎�H(����Z�f�]evg�;d�| ��X�Q�6�8x�IV��[Ir�/�C^�ǖ�P(��G;����O�2��K<Í#� b��f��݅�:c���?s���$k��D�J��A/$��|����ˎ'���k���Uu�a֞���K���h�T��F�ӡ���e�����2 N����#Y�� V���a�jE0�G��/�j��K�Qu���_&YV������m5F�`�Q�Q�ވ����&����7>Ob]�����+wI ̯b���%sm6��@���%��(A�!f�� ud�����;m��-
h��� �1�EOÊ˔4�զ��w�$4*1F�)G����gFӎ���Mݪk��z]��|H�S'��QC$o��n��a?
�˦��!��R�($�g�S���vǗɚ��ԗP��%��2à̈7���v�0넀8Y��xr��V�#t����{�'�*�
�������?�k�dߊ��T=����Bi�K���+��.�^�ԜѷzF�P�J����:����J�� V�{"��s�����z�t�l������e�U��p�5�bf�ȸd�����,�%�l�cv�&�Ӈvi�? a}kkP6KY����z,�E������Я��m>��!���}����:I��1  }}�RKF�V\s�y�k��k �ф*; %��>p��r�� ŷ�%q9ƮR
(5�@���U��
@[}u�5z��]Q�7\^CC�[Ð|��8Q��G���#%c�u�N+��]�{��ю0�pQ]�N��f�����;5���X�+���)9��1�H�/�4$r�+�7P3_C*�R�*�3쓛᫏�]�&�����[%��Puޗ5���E�b8cf�U$)�pȰȋ��$#�/��O�T�_g�󄖟�t]�����yx�&J�@�/	��>e(meY��V4�$�*c�{�^����A�S"2�| 3W�����$Ҕ�������o	����VpȡA���NsҢ��9�L}�����ʓ"���D/2��ڽ���DXj�6��w3�)l*�=@|�����s�шl��)Eo6�x~'��&�Ö���=����;Հ�50H�8�S��}L=A�R��֩S��1gdO��h�V%@�~�ɔ~����tr�n&�ͣ���l��r$�%���:�h�3Ͼ�5=��Ђ�����m@��-�cϤ��lp�y:|t��h�� q�#�����{v�)�M)Ӻ�V)��]R��˂����E"Ĝȱm�z��~<��9h�xN4�����!--�J�Ww��Z���p�D3ڵ)^e+ �6z�J	>�&� _�'�� �Ƃ�t�=�e���!��Њ�c�mt����l;?����r��eMv�+3�~r��-�_d�����_���
\Q^-5t�b�����)��?���rW����@�i��"Y(ܦ�t���5�}�-↭D��Q�w�	Y�W�I�zCL{�_���'����n<���[� ��1G,��&1��:/&U(�(91�&�"��ٮB���{�h9'$AT7F�|ݫR\�<&� �.-�k��;*��ҸV��	 �
*$AGtN!/գ�)敄�]��&1p���c�F��+�����<����������-_�%B8�3�r���\��"3lO�Π�.��'�3��ë,��3h�_���u0h����ǩ�잙�5�dS̜�5B.d׌�>��)�!�
αւ�[�~��@{�B#Ӓ/s�9I���q;�R���rN�(5���L�ei�1�9h�#�0;��v$��~3_Q #9����� ����h�wWV��;b3��RqGt89&�F��I�+��>��TEQ�.u^�E��f�"��v�� ��f&���r&�#��יs����qW�Y��a�K&��l0�C�y�T�����6S����~��=쌎��1�����^��kuA�ƃ���Y�����3��/���'���Y���,u�(58n���=��K���ơ	~ ��P_S�)���ޮH~9�Ae$�]r�LN���x�ͪ���J���S)��m�aH����3_5CK�Q4��N�z�{����vZ_�PҜU����X�0=`
����bL"fd���#��a�a�P�%��#���O��O{�2e��S&���� ?Q���x��v�A>��aB�2����J!+�*�����Q��({�
�xZt�"�Z����Y���(r'�nZ��%.6��(6Ѡ�]^y�����k?u�A��0�+<�MY��9�`m�)'$�t��d�emL�A0��o�_\0��wS��c�J�V��<�Z@���=�C@;���+H����Ls���5�s�Ԭ�xR�m��G�c=�2���V�B38��*cU��fO�`�U�xD��LK?�~�"-��>Bkr{bL�g�-��w䅭���b<�;όc��W��mÃ� �I�z��c��(���lM������ٛqSY�>�;�4���r��V'�j�$���`W���ʀ�؁RsЕ��>} ��^��nX(��]r[%Z���TkT�F� Z�B��ƥA��`��:�qHFD}�m����I���S�9v���Zq��>#��9xi`���0ߤ�->�Wf F�1J�w�W�]8O�P�̗5��D@|���b��2-!�bM<�|ZTߗC��'ϲ|斻�5�&�l7W��q���,8 ��u>:=�����j�(����U�#��SƼ�{ΫT�y���$u�Gͪ�Z��>�A�l��Ea�OH�yq���ƿ�4/���v��9����غ^�={G�����{<7�
-����c���r�M��9|l)<����fn�l{P&�B}����-N$�KƂ�3*�ɥ���@d0���ǋ���89�-������H˃�W ��)��&��Bh9}�<Ѵ����f�qaB.K�i��P����FL���~Q�}`�ݻ���p8W?^%�,[f��Qg�}�J�nb�sɚ��1|��%g�'�P�-��H�f��cS�eܜw/�,zN#v���u��3vi���q�G��PyQJ2�J}B3T��*lLBho��+�S;H2Bm�t�b�nm�nR�Z"{�b��0�7�<�~c�&�	�i���\r(��2���ܪx᯼����x-ڡ@p�t_�4����Z����Ȳ4�Y���ҡ�kt�ɷbRU:w��x�kQ���n�P�¡�3P��3�8�l�����fW��]Us������5�.@<���w3gl(�*�Vu��qGc��(#�Ȗx�aγػ��݅D�)� U�e��$/��`G�3~����F��P�9��h#L�\��з�3���E��sz�Pԣ�Z�������:��r�9��₱��k-Z��9ͮ��fE��_+?�M�����)�PX���p�Z��QH����E]�?�|�es��s����vx�[���'�a��	�\6�w���㛹b���=��n�Z�w��L��)���a@n��%��Ro����>�݆!��g��mU�Z��y�2/N��ѹ�ma�d���J>ޝ��*��9���a�cg��1��p����B�>Qf���~`a��̣��A��W��[`���d�H �О.��iIN)4��L��'sͭ���E[���P�9c�v�i�
\�ӓ���	����O ��Y_J�B:z�:)ٞ�-/j�A�p���v	��'�Qe���wFy#Ǫ^s#M$���B�B��GC�̬}����?�,F۔�z�����#O�+�M�6:Ҙ������9n����C=
�(��M�4�X��.���?�pE��>
6K)�͚��=�h�Ly��Q�L�cSlz�ZM,�jCV�v���n]"���;���v��8�h�)!��?��V�?<�����T8��%QK���AG�KU�3�	�EBWU�=�a�ڷ 	N/9=Oh�g��|�P����2�8���4��~��f�j�g�hs�ztr�Q����r���Vs:&&�-��"�IE�?�?^2L�0X�ېV�8h/F�-0�}	����D�$8����+ �Tx��8xK�Y<��Q!B�\���|2�aUU�����kf!�I�x+/�o������� ��P��]Z�썡��O�����U�l�Dהs���Bk�|:gD}8@"�<�az��
�g�(��v�2|��s
�3�opPi_�w��ܯ����N1̔�b��>:�=��D]��ڃ���S܅_����B�ʺ5FvM��&J�m,z���B��_zJ����_����!��k_�)�ݫ</%�����Ns2�ՖI�q��\K��2S'65mg4+Z�VE�W�p�.ŒL�H� j}>dZ˭Dd���Z?߰���]��h�H!lm9����l��<�JSQ��@r��B̴޶�Y�[��<���4:Z2J��\���F�$}����G�;����H�s.E�Z�#"��w*���9UU��(c�\���z�TU�����j��Ϳ�d*s���y�U�5�Q��,o6�c�i����w~���i_�f��� ƃ?Dg��f����udh��^G��ʷ�j�����远�'�H��a�S�k�Ɖ��U�dL��N�sWt����?��(���Ĳ&������ L$�iv1d ��F�]v ���7��\�P�-�^��M?l2jD`������:��"ΐ
m��:O]�.C��-�'EXLQF�E�I��v@Xo�мxe�_@_QQ�,"%�?����o�W���%�	�����E(���I}0�>�Rcx������&dR4WѮ*޵�q���<����X�ildm&⠤����P_���D����m��7Ze����E�Y�,M��	V@�z� ���TC�1���ME�"�o^7tM#H9��������`�)?�N���S�|�$;�����D�]��㋊з�>{���g!ߊb����!?4��N�̮2��<��7,��ܿҾ<J�u��6+�Ox�,��1���\��v�}�ƽ~�?¶�Y��9
��n�_�u6�I�5�H�}�eF��&Y\a���aNgf�ϋ���Yz�)��߈���X�Tڸ	y�\��n�t�����`f����_X���&xF~�yO
��Ӑ�F����Ȯ�������b���P����E�yu����N���pC����僊1P��ql�!�ױz�ա"���$���jhz�=�����^��E���M��t&z;���y}�ϯ�#�(�����j^#r_>��[/�"��u�)L�%>��u4|�!:o�a�8��X����gL0�v���^�5,����E�E4QVǁ��hm�+ '-N9<�x���oH� ���u��u�j:�)�����>�9�/��Ϣ� 8�v��"q�[��]y�y�$(n �'�C�����]&��W�M-��z��Q�9���I=��_���6Kc��'�������=�33���1?9b��+��V���b��n�D����C���ڨ�{��Hr,�R��4�/��.��;�W��f�܋h���䙗�`h�˓�y	�b�\-E'�{l���Csa���\AI�����̠q�my�A�I���L���C��s�I���*��zP�;4�Dg�񏕨#-�h�L��)�*��+_�p��Y�D�7A�_'�rAT+P�g0��]�7AQr�c�=�{��r@M�w/�j
������ZB<��w+�֞�d��-X��4�ɼ�PX`�~Q�-Vk{�2��#̩�\���
�w!-�B����:9��̇���b��f`��y�
������u3��uБ!�W�*p�(�mP�QF��.Hs�yx�H�ȟ�xv�u'r�ٓT�'|F>��.H� �jV۝i *Z�&�B�����歪i�G�@э����Ur���'�i`;��B�E�L ���q��;;XkFF6�ȗ��{��v��៺j�[}��㰐��r4�����R������$��j��bSO�,U8��27�N��
'��Q?�)�*_�:Υ��Q���<[{齝�U�NV������ɺ ��O����*	I������X)n�.U����aq*�6���M� t(�j�_�ΉmAh��^�O�*kx��Yol(Պn�l�ĝO=],]�C����=�R !��(�|�I�Vl���7��0|a���%�Oa����s��s��&n�2�,z�ҏ��U؇M�ґf
��
[г�;��O�Ӷu�c���"�����1�n̜�V��r[���c9�j��Z)R�q�ΖLO"d{�:����T�:��~V
 K�['ɖ�����?Z��gv��ry$wEo��g:7���^V�Yo` ��t)o����5f�;�HU��[���J��#x�z�o\��c�����n,��m?�DyY�A����<^A<_A���)�~|�����1��%�6�\՛0sB}�����6t`���m�ʓ�4�x�,�*h?��l"|����Z�u'ꕽ�fϬʄ��=#��sa*w;�n�	�:�o9���C ߝ͚��$�|�[g`�f����=���(���^�M���e��<����W�>Lg藥K�l����_ҷRW(d�aC2�7�� �22"1��$Og蒞2Ō���/*/i0��Q�>�5�<*��(���p���d6
�n�I�M�'��n[4/��%���"�}����oj�`�@Q��2�G�:$�"��o�D��j�}�Q>��_ ��VB�-�Q��=$��_ٺ�t�hV�5LE�KA�sx�H�/Nw��
�읙\$�Uf3���\�\.���&���m�)��^�,��ȱ���n���Df�@C�x^+���f{g�E��)�����I��a�hJ�5�y���Q!G���%u �~Uj��hY=�i4�#c���窃���ڼ�k�Q��=U�֐5ϰ�q�)�<����Jݡ��+Snk���� �h�}ڟX'1�QV!s�\{NT�5�Ee?�ɘ���kBf~"ԓ٫�~���?A���N��=�8���1�x��^ޭ�y��q�}���� 9�v�?��"3��?g��vj�0�ax\���Q�iW�C8�����ݟ�z! ׏�qxx�+Ds����D{n
�?��a��.�ŨB�#U���7:)xq1ş6�EE]p�y�΄���i�oеviu�^pݯٍ>��dĴf���id {�1@�����:�}��q2��s���u�$�Iੋ�����̅��>��f��.g+��V	iOU�u(�\+(h)i^����3�>�;Q�ާ�2r�j�Vj4�Y~^S�v��q��L����N����+�������ô�_��)H��M��ݒʢ��wy��EMV���1@0%�m�с�x�V�i3���\��sYkQ�����h�)�c��6�϶�����t�S#�=M3�H$�QuΡ��i�$'U:Q��W�+O����S�-��_�/�K������J�#�k��ڽL�Ѵv8?��)��@��ɶ0�!�;n�Z�= �awϣQ}��U]4@�,&/^=1�zr�֚]�v����d�WM?_���!َ?�����ږ�@��[&���ە=����4%`�m�H�?�pA �<у`��W
Zj<zj\��p[�S΃k��f�����]���R�g�q�s���P�p�JW�3sQ!��[}igE�	���i12��Ap���!��s����Ď�����TwGa���YC���;��8��*�
Qn,�Oc����5�+2�b7�LK{X���3>w���B����K1�����p�{��D��6>9��E�؃��-�'�8��E�В��w�`@�\|Ɍ��J�����1����
�5���f�T��SVW��7�/NKk( +��A�5�^�Uf�X�B�rr;b�L ے��8rP�UϢ�����jA}jɾ�(�t��6�������� �P���4�$nk���7�I0���^��N�C�n8���'�k���$�;>0<Fz��ɩ��Q��ʑ_�[r��+���{����XU�A?q��>S�2 N� ���e�����.�?<�Ew��,!��[l�Y'<�
qS�O�*�㧇%3u����" O�vg��@��\h���oe����9�{-[�l��ʻ��F�
�y`;ﲿ��	�-X���y�� �N����F�Ì��Do�Gb���hk�U}P��v�l벬����P�z��gG0��y3t�*�&���L�W��o$�kK�p!�.�<=RI�V�%�|��xJ�
���>F�SR/�:2��40�Z��7Ե������Md�&Ѫ�����#)���F}D3���s����s�+'�H[o�=�fv����6^� ��~;�z�l���"ԫ�I;V�@(����x>ݣ�Ml��%�� ��eh4���%���^  
W)A��(O&�$|8�� ����Ρ�M&��fڠD��A��go;�2�$�\�"ԇa�j�9ُA׫�t/�G����}p�3j+�R\��da�L' ����q�c=I(,�?ؐ)ݮ��YѮ�%.@L�}�Z�;�
0nH#�m-zly5�p���;N�U�j�%���3�OV�8&�`��K�3�8�����2|fZ����ϼD�+�ƕ@?TT�H�&�fsBRI�ŀ�CW�H7	�To'���I�/=H{���\�[��I�m0r�E�;N��.����	���s���y��Nْ����a��Ɓ��]����r�<D1h�~&�{���͙(MlglI�&'siߒC\���c�v{��X��K�o{� -ꑵ�y"<J�רZ�
�Q��B?���G삶�����i�T�Ŏ��h���[�����	1ثv�@�aR��p����[YϜoq�3����.@7�a���z|c���`��kP�۩�q����~+I��|D�,K��	���� X���3��Q��^�j|��ۨ<�@u��7�e��;\��-83P�Z���՜��F@�k�����wO�͂]&�Nk�T��u�̿��N�ԷF���a�鳋����J{�}m�lZS���Ǧh��ç�qȽ�p�{0���H��˴#kM,C0G4�U�A3U�a�ZȔ��;��l�q�(�y���yz���8�]13UP��U׺�dj{��(y�p�DdFXq�?~�,���v�m>6afKs����gNR7t�G^��_O�u����Y��ʐ���vh��˛4w�쌶��ÎiD�^�Q^�u�lU��ܢA��R�bZ�\@���˨��!�)��w�p���1zs@ӧRZ�)���R5��z"��Ou��+8Gb����_�e��QH�qm���fVg03.؅��V3]����ܒ�J��C�x]Vs����aW5�w���`��tl����z�&J�M>M���DfƔ�C�Ȱ?������U26rb��H�b*{�v��a4w��W��Y"��Ц��Wo�9*��5�Q^$aO�ϛ{�h��<���s��#�Ȝ�W8�6v0��3�Q��^��(����5*�3vG���]��� ��'T䒲�%�߶�M7�v/��C������%�|�%��(�:F�O�Lﳫ!��W�b�K�o�\�{��V�j�Dc;�Bw������s@�A����ڨ��IФ�ɫ�H�i���=��[r*[��_&���a:w����#e�A}�q�4JΆ�%,��:��	`ܼ��&�YN�)���(�(դ8z׷�֟dlQ1(�r��7�]�o?���hQ�Z�� 5��2CV�W�ڽ®�#�����0�@|CBZ��f�G܍���pf��{ݯ��54DQ�e�xO�����ה7�X���j�|��V�D�rd׸���|�V� 0\�����Ѵ�Y9/q�E�����u�OoY�D�
1�<1�r�sЪ��(*j�c�%�~M��엮�C���	'[�<�$�n�"�Y��� ��Z��iُ�M��]~+��^����Y��a3�����LQ������o)]0F����ȗ�5�aJ0w�u ����D�om�-b��w�s�����!��2�f�B�W��O�"͏c݆��x����ēcE���XQN}_X�Ύy\��F���9�vp��*P��.��Y���{�Γ�ي����.Wm����ln��*5��4KNR߼<4뵫�>i��7�����Y��A}qG��t�ĝa��'�bk�#���C���r�Z��IIQ���<u(U�8��AA9~N�li!��IJ�y��DL���^�f�Uy�ʻ'�(gv��܁x�nNa/�`W+�J~i9��i�D]�ev0`��a�<,Mz������=J4�1��,"�p>�4Q��3(ּ;\LD��9�k�"Q��SZ���L	y�����ũ�������oSw$^���zC�+�3W��?Y�2�;�B���Ĥ�0����@��`A� �Ll�m���\�f�`X�jz'�����>����n&��Ԃ,����|㸗�E�F��Uk��-�:f6���ݾ�}��j�0[����\��Ke���
�U�����B&��NiGp�X����k�TM��fwîTC�j��؋PUo@`��b^�pJ�99{2!Jp����ʛa_��^�=�p�0µ�[�t'4��h�H�Ѕ Gpe�8�%����wM���de���*](Uqc�C����DY0_� Z=�	2��ZГ?�?g�4��xnI�����ISʉ@qP�����E������|m|2>��;���������6��2μ����$���I�g��������weU	��HEX/\�Kx[38��LsXP|rA�h���*��<��j¾\��;�9�5;3ǉ�OIp�����)�J|���m�ݣ�@���	ԊV��Ɨf��K��J����@���v8QF�ҡT�2�@R�Ap�W����j9Al�(gJ�!oPN���<j�gO���u!8���A��{�B&�a,��JQ����D�E�p��Er����}���)p�q8�&���.���扺 T>#�t+4҅��mދ��vߑ������ūwK��n�V�c��#�,
3�QzB�+$G�O��� Ů}"��:P^-"I�#sa	����˗y�W�:�=�4�g2��y�b�5�am2p�F�O��&��Z��Apc��0M]?Q�a������?kn�F��9�P�;�\^;\��p�;e9Q ���H��nѷ'�9�����;�g|� �	���Wb59��Cx�D%|�eH�YI�r�|іS���D_G/�	xr���?$�%<"mU���+�G�y`ʝ��Э�3cE�ʎ|
}�a\��O�9i�Jk�����Ң�y���[|�=�!�`����E�_L�[��%{�u�0e�h�wjlF�_�=���g��z�d��
�$���{��>C��x�,.)�����Z"���t�F�b�
��f� �_�3
I��N�{��#FѢa�i���[���:�|�ȑw��(or:8Z�[5<$�Z���H�U��l�ЗE�|��%(�S�yxQ������Cn�&��93a
��{��g;S�Z�'1�fnL�|���汦��]��nŊY��&iu�i��SN���
I�E��s��j���%����x�mG�������g8_�5g=�/M	R&��g+��*9����@}�]ϸ����8rMm|JM��)�mhi6��"ܐ�D��V��Z�8�󅾑��S�+`?Iz�#/��Z�a��-��m1(�9�l<��fD���IZc�{���4{���uF���b#��W�Zf��O�?�I�"��Y���S������ʐ�����O�����
�Q8�OEr謹�������P�5�f�}�˞�w�W/�kZz�Hҗ�R7�4,�wDÙ;V�ʖ"
6�G��0}n�2�;�?�ׅ�����,��WVDš4�s�~�PV�[��sԊ�����j�F�@PV�9;��9t�Z^���)1��[�m@(���Qk��"=�Ҿ�e�9	h��P�Q����l�%M��a�`�^D�3�]������e��wfp��ݰp��<�6�ja��Ea�>=������FÎ��`� =�m de ��  r	�[�s@��<���m&C�$\o�3�<�p��tI�}x���0��,>+.���`�(�Xx�a�,�R���T�u�3����OԤEϱ�)�m@!��u]p��k{�*ui&a@��K�2��g��qk��X[�S4�9�n�p�->�W[�0�&��!�����53���(w� CҷM9�+�rW���L{�Yq���te缆��0!T] ��l�w^��׮rWi7� BI����i�?֡v�9���r��︦_�da���.���V=���0S�P����q'̮�[�b����NQ����G
���QJQ���7gs�4K?�1=W��g����K�
h|8K��N#.W�Z�ڝ͖�sq�^�0�Q�ʀ�� ����޻��͛N���2�ZN�'c�L�����׋p�N𑖇YȊ���&\��TjE3.��{������=�|��2H��X��(X���L�u�J�@�KJ�a^�18(ğ�v��1$���C�VX�����KE�IH�)(�rE���Q�ᴱ���j�B�-V�՜��6A�([� ��(�z�?؍�a͂z;ͿQ���ٱ������=D�yRX��s���\�����g}���b@���\1���D}�%,}��ކ���&�MOz\5�	ʝ0cZ�5�ߔ�����T�~���,�^��KK$�GI�k>�m��#rҳv�]��Uf���,<	��6���&���j��� ����Le�IR�/a�n������|�0��:��)���3���3.��Qgu�A����YM�#|/s
P���fJ��~�#�S*��K=\ng�*\HԺS�T2\�����=����_��Ø�V\B;#�<�(���2�*�ұ9>�z�-�
�����[Ȑa��<��V����7x=��Z��6_�/����E�ϥ)�9Y�s�p�ֈ��{�$��dd��Es1D�q�㢛����Y"�m��
����FqŀHo��5w�9MY�~'�f��v��/5����p܊!m"A��l)�"�:�Rc��ߜ	9����)i���а�����+3L�Yi`�%p=��	0�⭐�]^�'�Br�aV����u{g����#��_e����nw-�ot�c���Ŕ-�7�(@t��o�_�x`,#u<������{>���˝��L��j��ƌo�Z)d���ո9�
�x+���:&���yl1c9���NU���>Y_�y��˰ ���'�eD���<��؅[68��Fx7��jr>*ϛ��E֖���H�$z�����ΟvÇ�@����>��d�� �)��ǋ.<.��O�����LD�p.v���B	.���SV��O�P-o������Gu+ȕ��z!��XWk˼�O{��z���$r�˻+1��U��QZBƖDM7�{�2;�5+VQ��5�kデ������ۧ�z���7nJ��l���g��� �UݻCo)�i"�
��|�2T
�o��=w�<Ä!#�uK���^��lC&Oܛ{�����_/|��;�`��λ�3��C��Z�}}YpH�Ezߪ�mB{�X�ү�L�3�W�[_5AmR�b#}�&�À�乶�#bC�<��筄
�q+"q9=����M���+2��%ghc$�}A�rG%�M��<Rܾ�5��o X��˲z}%��.<��ޓ��P[��G٣���k�<|X2i$:�~��4��+�@U��K,!�����]�;���,wu�6C�xEO��.�k�B.ɰ��=q������2d��_����r�Q�K?rj+�_��i~!H�c��M�#4q\�;���K�ox��u��o=����ΗN~6��;$F��O�r���9F��ѥ��cц>�.�O�1�m�!e�~^я�,$�M�5�.\��v}��>��@�zN���0R�����G��饮�mK��&L4%f�������C�]\9�7@`�d�Mc�M������ä[����&v�٨Z(���ij�<�lr"�E�t_ $F�noc63���S����w�6c�o��*' #c�K�	,r��xՔ\���2�U�ޫ���V�'^G��T���u𩪸�:ԏcN�a���Ւ����G��\b_2�[����ٹ"Z���ja� Y��	Cz��ǀ9'w�.@���
M]��9K(�lƵ�Å~��/D&���/�#� P��Б)���vOJѳ/�Ai)��M�dXu&��+�����uDI��Y��p�6i����tn0�st l�],�-�>O<��W�� ��E�0�Ɇ�E��BQ����Զt�&��^4��,A�j�W��� Q��Aȓ����_T�9��U������3h��֕<�&�\���cF#���Bl��i�
���sm-��vt3����������K8�j�aP�k��z1V�3ˎ�~#��I?�Cg<?lM
��ؠ%j0�Y�˯�+�IE�.�s���?<n1Z]�0�F��o�8ђ�)����&�t=x��oP
�w������V`���!��1c=ިU\��o�Cs��G#J�J�]A>%h����E���^�h�4!nu"`��m�6+�8��m�lV)����_֥6�!hƢ'�1��!t.$�D�h�nV!{��wq;�E�P�(O�/��ZiD�֣x�6�O��*�hzX;��bK ���J����w������#e�d��O��9�K ���ǃ�?���T���0����O�p�|u�U�Vq�� l�!�)Q�D��q�K'���f��vQ}��̵�:]!W�-�s��o|��r��&��'<ćYjg������7�"������rs��!���y�%�~O���hJ��	y(d	�K����2{z��[$I{�=�N��e|�5���>��P�1On�W�n��_D�
 �d5�6R��tom,</u���S�祒���)�[��Ǔ��k�;��B��)/��b�1?"8�=����O{�(_P�\��?�W�����	;昱L��9R8��Y6c��?8 巐Q�z�����A`e���ˡ9�����~��^Uⶻ+��B��ԡO�Z��V�p�xwl��*�U�s������"�,O���W���L�g���S)zLgF�{jS���ԯ��l+���ۋ�s;i1�`�҅i���NɅ�Fϔ�ړ�)��z�
4^yb`rP	M1>�p?i�Us�`�W[�������v	��e�����v�3�C>F(/�k{�+��i�|l�&c���#Y I#X�G�﯂>P�>*������͆g�$u�N�g�yV��(�(Dt�;�,W	|�A�Y����T(�N���˾�xK��~�=��f��;W�H�ia����Τ�?w>h���w�χ��
��K���-����#�3�c��^���{�}S���_|��wk ,g�klf4��YX��!�fֳ���"�	'�7�/mS�ǥ�G���既Y��1��'�A�al0 q��7��ñ'���.��@�t������p��|*S'�IS��g�%f�l���:��m�,�X���XM�V?��5�G
�	�6fB����ȥ!��Dy��N��[Y��ЮB�r�rХ��k��1�{�3�ֽ����(P�p!*�79>!1�%_��i�i�!�[y�t����r���l0ut 
4�x�K�2I���&Ϯ<�1O��+ӧ�goT=.EPU ���l��5�Wh>�ߓ���q�{��^��ݥ���X��lq���wt>H� kΠę����?b̪AGܻv{����=�݌o������w���6m1>�A������xXI��g6V����a�e��<�ڭ-�n�6eF�^��������d|\�4ڭ����h��Hl�Y��V$no�1�Q"gVB�����@V!�Ki������$���_�a��L 5�F�(1��4���_���>��޳}:�c[`-��ZNL��g���{��k��X���^|uN}�
�lo0:���<f���hx��f�mM��qL���ǁ���;�5����4����'5R�d�
f�UH٪q5\��;Y�O�qEJpx8k�������G=q7�)��V�\:�a��=5}<`rt�p�e��bkF��EO��\�'�8�،���LWE9�L�f��8ƪ��bڙw['[`���(��^VlZC|sV�4�J���� 4X��"6kx;|#Ē|Y�u4���֭멏l�2�cvn�
��7�
f����&ճ�Z�N��]p������I%�5>8M��i���q�U��%!�\�考��k�]6�;c���)��e����ƽ[�W< ����x��0ir;V������z��4@ō��h�IW����od�P7�����J}���o�Ơ;�而�M�g`&���8��w�V5`%����<���w�4��ΏV�0�ùː4��0l �2/Ϊ�LGF卓�J𡙣�!���>2�6Վ����y6�P��E���P ��Cp?'�d;��Ŋ���F �ʰ_ �i膑��뮐R�}`j� �n�q?�e.J�
�oa��P�f�w����]�j9_\ .�D1�Zs9�S�k�=��=�Nh����1@�_�^����y9��Ȯk	��%�e��{C�^�(P{�E�ս=�?K����1��
8� a�#��O�ʶ?��{3�_�o� ���
G�z��z�"v��U�čE��ا
`�iR��.�E��{��x�c�f|A�"�7�z���(����\�\�Y��T�+�\Zi���L��u֒�H �"���.�>h�����wpC�
y�\q���!_�ޥ�b�=����l���u���(پ�X\�r:�"��p�]L��ӺA�Ԅl�-r�U����f�o���fa�Ϥ�Үe�y�y�T+a��~��=�+�U"��̑��k���*��3�5�)3�i(��2�c����Ȣ���r�����ܹ�����[����ɖ�\{`'~�lr9��g��	�d ]U�S�(��Ĕ$V5Z��迄�8bȻ��t-�c��;$k��X��Ǐ��w}[S���3L0@v<Ke"���	�Y���ĘE�I�`7��{�Oȼ��]�#�b���@nR��Q�����U�bv�#S<�w¿��aKD|Z格H�^-3�',� [����cA�V���|-v6�4it1��ϋ�V���t	Şh2}̻���R��Zh�}���@��ŧ?�qO��-PX�,�����W[Ji������6t�0	�K�y�M�a	�ԉE�h2��Y@V	�λ���@8x��@���K0�o}�ކs��,�mP�����<5�EQVi�l��M��������6�����LN^�������UE�4���c�=Y�!���Ce�N���ɭ�Pi���w�8q��e�ǖ��)��O�"D�H�0K������f[����vh�̌��^�����1يɳ=?`ۀ���I=i�������z�&��]ou�'�օ�hteЯ6pt$��� �1�J�dT}����������TrGҎB��%���diz'�����=y�2��T�Õo�Ȇ���d�ns6�Wb�S��p��cN�W��~�~��5�-�_$uN$�ѹ�5�ݮg��d?��<*�N�&��Q�#2Z�68܃�m�J��[)̒�cQ#$�!��u$,�$�������E�pR��6�~�Ҳ3 w�k�H(9j-؁�L��V���wjq����'\R��`��>�*Х~h�;[?���\`M�6����T�U�|��>���#z1F3K1��zeq�,KT'~+����� I�����Bf|�
��WE/H�l�w��:0TWJ��"(�(��A1��,�O�U��TQ�A�E�;5��b�f<d#���B��F�댴��e.��^ީ�B� u�+_O$TkX��)g���0RҔ�~p`DͲ���e3+t�a�P?QRK�G��&�Oّ�s~̉ͻ�W������}R�^e6�C���h��a^���I �v^櫤�/��aW�f��� �_I%VH�&�=�����"^�+ӋV̦,@x���ҷ��gT���0��D�X��7�PI#���z�ɿ��X}gd�����'�8ܟ�=�:�]LH�O��$~� *1�"bn{t#U�V�PL�Q%���<�߿6*q{}�
x������H��r?t�y��N'����i���^�'G�2K����]\�z�(�-R�}�5�9�H����M`�p*�e�Η�+�)c��?��p�W�Q��ܦ�s�K���+
�%��8�%�X��daHFҫ^O9^��$���'e\�c�YJ"Ijߣ5!�7Fk]�e�����Z���x��|����O�z!l��e�9�"zVݰy&B_�s���u; HnҺ��M2��c�n=o9�f���ǩ������a�s���̘L��kpY֑�PK&�u������5t���]T���K��YC�{��we_|B�W��<��0��^�����:b��;�f6������HBW�i�S���N4�G�S�=Хx��ا��Ϲ�q<	��ov0��pD���˘<@E�&JDJ~�k+�\���K��CI	��3��-���+?K�n�ʎ�l��6��f%!�Ax�"��u;�?pai_��U__��sG���e[f��u;��y�:r��;�(c
t8�顒"%�~�cOj�z ����X�F�*��﹣8��%�8~�G���t���?坌��3�1DZWg$�;�:�w�i.������¿8��B� ��e@����x�!d�h�"��:>nRs�92�!�;�����A���I�g��&� #��Z�/?����趮v�{��ڶA��>'��.`is������N>kj�ٺ�"R����.=��Ϟ"I�?PگR��QL/��2V���8'�7��)�%Vz޾�VЍ,$��?,�B�8�3�`��Խ	�� ��<Z�̚�ei����y����4�1�EcE�_�t��X�Z����f�: ������~���o+BPѿ�����$K��jb��^�<T��$?����'����9<�U������O�wG.|¦��غ��'�1�׀���c줮������2y��Rz���ޤ� q'i���<J痭tQ��E�\yz����LQu���\������o�mO�g�AU��l�#k�)�`���e
9�3مfG�^hЗo��p�Br�6��^*���t���pX�Dķ��H�W��V�b��HH0���0��?� ����|j1~�����q�*��V�{#��>�0�) �b)�}�>ig�p����IX�\E�MV��wڞ���*X�R�<v*3�ło?;�SAe�q�|��l����GQ/3�vb�9�ح`M������x>�����I5����J��u���	ע�z�PF�ST�0+m�-��di�QC[���0���kUp�j	���Ĳ�����[G�����G����`5\�͞UV�F)���CDl����+#�}�R��B�ؿY&8?6A���QV�_A�oP�oĞ�)vY2�-#�3�~�S���l��b"���`	WW�u\"�p�O��^v��ɮ��cC�ۆ��d���<�&1"r�$�ȯa�0�sJ�ְK���7�	��[`��M����Y����`��G��=�o�h(��EA֙ݶ��>�},�
[%+�-�D `g6�m\CQy�m+�]3�=(�o�3�)���S4�$ZŶaJ�#���KQ�N죣��+Ѩ�p!���.%&!���3<��=����KAy���x�޶�(��2V��j�ϝ�-\\���QSe�����kd)��!
28�5 �_&߿u=�8�Z���\�h ��}��PoH}��������*�g�����!+K���"Djh��sod��d�ּ��gm�W1�}";)���s7�ST'��e�2��>�Z��s��U�>��!#��`[�NJ��f8�J��&#N��$�B&�l�P���t�|�"�)3ю�2�(�������w�f	��by���ߋ���rp(��f�S����̻x��Q�'�o��,["ǫ0-`;���E��E��	E7�1��_�mӹ���!_����R��15W-��J�J���%���-����@$_��Ws������S
�_>�����0v�=٥�q,��H�X's/��x.WGs�1c���S/e�e���U�9�[�|�ML�uA;�q��E,�{�T~�16FGmG&�{7m�5�|w�1��Ŷ7R ��_���:�����b��]�;��y�Ë�ߍxל����qf ��D0By��I�ܐ.��>�<��fR5�n�ݱ#j6�Y�z�ˮo��B��>�fhEiC~� �n &YX�D��{�h0pQ<a���<C��U�6�j���'���z3y	ؘ��AV�M[iU�(��zH�킪�T�L!m5��6�����J�uVCDqDs5_�`�z��єKn/wuF��g�Z���ݎ��4���ѓ���b�}��𸝇��R�?7w�:�c������>S���u��k��2��������9�,���l7	�#� ��!�����wj�]Z�v۵6o�/i���K}��S)G,<u�5m�]˩��FJ��	-f�Y��~��>�Y�7"h��)���]��,\hS4z����@��IRq�*��Ru���>�%���4�g2H��l��z��
�1�C������*�����;�&,����F
 �5=�����ޗ���q���$�H~%�=[,�Ihp�S�/+I_@AS�>�|������2�U,�!�-�Rk&\���3�Ҡ��!Rl.�S4����*���5jj�[��;'��Ī�{�704`��P��6�Q7w�
`��̨6�����(W�M��7�qP��VX�T	�P�~��v�j��q7��ʵ�ye�;�'*t���"�s2s�m���L,R���<�j��ʔdߜ��0���E�������f�&�t��o��d�C�]R@ϱi��\/_��_ �xc�:�(�m�P#�y<	R=L ��v:��'_"�
��f��QE�ݚiw*J�A���K�S]e�o��9}��}k΁<Y-�H\lM��X+L���>n�����0����w�y��[�UzS]����i\-`�P��i�+_�֍�a�p�������.$3�3ۯ�����b�i���-V	_���|�\�h�b����l��+�'ԇf�@�������`w��<׬�O�Z�� �>�P���T�	�
N�O�m�Z�]4���'�[HZ�d�9\HY���^@2v8�n�27O�W��+�찮k�#C�On�e�&�A��}�r���Z��L'_������}h���dY�o�ퟡثp�-�LBV�q�]Zk��^�>�Vg�V�@ aE�o��$���(V��S�3 �đmt�P��[wG����m���uxY"ߦ�
�q���K�;V��e����f�j0� !&|O���߅C��L�|R�q�˪&�����R�N}ג�#�n�֫�9����*��6�zQE��G@&��FN�B�� ����q;�[v@# u%WO�������o��j����]�����%���i�+�*fȹ�G�9}M\�; �FU��cp,H����_�~i|/�l����0u���z��B�>"���Ǡ�D��Rb��#�^k�����i�jV��eI���}cB�c��]/�9%+�p����F����꣔��f6�ڵT�F�'ͥ(�̼�@��� (��?A@���v\�)W��C9�ąf݆l����6�%mᰟ�����8ݔ%�5��/�c��G�e���>�A������vj�9R�kT#w����P����	7�q��͌@"ș�G��&^�UI�|	�����K(�QOxY�Z*n��a��P1Ar[l �dh�!�+<S(3;+�9�E�&�ѵ?��z���S�����7g*[¹_��S��ޖ�3f�wޮ�#���hP���b>4��|�˄@f���>�G$��_3I�����;&8?�"!�������0�;d��_AD��n(�҃�;Y�P䃁�m�gW6a��9=�jA�!7[b�X��W3�,Z��N��@����B���Fܪ��C����H�/�o�$ �d�;3��f��4O'I�`[�i.�r�U~6!�p��5�oQ��GBQ��c ��\ 0P����N��_1���W��.�V�ݻȿ	��X��V2�{U;�X�`Y�d�B�K5�.�Q!^��L��QP��ѡ��P�V	��՘���Z�����)�wTx�;۽�sЍ�j����5��R#)#�Y(�T�Pn�����ŖG7�qi*wfnU���UW�R�wKQRl,A	F�W^�_Cp��X�X88Q���1�0O�B�ɩ~7ژ親"�dQ�c���V��j�%�`Z'��s�ne;o��_��%��6k��o8����٣y��W"�+��J��_�X�1_�A�ӪT{q����Ċ�8p�ꭧ�!\�CI<�Űv��:���Z_x:40�Y��?�MZ�
����h�C�,�|.��!��?D��bq{ڐ�uBQ�k�ڞ]h�Y�<�؋���K��%��U��`���PYыUe�e0A����wI�/6����5��}�J�#�b4���跖Y�ª������:�d��5��P7���������(��A��|�G����(�QMWf #�`\$���5�q�l�L�b�z+�]Ip�+�~��gրXdք�#]L�cE�v:����Hk�hztC�'�U�Aw��]�8�_�M�������څp0�'Z(��3�7[�q(V���Z}��T�H������m]��Qh,ѧ�ʟ�YlF�G��U��ۄU7���(U7�`�ם�]Q���|��WnSSk�yӆÌf8�zU�oRq������n�bgm�φ���e�旡�����R9�fě��TF�K��(/�G����mzPhL��SM�n�e���k����ϲ��j�細*��)��ZN��_Lo��*	�[d5C�x��w�s��9"6"1�X����K�8J�HR^��T"{Z�c<���yg�m�b�＠ca�����S�$��T�~�8��g�V�z�\��Ĺ)BI����QGIsy��҃��ՏyBj��v
mk-Am��E�~ٲ��2f�z��Om_� o�m�ZH _�l�Ö�,���} �,�H
�5KEl�ks^?R�Z)L�E�T�n�36/���Ǒ��9��Eg��1_��S=	��m=���7��R���^�_.���k?������+�
Wj���{�������������PhNO#�s��8�i
�0�F��Z����h��xpݠ�y��Ϟ�!��� ����z��E�����K3�P�hZ˹50��!���fO=5Ժ����N��J�޷�e-<�U8^�c#��>��yr�������;D�@ץ��ɂq*۹� ({�/�,���v���?�hvh���L,?y�u�G�vv���H�1e�<-B�`�t�5+֮���N�����h���A����(��T��I\�]#���{��x�ŔC��#%�I�M��.���_ڣ�2k1�t�u��s���a�}d�2�������Qթ��g:��=�;fF)��*�yh��e3p��5妥����O��3�c��׹7�q?c���۷�����g*�+\7�U_ڎt�g������[���=Pd.��c�ho�<�ɹ^�yr���d}t�	E8�G|&�0=
�em���c�:�T����O" �����۲=��?�O}����'���G��`��)���C@����h�k��l�Rִ{!�li�H�)�Ȉ(�krh���3V_L�c�f�#S���I�b��Fys����fCsř�A��`�e�g�+>�:��χO1KX��Htd��IN��j��e����TM2*@)~����}��h��ɑ/�s�I3S��-�����_4�F�fS0 �D�^zG����.�R?�xHM����ϸ_�����+�6���=o�W�o��&jH8:sǆ<�8'��������8Tn�ٗ{��Zi�c(�21���۹@�Ol�/�����׹��6<��8p}�=nߕIB��d?�K������
�r\��4"�����&����x(T q:Ѻ~3�q]�1�<�c�E�lu�
Y�.t�B@���Au9�l�����`�BS���8��**�ɧ�a�QE^	);.��� Bf�sͥ3m�ƨ��k�����kf4��Av�fj$"(����}GĪ>=M�S�s�8 ���|8�����,�}�}��)�f�@���6�����$/�NA�M:�6���1�9��_W!ql�
{�r�6� CA���e�,�E-�~��J��c$k'�Pvx���Wk�r! 5��uY�(
f5y�/���+�PJ�g0�ҷP�9�׿�p��ޘ:Q`5�'Up��WD;b{Zt~|8]�3��V<����>�+V�H��+OYۆM� �4j�9=�)����G�?	5��V#�+"�d(�H��_��ȕ���?�"P������dzo}��\O3���I�k\�]p;�d���L"�n��+B�^�@�虛�@���[�-�|�P��u7�(g�[K����}��@����7^)v1D�y���B�d0P��b�a�"�.�}�0��~��{��Y�O4%{1�Q%����2-X�R�g�r��5��1o�]ƀ��n[I�3?�g5��3:�H��/:�}nzŜ��~Aw��&-�ur�;]ͫlMx��K&'�rDJ�a"�´�	v)�Ո�\��������rke�v[X��Tk��������7?�� х������X�Y�L�nSnMuP�m^`ӏpb���%lO�I��������yLD�ώ�W�-�+*@y������_������M^���O������}*Q���T���Bt�J�15�-D��[�\.��0�<�!�̓�šVj5�Hmi�}J8�ъ��ϢBz��dj�o��u�6$5;�j�.{��M:;�{����\�M�:�ux�|�Qn����S��7$&��3F�l������^�Y�w)y�X��]z�ר��K'�j朾���#��h���o��ڋy�e�ĝ�Z�/ґ� q[���%
��}C�:�g&|pڷ�D�W���o�����\ʳ����^�U��(]FY煕5"w^���}�g��܌rL��hIC��M�t�(��aG����.������}�j���us�^x���>��y��[�L^��|�W�h��Kl4�J�AƋ�Qe�,��+�N�;�7�֘�:�Hz��~�g|.a���8��vH�}��J��Q��ٰooyn��M��/w@�#��e%%	�,�:��W���}�K�4`�mB��A�f�C�4W�졺D"�B0&*���9Rd�T���?���=��w]�f}$���$��_P;�mt�i�%tN���W&("��w�_�����u���^�jF�mX���T���m5Qi[���oSL��L�0�.���&�����.�%�[�}7)�����-�_��@���Z�\�g����fY�J5c6�lS''XX����I*kq��>��Fn�IՔU2��+��ȅɣV���T��/�"u�d���~��t����/s!��a��4Igm���7� �{!��@�N�;�6�>Kz�h��޸�T2��.�fV�Pã�w3v��c�׾@��љF8�ח���u�2�u����v��GͪŉA���9���d�[�z�*"�FG1�MGY�!V:�%��I�կ)9���p���&�������0�i�
�;��`d�U3���_J����Ǉ�?�,����b�|� �89��/���)q)�w�;V?%����qT(t_ �&���K�n��!?��)����<�X�]���~�a�B�nlw�X"�*|ڢ=B�\�||�t<�_bJZ���b�F'��Yc��͑�������L���YFqY|�,�k5��{ Yb�ŀ�%��$&'|�z���rv�b:�L�,�L����r�����A�*șH���5���������Rg=Wb��Uy�|2u��	�R{����!�\��!�d�ٳ�`C�w���B�242п���Ɲ�Pc�T�� *��!���Gz�Z��w��7�������Ű�ݺAp���ɞ�]����?��uB}NQcf�R�"�����ᖻ�&0�_��Hs��Gy�Q��&HyJ2�	,�5�lHlk�'t�p�:��JAl���U�(R�>�V3CnC�܌!����L|Ǧ����o:
��ޣ�54&��h��W�6����WT9���c���G������h��3��,� �i@nÆ��fj_/+������?��JE�4�l�f����m�kS�qQ�L7�$$��KĢ�[���UL�N˚PbN�5 �����$�V��{/%�Fgﵪje���
��=����G+7L�F>�#0`�X���h�[Ż�|T�Y���JK�Muw����b��[���o��a�F�C����[��N�����~`��v���
5�	�d��qg2�V���X��B�����x���]����җ�}��Y	@G�>QlN�zb<XH�U����Er���XFL�hj���[����'$�[���Rt��z<O#{2h�B��	���[{�4\���\y��M{`d9��"s2��p�'O�c�����Y��������M���耽;�<���v�O�ٖ}W���@�g��h�|;8�7�Nڛ'�$\t];R�?�y�X���������7����,T���Ge�h���N�;�V�1**�T7�p��󎝠K�+�[�������?�Vg���ĕMx�[�����C� ���4�K�:�1����@o�C=��Zx�~���6�c�g=�ǟ��-Q���*�'�KA�GmU�M�	�2�K��EV`��d�S���Bz'����n�'[)��z�^�ɵݶ���$�jC�込tL�g�1����������:GP�G���ߊ����Yu_f6�l�|�|2���L���_u���)�i���]�6ޤ�(���K��Hl	v�d��)Y$gϲ8��+*h��aN[���Kk>BW��R2���(!X�{�5^���/t�*��TS6�-���>'{�[;e9��u6�j����)����2m�h�����V5 ��؜7�V����T+V+�6M��1�6Y�&w,%��d�2J���j K���Sm�L�2_����Z.`��-�9ڶL�R̗�/P?5�(�0����h�m�4���K2��#�~��J=~����0��iA��mD�y��D�%��$_$��A�`G~�Z�&J�[w&e���`��XT$����}<˛3�ʲ��7@$�#��pӱ�
8F9;w����7s�B(�l��~���vg�^F|'��w|8�F5�8���I6|�R%'� '�� �@Q�i��ֿ����v���:�>P		����Hׯ��x�@��0�p�R4vP�3Q����=@�	�.H ��c�V`����,�����P0 �8,;ޫG��M�ϧ�Ǉ���q�r�uka9��(�2R8��@�2� ��̐Uк��B؍�o�t���NթWts�����ã�e�X�'J�B�AO��	.�+}c,�-4I��ſ���u�l\��Ӎ��l#���)��$o��ڞ	��u2��bS��	$��6_:���~k��p�!�s]�k���A�2[m���V<�Ծ6����Ԕ�Z(���UW* �v���I �j�YP�����M�q]0 T����X�o"�E-�BIaw��ȧt	@gR�3y�);{o�y��ʛ�`�t`6;�>�5��`�9��wg�Z9!��˛�����=�T��z!w��c*�<05�^Z�y�B~e��I�J��J�ᗧ6G���gVN���VYP�l�ljY�����䛙R_�߭�V�)�+Y��c��J��I6��ɇ��"�����t�z�"3mʅ^>`v��hn�ls������/��{��6r�ߎ�ra��?�׸�K��G���Y4Y�G*�9�[�g����W���pܖ���Y�� ,�a�bJ0�}gu=T�$���1�O�W_\�����;&4�O�ea&�@�q��>:��A�}Ã��	`��J�[���i�#U�M0�
U>�
Vżr����9�1v�YsD;*��\p~�K���8t;�����(�b~"�*�@�wQ�6(����i8��RAIq1����|s��R��i&�q�G��fbV�#.��	:w��=�A����P��m��4)�I��Vk��Q���)m�}F�k�J�\Cp��\�!���)܊��]�+b�z��s"Q�3�o��<�.mAil"s���Ka��F�a
�[z�h%yA�Z�L o�-/��;�2ֵ���Nw��.��~��S�u��$�7����r�=����
�r}��巵4f8�^��(�xf[�i�GO���ڮ�����S�������{�n�	A��V
�w�p�i��}��2^�7�L o�X(�i7���3��{�a��D�`b�3�7D�9�>D����O:�,�ē�ਟ��9?p�mHCUiN���w����@��I�Lo�,�NZ���dl��^��Y��iZ{w�%#��5�>��v P߶ڝ��|��<�&�8�	��m�p���{�};�D;����Rd�݀�03���S$�'kAՌr�i_<Bp�u��յ��0�_EԸQf��M��A�*R[(���8����\͑�nq���fXSn<��6���R��(L�<�<mn��r1.�C���zv�g�[��M[���9t������\�Jk]\��u�G��|�ٖR#c���[ț��xb�;�P�(ﭼ+�f��v
�e�Cl}
�v�����Z�U� wj@p�I0k���Ց����W�0>Z 
y-Y�CVS�0(}���&�F�k�~�:ss�b^/�&CA�H��`E_m�O.�bkPn��矗���5�w���Ƨ��8�:��O��@mVb�n��7N����c;�.[� ���|~ƹ��h�g�qQ
�@���{�qWl�3�����j�N��( ����m�3yړ�R8�v��!7�}�e�� �Į�s�_~�����R⢆��іR�7xʅ@�Y�(:��/ե07�E��n�1��2(<wY���:�\���J�3,y��S�t?�0s��,�f�%��<s�/�Gƈw4
�G�K����mB$oXC���������;H��q�cl�jKM�1��<�O_��y+��q,��j���K)�;Ak��3&��5�$�J����KNn�s}'��,�oi�L�%�t�M'�,$��=�Н��8��m��7T>*�(�{t���,`�a$�C�6�*K�	��_?����(J���C�����%�]gRL'pq;^�2�S�ݿ� 8��9ȈAo�i��X��^XĜ�����9�!�/����'!_�՞�3��X�)#Y�+��r�2,
'\#�q���J�2��:^wtw�X��Z��~TE������`p�E6� �芵�8K��@�Ce�G��?����-ɧ�Rq���-������ K*�q���Q��'kñ��8�l<�n0��rd)!d���K�e�%���4������W�b�6W 4J�����d'O��#�
�1*
vN��lf��'D��?B(o9�ʹ�~�Q��B���Z9�� qc��F]�Ƣ��+�n��=]�Zب	!|c�#*�>Ou@�O�@'ʸ�\�ݯ�����+�k�|�H��GBq���x�Xb�pz�:;���U��6����,���E0�X>�lPѻ%POυr9�}��ދ�Dz�����)�KJV�f�Y%��ES+�nG�p��Z���lx��7+�l)ǀq�O��M�z�l�9;��������W���լ&��gǡ��	��`��h�*��BD�*<]RpA]q>`?�oj�I��Z1fh�����X�������4���k7�>�\�=��<W|t�����b:�^.�J7a�_�f"��6��m��[�tI�������h*�<,>�)<�"A���~%T�PP4���Cĝ�|⦚�����ZdLf�P���ƍ/3��^��b�T����n��L� ,��:���O��J}t�4���g��(�b�r�=p�3�I�f6��	+���#���0+�-d�Mx�'�ut��U�'���Eû��<T~�·B7p�@�n����+��j ީ��%>k��t`q�"Է��E���O��l���|i��?�����$]��F�`�.N<?Ѹ�Ő_�&B�Y�J��h�-�3��p�,�ߊ�۷�<�τ��ĵ�%��mCq��g�حA��Q=��whI����鈟#5�R���U��M�%��p�j��^���r懊a)�A7�)Z��XA��yX�x�A���{t3���X�G�w���]g��X����0�7/�,�1�#�p����c�x2��e��k�4(X{�QX����E�m�4w������eq��[7��^����5c,�� q�P��	B�u��Fk:`_9�%?[��q�AM���P��s�P�y2�s$Pf��r��h�Gêd.������A-o#7�8
Hh`A=��EV���H�da�61c�+��S�̍��̈d���:�4�V���(�\�T�ZL���k�+����z�F�\��
�L����,5#Y�t�Ë �m��kR$����V�MwE�Fn��ΐ�"��j�K �\��4���m���e�7d+��	�q���bE?�3C1�Z��p��\��"�qaC�ӑ4�кT�86�,�=���G[��7���5��8��ax #�|��<en���	z~Y��k\��\^�ۙ k��9��ϙ ����ąf0uc}�3�ݖsz^qZjA9�vd�_�$Y+�����6#��2^���.�z�����`�]�ؾ'���p��az����p��ձnB���M�b�#��`Z\o3F��b��4 ���BDE4� j��l-�W�,����`t�B�����udg�8�sS:
-R��g3:*t����h�5�M��־�ڱJ�B��edKX�U��]I��:'��df��(��$�Ul��o��#��Yb/��bJ��M����䥍*�y*��}J��ȇ��Q��1���R��5��H5i ��7<��r;<���`4~�,#
�1®b/X��[�t.U�s�Z�R�J���w�B�kO�?��0�Dt~I�0�������,W��6�#r*(��\�a卦 r�^}�]uũ�0�S��|E<|�C���*��Vs_G�p{�s�+�^Ĉg��"���Ϲ��(����i��51𽦖jcX�t�ad�*'���\rݖ�hqm5"������e�A�x����4/�aGF����>|Ǆ�B1(�Y?uu����l)�7��	��z��흤�v��{�]�
3�4x�6)L�@���~
��M�Y�V��]��*h����N.�Ai���s�4 �t��j�0 ��E�gFnH* .����&�f�[��/w��ߓa6�����"��C1��T>AQy���G��)p��9�����5�N�4J6�[�6��4�f$!r�o�,{��\��e@|��s�M�w耍� ��GY��,��p�z����A%�p��3�]��~�#���xr;~ךB���ԣ�Y��8NL�:2���G�w"���Pm;G���-�D���&�W���BO�Z-&�[0�LH?���ظo��Ih|��:�E�2��m���6;9@4���h��"!�~�ϋ w��M��۬D,{���.E0�ۼ�_�h�O���E~L� &���R��ծU{T�G�zdrj���(��}����!r�q�T�oL~YR�v�O�):l.��/P�ʾ8���#�<:^Bb'&�K�U�G��.�RwX�V&�����-	Y ^�/)�<@r�$#���t?�Q�H�L�%)�_zA�uT��@��������?Z]0�PG��Cn�b�똀'�][Z�b
m��C��z�aTql��y�����TS���Fq<i�M�8yrF�q5���m��hx�W!�)U˝����͗�md����z�,������\-ײ+�O*�y��DOs�, ��Q��p.��A?��{P��[e}B���.���v�.�q�J5a$�R������lSJUr'20�9I_w7��VV��X-���);�7��Lju���DV�b@�D��l���{�O�$cC		�Ĳ���m~Qj+[�r8�.�7��V��0��j�ܶ��ӯͣÒ��5�Jˋ�W�i��׀����`�u��R���V2�a2<��
0?"	� �xw�-t�5ym�����7L5?#r�x6ϟ�Iu�S����S���}ON�:�Y�%WH@8�����:��u%�Z���.�>��y��O�0��nT�#H��}���/j�5�0T�������؋'9�������(�T%3{��Q�EZ�S�b>ے�Jd�撾�^�z���x��r�dӘw�e2��r�S���4���m9f��v�9�o5���d�v[gw�!M���fd���n�����/�}��oi1�5�N)07�����8�I1���j��fT�NA�S���w�j�?�ðٝ��8����z��m�¨����z��m���{��mm	:���	�i��5f��453Н�ny�#�h�}���>�����o2����s��"�q�@�ł��į����Jpj���fY+ػW�Cl:�/�*��'S�hc��+�'Y~��"��]�n��K(�@��u%�%�ؕ�����;�e3Z�,v�ev�8�"l�l�C��e,6��,�*�<ӗ����*��K��;]9g��tH3�J� 6'��"��q4C���ћb�	�!��=��ŗ��w�ƅ��I`�xxu�&�3]mޢ@�e5�����XU���?̞�-�=���ᒮ�;���Gǰ��p*	��+�W�B�̩��B��\��]l@�B�����;��G?N���9/<�T���O{&��CA6����~��>b��N���%ÿ�]�F�')O����4��jPJ	Kyؤ,�WvԄ|��-n���j�b\Gk��$�R�`�J_��q���s��.9�h�"I�*i�G�)v��	ݥ�d�[�^�<�$�\ڿ��C-���R1f��pg��-�k~�v��H��yP,�FU�P���*g���4 �V��3�{�M
���_.>���;XR�*I��&�i@�����SL���e���^ۋ���$�?�S�cN\ػjj�R��h�i�p����i�s�|��$�Lj>=?:���[ K�����6qx8��CW���_C�_Oͮ����a���#Z�-�._eH�+���Y="������}Z��7S����+g]�s)а��$��A��	m�λ`gS��a3C~�k�U��H�%J���gφ]����w5���yg����Ӝ���p����oO�%�c6�Կȴ'�Q���*F��7k��k��ƇE���l�Ǒ�	s�N{���ȇ�ӌ�sS�L�4E2R���F"���]�ȿceѯH.�d���|N+�_��Wq�&
I\��b�!�K�c4{_�Ny����,A10W.]g�l0@�1f���_�� �*����r��ܲ��I�|�W�5V#Y�����v��	&�ɲ�G�H9�(�� ���lͭ���R<���;1�����Z��h��� �hur�����N�0R�$�(�������ȇ��*@�B~$��o�u��d���V�Xw�:���7����7�JwĔ�$;��R�q��=IM;~}�j�%c3��F��CL�� ��r� �?O`:����J��YM[4�>�Q���eeaH8B%.X���s���YŁڛz��2}�����.p��WJ��*�J��t���߮|;�є�p�K.��)�Zb9lTUy&
+�FU.�d�nPZ"�f�\UP�s9�<��#��Ԇ���u��⥳dg�8�O���������]$��w�3F���ڒ��K�2Yf��I�T��
e���a*��".�0�83%1 ;X�>�� x��!�_�0��C$����u�4�������>�[pH^�%B�����hy
�(�}ot>s�d`q�����c`еH��_�U�&����\��{�2���4��շ"ە��%v4mP`xB�����h�g�d��S �!k%��}�<�D 7�s^�	���������7mk�j-Qw(}���Sh�>��t�Z��e�'8�-�l�Cϋ�Zc	L߆�>,I���*f0̇������i��:��\���ݨg@QO�ѢCR������`	,_��/0��y[�Tu��Ab0_>����K=��[|'��Ͷtn��=�E�x)�?D��� czO�ݦQ���Cw<�6��G����h�8��J}��V�^��t��ܝ�)�d��m������%�jo;_M1��F`r,͚8V�f5�h@���wNFF�y7��BUhy�/���x������]0�o�w�4���MV</����tĭ�O�;�X%�0P�k�-k���0��F�G+ع>���Q'��A����(��
b�p5��3B��W�۽tC���A�1��Rm��K�� ��{s��ᚻ>��j��G�ρ��4z��S�IG����[#/�Z��!�śF3��A��c�)!!5^@29�Ӱ$�@|8/%��~��4yA�+���	$y�4:e��{xg������L2J��W8�z��8�p�	�"��j�z���~^Ju��d�&b﯌D�J�G��}M|��s�q9�H����j�Ԇ�����QKU!�Kf���=�4W�0�-Cנ�Lm H{���� 0�{,�M �������ĝB�t�Kvd����0U��`_��t+����Pw��ur��|�T0y�� $�W��Se҈��>�X�o�/�CK��1������7�[�|'��]��}[������吭�)�$��dL�+Sc���hʽ-9+�H�>9�'[�0<&�Sψ
����K�eKI3J����긧u�_o?�N����}9�0}[x�Z��=�m��<�����bN���Q������!�/�6��GAKZ����ؒ����Hq��K�T#1��4�e[�1�*I�Un(�����r� 	m�mؗ����%��#)�l,�|�JF+r�sj'�>)(�k�@�C���jÔ>|�<)���t3�d�*�}I(s����,�����E���ˢT�$z1�y���/�_��s׷��`�ƕ��q�m��4'�g���a�g�������(G�x^Y~��Pp�Ax�i��|$�mH_F���]4��u?����-�RZ�L%?�B�� �;�e&r��9y�-9����c��q��k�	�i�͕7�����˘�
z��Q��/����ǣ�_�����;2$�U��k���՝��C�s����_\�7s�-���<�����Gj��]���M����ʰ�?W��9��8�4�8�����>äbS�m�p���I����y�^C��vyX��B�����U�g��x&���(��=`WE�u̱?۷ �?�叁��{U��Q��C��oFo8���Z�#i��q
����s�;�z�U!�đ�3V�����,;>���|�ih��L�����PV�;�4�+j��e��Xz����)���3o|�Մ86�|굃N
n!��N=��t$�.����a���	v�� 2�#% ���
�	��B󁺫�n��Gl$�h�}��^�nY7���!��tZi�ST�(�����W�E�k)��Ɔn�C�2G��U��r����o�� _���'ۣ<U�X������I�<b&���XN�_�V��3k�M��Q�Um?�>5P�d�K�}��U�u�� ��9�R@�Y���&�5��5$P-��WD|O�Q)M��{���TR��6�4ڌrT�ŷc�ʝp�j�e�M�g;��'�XJ�?m���A��cr膔�5�!A�|�;&��/ڼ ư�'ژR6Z��>3��t,-���r�Z`}�ʀ�'޼�]¶4>,�f�4R�)T��%ύ���M�[��B ��uY�Dy�Ȫ��׈M��#V�}���z]�I�Vj��W�Y���i7��f��k)`��S-��"�	)V��|�KE��Ń#ݤ#�Wv](ϙķN�!`8?�X�s����,$���rr�ǀ���^�x��/��!�U����u�ө9<YYǬ�M^��*���IO�t��O7#�슳���1if�X�EP���q��ݐ�]2��m�V�?	�>���s2u�M :�*{��^a�?�$8D� �����N��X-!����la�6�I�%S\.N{����w˺ARls�8O��\"Z�l��[q	������^
%5��U�6:���{o��^/"�ڌV��!��Q�3N���5�!� �����<@��M�zB��/�Ɂ:�Z-�H�\*���5�R������_m\h����Al��KY���õ��y%&��w7�\�w@S�}e��5��>���C�EfU�@��mbqT����*���QćR�!�q9#�g�un��3h�@T����c�L��p]�|�Ț �;��mA�Y�w����]��o{f�)�rЭ�M��dVt ]wW�������SgR�.�ȣ�(	�F�TXk�$H֟+�IN���ّ�
�B�O�)6-���	9;���AY���و�^�ۖyJc���e�s^��I��򪐑�k*S�5��2|ۏRy<�<SkL�4�`
�����~	����\=tV�%�x'�T�O�3޽>�w�#;�<����eF�܀`֠�rzi(�Kæz����,�	/�#0$�n��@�N�-�
t"&�g�K�Co�T���%���K=5���dl����i黎��7����^n�����۔��7�ݧ��8=d+Qݝ��x�j�uT��#1G���Fd��*�$�N�/���������d{��b1!�i�1�uhDt�a��>���7�w[5����z����Z���u� ��ܫ
"�T�FN��|ؗ�.���{;^xJ����Ė%��
���q$t/>��'�^_���>,�v�~�?cS.w�������nV?!��:7+?�!�$l�,��o(d��.?m1��K:�B��d���C#�kȍ�I�\�3-[�{�rq$!e'_e
8٤��v>��	���2+s>=gKx��W�"�FJ3��Uh��y�ԭ�q�TC{�	�[GBbc�~��3�M�\^^�E�!�3~�R�Hi61ц��t�y�!�QNӠCd2�oڕ��i/x<����^d$�T��t#��n��'��T�)��|��t�T�^i i_Kw��)�>1=-މ^�^�X���4-C�x�|�b���*�'$5[��Y:���]3+ Ƙ�V��mP�F�xRiy�HJ�􂕢�LG7r-�Ɨ���y��=�6�'f=�%t"�/E�}��~ε�v]쌗1���)5C�q�m�i��w|��j�= �q(W�V@q��5<��ʆ3^)a`�K��{������c�Q�G���v3��Zl������Uk�ӓV���|�{��8gS�"�!?`�8��z�F��u�rj���L�~ �$jH3��\����&g��#�t �25��:��g�բ/�׾X�U����eC/<I���1��{�_�v���-e�큰�D�_tA%��Z��_�^e���Tρ�
�C�U���MT�JK�n9�7u�?�3�[C�"0A��5(���Z�~Oo
)��o�w��l��Q��DGb<0y������%�i#��d˪���5�����2�ټD.n�������]f�@Q���ٮo��+��`���G1W�H+U��6Ԅn�1-�$?4����5�ڙ�ʩ$��^+<��V�L�ÑM��<���Hx ��� R}�C���F��4G����|eE��82ˏ��N��=G�OtI�Q3*�w��?��
mH���P��5����MDZ�0r�&��GŘ��I
*y�o*o�7��o`;1�'C���gc"�Ǵ��$2�#����[��0��n�"�F��=�όA��ȸ��T䵑�ɤ'~���Wund���d=�Gk^�q�xߩ�wy����e����AL�Ə`����ڞ�t��o�����&��zc�iNG���}4�l.�v-��O�$b-����3�Z���s��7����$���u������,e��\��gx/��⛇EG�`L���y�ǢR	�Q�Z�g(`�����ԶA^�AP�<�#�ǰ��0�M��E�������5&�-Ѡ��ڛ�T��K:�3�F�9ŕ�y	��A���T�h���U�YRWA���Le�������*'م���ʃ��Y�:!F�)�T��6��V�]`�I�FE��λ�ĸ����W���}�'MDtL����bM�3���ǽ\�g[����h���L�<�]��l`#��o�����o�y�� jL�6�M��\~���5�R��Il?
^=�N���P ��Hk��N;Ơ��ERR;��l`D��?�X�V�k�Y�s0����2���hѩy��d��#����հ
 B�	�h��d�O���78�>ҝ>c W���s t?�Թ�Y����ݼ�ۥ�I�vE߱�?A��<p�	���|�Ą���}f�@��Aa�,b�iA~H����E�6L�d�R���ϊ �d���� ��yM�x�4���ϻ=c'_{���*�J	x}��9�pzk@zF �������Gߘ[�]�l���2��'*@}8��U%W據�sj�X'K.ǅM�W����q%�ހ�3������m�uV��]6����[u��`4�Ɖ��]��w�WY�'e"hL���Ї���]T��
�������r��˓�H�%'��cz}4�:�/�e��19��&�nPG�Z�6����[�N��ެ9��u6D��͑~��̱�����r���S#X�Zҷ5���;b���`�fbV Z}�]tR+�E	�'C<�{x���DiHhz�x �Dk�\��w�Q|w�?�@`Mi��j��Do�b������qB�+�ZzR"��8�9F"6��HZ�Qb@�"��� ��S'ƋΞ���]�s�D��Ua�xЏ8�a���[埙 Z�Lz%y������`�|�,�w{~όן<��=����m��8�q�
�F���v�T*g\��1��0;��� `=���،��iz���j"��%Vo�_k��όᱳ��x�0��0�$�Rc�g��*�6t���م9�)zCz*����� ��+�Eb)9m�W�C�?��bI�T�]d��4/ҫ]�\�q�\��i�l�'a�,�q��%�O�H���*�u����H[�?s�ZBn��R��84�t��2�*6b�m��p�У���f�թN���dZ�0���haCQZ����ӣчI@)]���yW4r3��{�5���\�������"m����D���yG_N"�T9��-�ǥ�p��+/Qr޵�l3�X5Ar��l�9V����^RI����T���ޓ�Q�'3O��e���X�9&�RP�y�����<cM������E�����(R>bz֍�<�b�j����a��F-=9iEm�M�x-�k��񴉸;�v�ͯQS"�	z��'�e�Vu@�y֛}�YW��\	��/����`h�ȾQ�i�hk��w|`���,�8�i�iѲ3�Q��/�+pm1�䱚:K�^Vg��fy���bᗣ�M���M30��9�f5#a�&���G{/�ΗP� �0��r���2D��FS�B��f,��5�H��I��	�t
����y�[�������R�f��e֑�.f>ޡ,�b1��FJ��x�����?�Υ+���j�i�3J~����o�V�%��=Cqz1�2J.�o�1h�?3����
J�Q)ya�l�_�����_U~ߦj8o?s����i]D����q���6���kM喦�!ف�1a�B[���	9��4����x��c��N/��@]ն`���nrI�Cx\A-W��t�*\>����\;zR�7�������
B��؍_ ����݊<C������ϰ�����1�L��rV�M�/7�N�zi�@�b~	&���JQZHB��ho��3�&����)�j0V|V4`�zQk����g��%��!�:����]8 �ƶ�jqh��U���3l�WVe̼��0{�����2���]�RM���g�l�3X �I�]	��@��%mQa[-Ԏ�?A,ͧ�L��Uٞ������M�g�<�"�KWk�2�����i8:V_�8dQ-��a��6�]	P2$�5,#0e\�}*�ꝭ��ik_�{�hLBNgƻ���9m�b�o�{3������n'��i��h��Or���i�Q���~qAv����đ)P����}S�{	(>��x̢�OɈF:{k����ָ�W�o��T�H?�����hy�z�_��荄^_ n��L77�ο�(��4{�j%-J��#XQ0#H#��F���l僧�>��~��'������ߜV<��km� ���]���y�������U��e?����.��\��W��P_սᒿ�%SI�j�|/~ǋ���f�ٱnM�|�@�W����&/� ������n~�(��>�XqęB�O�r�+&l�yZ�=G�x8e�\�_��j;���Y��e�ެ������y��x���ѷ��G׍s��/R���.bwia����ͦ7�0�.�A&���:1�;LP8ٴ5N!d��Mg�c�4Fr^f�uٛI"%�¼3?)`��w`h�`��9]�ΡZ��(N�U&��o�4���s���tE-��;�I,��,�	��ۭ�vV<-A�X��c��u��R7+�{�D?'Ƹ��*�w^K��`�IS[���o�%�H�N첓⌌d����@X𰦄��3ą�cI��CH5��,S=� &Q�t���o)q�˴b`�E+}��ܖ�\�I�6�_��(���T���$F/_�t��RT�Ik�ShE O��P� �7��	��AC�B�=z=�\�my���5����Vp";�2W����_+�����|�~T��A�R��L�S��D�KH>Z]��'}&T%�BG�qg���˳�ܶW �^)�J��%�ے�U�e4\G�+]���Kd|Uә;��vrۚ�s�<�Yw����L\�n�V#�63p�ST�����w��]��>j�C��^�֘�%Q�R�������q�v���lW�o��*Ύ4��^�\�8@�ɺӲ����ƖNf��I� !n�>dω;�	I��3p�+(��Gbb��vI�7��̋��j�XMB��wZO��v�q�	����?E)s��JM��%����J��M�p�(O��7��ß2�U�Ȑ�k|��%s� �u�b'��>����˿Q���A[e+:���wT�S;òi��6-|z��5a\N�(9�-kߒ'�р1��f���V�3��a�UZU`دQo��ݬ J���F�↊<�|tt�}���K����ԤÙ#�)���p��!OdS��h!%J�-A�/������R�b������:���z�9r*n�΄Ĺ��(y�UxO̾ҧ`���p�$������M�q�����l��
�H��������`�� Rb���r��f��N�P��B9�R��+D�a��y��!)/]:l���6����
%�L1W�&��av�F��y�VM� �����U��烂�o�Rl��zP�� <�_� �\�]�c�a0����M��Cx�gn�;�24~�#�g�'��J���&�@r�*�ڜ��?�0I�FUc��k�wA�Ϻ��K�}���Y����C��9�M,�\$��nLsRp��7bԆ����;�+����6f� D��+q��e��T�t���yp����6�uF����?zh{��ŧp�g��ܜ�eH��w���0�F6��؇SO�L�mg�ti��?MK�;0�� �h��K4I��Ǎ�#� ��4ƭ�"���P�7n��1E*�R}��K>�>(+��U�2������
���$2ͻ��k��
�Ʉk2���H�Z��{�T�Z�ٰ��d˱��L������W�e>Y�{��&U��,�C#kZ�*�̼T)��j�A1FQ���c�5�niL���:~�?CSyYr�Ӳ��в:�؀�P�����O�e��=�əT�Q�ˡU���4��ڈ+_�����ߗ�\�������d���)��;�m~�::B�,��X���:w=�\E	%|qB�2�x(+���ad�����s�7�zZ%W��t�z���o��Gm6�m{�D'���k���]O6{���D��G-yd�zl> �1������}[�9�M4-EnZC�n�����
O��m�w˗���f�$RN��d"L@;�/yT�fɢf5��p���I�? �k�m�󶹤T\���i	��$ˑ�� ���zrLJePۤ�r!��`3��`�dM��&� �fr��j�����t���6����Ƴ4����ܦ��Mx,ҧ$�B�y(^�Z�9e�� '�c��Q"m�I�5���,�|��+_���򈈿�`_��3I9�����r��Kx%
u�cp%�v�K��~�-;�Q�ǚ/|�*��&d�\M�#k�"�XF�FW����JD5�I���k�Z�3Dk�:$�t�9D*&{��Z��muZ�T͋x[���)ouh��݄�����W��ص�UB��;�3Y����?8����1�bL�J%���Z��[��l�Б��򔞃J(>?�9�Ձ���;�:3�Tq�E��\����4�h�pA]��v*�_{8����i���I�[��[����R���h�M��Ý-�`�eN~���<�%c�������i'E��G����:��g�\n�^T�4
0;�'.v��-�ނ�6��~���:.;��k�z�л��ؔ�(����1�6��.g�Lލ��1Z?���H�5�]Е�� ��*��B�y����Dg�g]s��Ac4~*�Z���&}M�^+����D���Y�
�.�V��=��=�rRh����OR��h��#�[ɾ|�'���v��Z�k��8�G�]Ӱ�.�����.V��1{OM������������;����e-ٝ^�nOu0��UĿ|��L�<i(7�T�$+pw����
��}�܉�@E-��Z�e򸽱v~�T4V�V�ĕ}�lD�T�(n#������C�0��@�H��
OBr�F,��s��Xs�Z:jG. ��&"^���|ګaʗ���e����W��x�%bD�Kh�c����|��!��
q�5m.��\��@�K�L�,[��YK��P�3
�@|��]��|e�_q֊��}rr�*�9�*��X���3��v�0�0���}~��u�Ѩ��l"�5N��MRɰcˉ�T�TU���QM�>�I��,�
���A%�NƨҌ��Р�CU�VB���Pc�#`�Pzd�K�&P!��;x��fM19@�\R21��	��[���Hm}�#�0~�ҟO+�r�	�?�����H�'�#���M�R �#��դ��P�k�����	��F���I�PI΄w
Bx��rg�t+�@����*������*���E����fn��?s�D���EW��2 I��&�����5���`a��7�4����:x��S�H��\Mjq`+�!�wҾ9�/F�0Fe��"�ϐt*�q�"$�����F:��/�E����t]���]�f�Dw����BrM��������Ct��^0���B���i�0/í�y��*+O� -	�Lb��_��%c4��>YF�uq)��k`��z�O��W0���r���l�k(�yI�N3@T�}���H�̔��vc1�2	����_��f�h�5^x��³�0������4��<��3��I�f�ռ5KrWY��g����<=����U����\��z� �<�%ds$����홵�$.�Bh�W���T	�H�TA|�Y��رR���Αf ��[/N�X���3����K��O6E�?vּ/_�]�HSМ0'����E�#~[����n���e�槌t��g�t�<��6���Z���&2��Oj�}@L"V���m�io�����8 @�
�<o��.m���ɕ��'����#���-W��qoB=�ރ|�l<-�iS��ki��|����f<T��_-5�K��
O7I��s�؀dʔq�zS��@l[|�Em�u�����s��H�����lD�?v�"a|�����aN����ڝ5�(g���j{gj�P��}��޶/N��XFQ��r�1�D=8$�V��~݋��Vi��J�XQ�����eQS�� 1�-�^�CVv�4I���MSs�,@Ӌ�p����n�ᗐ�K�'����-�c܅�Q�t2�fCI���i>�li��m_F��"��SqÁ�B#ݨ��l6P7cU���.��ud9�}G��R��}S��{K���:z�'gD����a��t����^b(@�n��xp�QC� ����dؿ��/����iJ��#�`��{�7[,�Ȅ�A@�񧛂B2�DUTX)�W3Tp Y�d%�w{3� ��(K�N�����Դ�:��.&����<��K��!�{%���N�����!�����*Z�"�'m�08ѫUu;�JK���N�+�
�v�~=p��C���p�X(���Q��{��~�pAB��~5g�Ú+�;�c2�;u:�L���7?-��缰��i� ��!��5��;�x��͌n[���X>`7dhN�#C
�<���&A)��O�Hd��t:�R�8W���M|nR{�5G]AC�J��c( ��=��^��
"�(��vk&i�e��ʕ8���ug)�Dx���$|��������&Ђ�{ء�S����ۧ�Ø�S�5�'i6u�}62�Ѳ[�-��o'׽?X���+�xm0�޸4�Q�l
����PfgPju���Ɲ"0}�M��4�=�ONs5B�A��2l�t��,T-d�����+�o�����ᴝ�3�,��x[9kv&���MP�*e.����:��3%���6��ķ�l`ϿXӒ4u�/*�e�1}�<(zu�6'�i@�9�~B�qLFx��.���,]�p)�:G�+�L,�[�J\AW'0��<��bo��Lp1�J㑀٩у�A�#��4 -�l�Sؘq�0��	��.��+� 5I�Q)�l�������zJ��|�z/���Na�3ٽѴK�j1�X�č3��rU��|�rQ�e�ōmE7S3�U��f��7�:���AB'�K^��.�4)ZR`�"w��2 �����}7�����Uﴬo�(fꙗ�<�f��.g��'�/7���}�~h3�_�6I�W'�UjLN�,u$6A��g�k�6!}����{�hT�h���2����%��R���SX5����7#�3@Vx!5_�&��w���;��F�	Dß'�
���0%V�q��gX~RS�i���n*�]�azq{K�+v��o,%H���H��=��Q_:`��0s�;�f�؏��J�u�)����Fq��!�L�5�&y
Z�}�C����4���nP���m		�pi�T4Vv��=ލa�;��B4ԇ��Bo��!��	�"]"�+r28��H��_ώe;1�~`�)��=���sU'���1�M	��(Ad�d?�V9
��˟L�Z��ϴK�sz��^0ոR���پK`wn��?X�T� ��j�<�Y�3�����i�l�ms2X*mJ�&>���b�s��D�$đ��Ĕs���~H��e� [�ǓCm!���[���( ��keZg�7K���fa9��ĝ�C[�M�7�s?׏�	���P��wE�pEVo�`�����fo����ՙ�c�T��F߉D{���nG�p4P�xV�ip����'�P�k�a6y(^�tfս�,��]��Ǭ.\��Z�����5�N0٭���M�	� ��/)t�N��;�D�u���,�}xrO��h�W� K`�V8{�ޭġ$BV�D����1�	������pox�4�Q��(֦�B%j���/Q�8ݽ�tk�a�o�s�)��f��x}�Xv�s�"h��|��mU�7�˩�Ǌ�bR�0�D���l�d�Da�w/L|���N4}�?*�2o�s%M�'�I�߲O�"��Q=E'o�23��-1�)s�Vp���eM��@Vu�m�,����ځUe4<C K5хhA�;Sh����(��D߫��ܢ����ܫ2��6� :#��"�*�����fXnG&_b�}���g;� �#��o����
�Co�)F�Z�� !����k�#7�pլ�	r���-g̊|�����U[�u ��\e׭}�Q?�#y v�O.K3�B��dxB����!���)#Ǧ6,@iT?��О�b,�{a=����;cb �=��-�솽e(Ւ�h��b��zj[\
?i�x�;�q^�b�������
u�Hx�X� ������j��2�h����]�Mw�؞���Dfni�,O`C!�C�rU�g�M1�(�=sD��g�T�L�7)���W��ܛ|L�ր��}Co#۩
�by�j��-\�]vfH�Ahk�AM� (^bݺu����zH$�Bi���]������C��{Ƶ0����U�С�,��6~{�&��aĽ�:�+.�R�oy�V��f�C5Qz^l�s����	���x�qy�!t��d��ʀubN<ȣ�v�ᵘ���	�ۉt'��tq��;����)uP��>�e������s=s�"�R��_�x� �{���G��&���֋��i��R���Z�%}R\W�^Qj���
��am^(�T*RDJ�"�tm��y�ʊP<�YZ%�*�Z~L�R��c�(F��>5��c�Y:w.��\�p,����rY�����\rh�z�T��S*�8=�_��k8�����m��*��(�/�+�D+@GQ�)&vm��dBy� �v�%��<p��14�vԧۚt��/�T�P�^�\��䔷��=(1���)91���V =��v�M�j�� p�vˎ��g���Wx%��b���,�b��M$	��Z;��	�>�*N�!B��ד��;��^1D��)���tŎ�2;�n{L�D��}�\#���x����'������Q#Q^�9�N:D��2��G��d,��Y[#�@�A$԰|��蔫�x�V�)9�F�mWġ��k�Ӱ߇�ޜ�{��ܕ��� �T��흲vPU�_A-�߮�~�^h���(���uO�a85l�����g��]џ����P��`�Ͱ ����~i�θ���M��wo�KR��m��e,��"ҷ�o�Lg�k�S:Hc�KJ��-�ԅ��l�g�'>g���߽4�ꦲ:��@�����s�u��#޷q����t�T~ms5�y�APY�B�~���'���j?�u�C��L�	�g9fK���<�;_p�MV��L/J~׾�]��&Rt.�0�
W>Ox���B��˔��(d�r>�v�模���r$��T�k[ρ\�є:���	�\^'�x�y����L�g�+�P�-5?Y����0g���GP`06�j�Ù��"H���h�l����16� ��r;G���Z��3�m$���#I��>���"6�����i"�wgOt���pu���K=L��>8��΍��M�Ү��j�ܬ>c]i��k�o ��X++���֦
���/�{猎o�������S��h�:x�5��3����i�o�
�D�@��÷u1��\���	�.5���4^��>/�VGF,s"Nٺ��/���Ǯ��ܪ�=��"��(��Z'_�CU�� K���
�6�� ���wݔ���>��\��]�0���ZK�ԯh�?��=���[�&�W3��7��f���(�k�=�\y|J�F+�y��5$���Ƨ�����GB�ڷ9�p��00g|O�y�`9T�Z�	�+���A��Kr],ʗ�?|ß���;�*py �WQ�DB{c�ŲJP,0��o A?�Fg$Ϙ��B�+>���ǜ��{eg6��=��Jܠr��W+����ّ5�������e*ɿ�k����ĝn��[XFF���=�d�@��r�>���Vy�W�M�:�m��}�&������\�S_��7+�K��y^/���2�[����8��Q�W�Ԭ���_Q;�3J�5�5�a��B�-:�cUT�a��7p�S2�At�V-��r����Ds^[�m��I����,���j��r�Bp��������G��aq�IE_*cC�A/%h�p�[����8~-$��@6A!�|�с3T@�5��J3Z���FD��gf�v�7t^���Ӫ��$���Դ���[���Kg�ށz�����RÞFɧT0<v?��7��mbXr�Y\�ȱUFR���l���͸�I��)Y��7�2���O\����w��i��M����bqVz����G��1@�\Dܜ�%'�èc/v�%�]X�k���N (#��6dBJZ�sIў�&(ϒs�b=k�/�l��-i�������Sh`��D��8������t��s�z^�g�%�toSq���6�E�uLAߴ���x&��� ��i���<B����$(�e�3-��E6\��c�tq���_92��i|�~`ǳ��@C(�S�؜	4����>��3����k�Z�W�yk�i!�����2Z2f�Y{�l�]5F���EU1�E��Rs7(��%ŒD��2s5�>5���>���TۣB9a�k�O��z)Xh^>�΍.�V�e39cڏ���pr8�=��:4��A�;/f�8�rJVaC"�Ƒ��v�������Z�I87=��g�ͳ�[��3Q�(!���3D ��#�"���o��R5�W݀|fX�˼˯FV>Cl��-�0|Q�,o5+;�8����������,�W�.ؖ/�~�G6dH)�%��܂��tW�*��ı��~���j�Ӷb7����AZ�)����j<����۹�U�(*V��Ԥ�����>�y�t�,U�s�.2w?s��VK+��]��T���=�H7Y�':��V���_e*��a�_���x�2���?`f�mH���z�HhG1������4�����	��I����;�dE�mcA�}�����Y_9iN��(�	���S����jLE�#����(י&�z= ���Sl���
�B`���,uA�cE�zJX�+�e濃�'w��`Xz��`ʿ�Q�!a��5�+ݗ����M�-�C�)��������0K�C�8=�m�c*2�͸ni�-�JK���%[>�+X%�]K�l�4 %�&U~����5@F�4��eY��$R4����8�"C͓�/z#�fG_��>Xiv9We�S�A�
���2i��o0~�Oh�����X��SB ����{�%M.���6�v�s���?�Mѐ=�r��Ql�Rf��a���5L�xxQ���5�d��+�6���d~��l�-���~�ņ��_A<o��E�</q`8^���O�L/I%sc� {)��&�����3���O��x1��8��Mql���(VZ��J#�l`�7jJT�X f�����������E���LEym�fъ?�A��)S'��efn��ME�sl�K���gBa/-"q�Ǩl��ϯ�K�hb�<�X�	ڄ������n=�*1����\�n�1~3j����.G3[:좲E�8����z.`�D�VnN�{m�\�\�i7o��u��.�����֚��vf>��Đ#H2H��*U ��d�<zE{�dC���՛RV}l�x`J��A9��E��#��d��nl��fV�]�<���E���� ��RE�U�C��7_r�R� b{>t��9�Ƭúk��wV���l���r�; H��i�����sw��^�{�cp?	���z3�;�A���D���?�v�G^NǴx^yjW��~.���^��S�?93�ؐ���X���J��P�LX�z�
�u�X�[����;1����h%��JoV��PP��vw����O<
��<KOB�M��4���V_�����[	���E;���������l�a��ϖ��-��G3�jI�ͥnQ1�U9������4�x��Ҭ������|SU�S�8O�*�xS��F"�V8�YN�h���b�8۲1N��$��\Z�Đ�F�8�v�5gJF���Jrl��-�N5y�z<U �'�$S~=cE�ӻi'�Y�9���c�A�u�D��>߫]��6��fa�}���'��!͉�b�@�P�6{���?v�����p����|:���u�'U+nU�y������%��uĭ�/�7�ʬ뱡��������2'�]��mC����F=ɺO��иCh��zhP��T�w���!��=1�5@�p���KR��@��p�:�c���fҢ�)����V�u��]ys�ihҹ��Eo�F������Y�Ò�^�4� n�a�[�*Jq?T���rY0�<)�Է4w�Gbj������7�.��8}����b.9q$6�Li�3���n�+�w��LSC�J��?��x�-�����}&Ǆb ���6s&<����g�%G�0}�������
��������6�Ĉs�(6�o���BÜ��˧������ˠ�|�F�@�-�~�Fh;�x��P �D���v�z�N��yPG��F��@1�jPs~�h*�ݗJW/r����tS�#ڶ�i�)�mB*�5���ԁ��`��+�H����"j�Oތ2(k��{&�#���l�7�S��e[c��O��y83�\�3�4�	)G�����.$�*��8'�<�p)0O�X����EӲ0�鳛v�?��(e���#! ��"���H�C�X���j��q���舽��s�0XMq|�[a88vW&-�Er1��`	����,E�e��+���t��za�T���p�ZMD�T=�,1�y��o3�KȡIc��^�sw�(��� }��},װ肹�I�4�+]�cq����|2�YD�g����9gVj\u��ξY���Xcg�V�XD0H�zN��+��DA#�FI�y�_�H�.���^����7Y�!�7�UzY���SR�hf|�ge��vN�=�i̅�`1-xr��i�9�7�.f%xOR��L����\�J�H3 ���]m֘��,���y�Պ�+�b��Ŵ�T%���Щ�*�C�JcDbE�I�4��]���I�l*�O4�(������c!n���e�\�q��ctd���K�FjZ��KP�3ڟ��4}�F�%9q�啒mW6�����g�+�XQ�bM%ŋ�a��jy��}�U�Ŀ0�^˨x���$c	��׽� �{�0�1���A�4쫯%������©�M$�v��2��E�sa�־����E�ݤ̅]A�����Q_�i�6.��MB��&��z'hUl;���j�Eƃ�揽� ��a5�_;��B��>�J9A��1J�}�����<\�/�g�ػ��$���jPv<�1�(�,|��C_�2��w��7"�$PlF��� ��A�ϵݮ�G{a;��ur̤�X������4FzZɎ�����x�m���d��n|2�S4�y"iȪ�:1aL�}���	)C��� KY�`pN�5��6�%m-hΏwj�?A�(-s����m������4���<�:�%�'��mC��B~z�!�Ηb�>����
G$v0�td�ݵ�g��$O\	�T�ԍ�X^���PPR��ZSGj ���.�jA{�����f%ɪ�mgޣ20�j(�I7����$:���$�����9s�(�߿�֚�3��ډ�����?�o.N��"���7�O�Z�7u)�@�@r��a����p��^=�[��*I�#Ԉ�����y���z�`�Nc6�L-��G�-e=s����]����z��.�lF
K���U�^��r��;v������Q�)z���5���h�7Ӈd��j[�{�:��K��x�������Y�s�������u��� j�}��m4U�B��&���[���w�B��D�,�)
ekK|�R���U�����P����G)v�Yqc?��P&H��Ț��/g���g�݋������Fc*,�M��z̹̬�/�!�/�C^�<�8Mޔ� 'c|��1�xy3�t
*�~<H2�!�Z�>�#7�1r�"G[�2\�[!��&��R���@W�3��q3�~�JF�7b=���,n���%B1Wh� 0�|q��#�f���qt�����M��c�A��]�����BiP�x2���A�������|Lа�oF?d*�-G��r����i�X�?��'�`�qO��`�M��|>Q�گ�5z�
j�}�����v��s�Y�XH���b�ј(�h�
��	sV��@ �B��h���.N����)8Ԁ�����8�������U�=��4�n؎��a���>�¤���X���-J�@�zTyȏ�:��Ƥ��"��{�(P�N[����v\��v�Ph�E$�0g�~mj�'��&�O��7�:������9]�~�N��䠬gv|u-����Cy,9íߗ}F�g�W�a���y&�xJ�aA�`F��i v��10N�����yC�A�Ɔ���{�=�.�K���b�$�t ����R��F�[|�NUuѝ�P��A���� ��'���Z��<��;�$�FO�xݸTBS�ƀ^��� �о�.�,�z�MGR�[25ʸ��F�K��q��s���àdJ��4�Tx�D�f����*w����NRՔB5�^ƵN���5���~��\��/I�B(M���`t��nix�� M;GL��� .�B��U>Z~!�@����2s�oc���f���?�Ҷ���s���<���&��a�����o��Ƒ�^����d���Yk���X������H�rQ�,�>@cvw�'���T�k�»�[������_��.������~V�tCM�Y���G^�	��lF�S!Z닷��Zow:7��½�/Pă����ܭA��yx:�l@���z��7�)E<� 堎
��6yi�8H���~LvQ��D i	N���K@��g:i�	��b?[I��e��ʳ
�"�!��}����t$��ڼm4���"�6I�uf#x�=c>ڭ�>�����Uo��,S2�a�K;�H<����SO�J�~�K
�Ά���0��ly��N��`����Q�A����zj��� ������I��&s�y ;g��P RawKK4�1-��;��z�u��P7w\��qf49�/�ɲ�V��} �c_e؏����8��s��w���{�'�f�Gca��I@,�F�jC�z��O��'ij%����؀�q��[)_�Y'����q�pu�+��� ;����}3iZL�wgR�,A1-��\6��5A�"�R���R�Aڮ��T���Z+�v��L!4`j�����suW��O#x�p�<�f�|Q��a{�3������SVzq<cG
6���LB�'c���	�ߣ��r�\��T�W�>$�\��Q])�h�C�A��#;_C��5�t�]���P �3�A�T��P�4��v����[(*�,��Ӭ��B e��w�C0�}b�㎨/�xщ��M��0�7A��]����u��5�C7C���ԕ�<�Q���e�'�C~d*���]�*�j��"�IUu��<�{�V���-O��	pS�Y�T�u�6�q��ù	���N3��+rs��<C�f�q�	[��;N�~0�	@#$('��1|^3Y��#C�X��b��([��goM���ڲ㚺z��W�^ $&���ff�!
���l�����VR��/��֥�%俱�,�)h�� ?�S�V��>(��YL��5��ϐ���K���p@�|�c#��6패
.�btZ��=�P��gu��\���%�C���2�	XTx���&uWm7�`�����f	�M�[��ȨkI�y1"�h�b�dRȃ'����ۡ��i��U���&	�j�swnF���q]R@H��6�2�����:Iҟz6�*��)��l��kz�TJ[�,Z�[8-7�ӁQ������2ǔ���
o���m<[��	|�WrsŇv���0��.�gȚ�۩�M�4:(G�j��b�]U�n���� ���]Ϣ"&�3d��q��]�8�V�
��c�>�����Q��`�&GC�[UY�U^����$�!P��8���ý���E�R??��N�"�eC�PzG��^5�Ң�zP�}@ <�"��{Z����-/�_r_�Q.��z(ŕZ��!@8���.N��vu�" �.4פ�&t��j��BS���s���b�|*��"ą[�Ԃ��ӨR��ǗYZ���l���.�j�������������io��|o��&��Mϋf��(�Zrҝy+�LI�_x�VW�?+^�`7ދ��0���^DY��*k2�����9�Om�����Ӹ�ڳ3N�c��/apa����X�Zo�.�L_���B���N7������v�J)C̼T"#��T���?a2ˢ�ȣ_��Y46u�pc��C� �&����+%�CG-[��>���m~'�v�)��4��X�嚜�W� 
ƕ#8`��d�O��b
��&2gqL^�mDp��N@��S���D*ݨ�ݟ�O���j)p.�ar� �A:=��pn��׫�>����^}g�˖"�tk�3nh6ȋ�R��-+��1�E@�79�8����_���x��s�o��랚g4��~���t��+!3(wXL9I�b}d�L�+<w&�-�B?�y�2��c�6ge������3����~I�mWi���\��������U�s���!�4�})Ҭjl��c����-j�WK�����t܈Q��HT�G��������r։���a�:+8 �,&��!���9K�gy	a�U� �Nw�G�B2�Uݎ�Ŝb���G��w����Vz��g��p�pO%��%�ӎ�n��_�+@ʢ�8�_'|gˋ����Ћd1ƪ(d~J��[$WB����]�|c�1׻}6�[MP�)�!x�s|=-�(�2)�
ݏ=��ʭ�:ŀ�pQ;@^x�:K]�!�On}��_�:B�9I� E =y�ٴjJ��قՎ���B����!7�h�T�C�;�3�\��AuKJ�u5�����c/��ū��H`�c�G���y�����x����']Z��F)�u��$����!�"Z��>��xZ
��	��S��g�+TC��g���h�G���C�փ�C���+��K�lz�����q��S�Zj3L����-�$�G f�����SA���|�Ë�=K���tA��}�����?DS\ۀ��Z=�*β��H�����	b�ڒ�XL��f\��OE�y�F�Z�ŷ?�?��7�9޽��1#Hxk�0��!筞�H
�Ꚋ�\��f���|66�������9��Z>/4�^A�Nؔ1���FVLIZ��ԨQ�AXG:#+I�x�DK古b���AC�a�Hm�`^T|uk��#�l^�ܥ�q�ԥk\�VAu��,���=/��� �ě�]R���q��L����\|Z�"i �� K�ÑEb��d��3�>�`M��x"?v�V�:�2�������ִ����R�zl�N��nh����c!i�ex��/��S�{#us��%9���������L@�[�F���Z�����{b���0g��a�J�'�x��İW�r�W�!��������Iƴp��t6z8�������s������3�?r;Sю.��%���%H���8�uh$q�c>xu��4,{[��s�ޘWS~����}ѫ������9�akC�#_O *�m��[}��uH�:�D(s9QZ�cQ��C�>x�~W���_8^�-�3p������z�I�PpP!9�b�������d�C��G���N߲'�q<�aH�7���C�)>��:���WI�[ݓ�>��[�$�ήٙ�tk�
��N�)�㎮a��sN��n7e��7�Lq/E~l�rE��XoW���<�z�nt�Q�="V��jnA�K����;D޵�CH���sߕd�8?+P'��pPb�b ��Vi���#���V�`���G�Ex�8�œ\���v�)L����5+Ջ�
	M:����B�y�׈0�q����wma�m3]�����\�{��<4�2������D*l��mp�� 7M*9�y�����2߻Zۿ�4d�|�a�(c�pn�5�_���� ���9���?Đ�[o������Ԇv}_��䢙nI�6��0 V����/a���̮���5�`��W����b�u��q6Gw��y���t>�fU�XNީ �8�u���C���*���YR������m�1��GӇ졮�D�"J��4���Y���'(�qr'v�۪��,t&�0�� ��mF+�6�3�R���G��w=uK��e�)��}lA��4m�`'�|T>Q��/�ѡ��CN�w��-V��\!LQ�����OE=l�64��X�axL���}�̑H�9�x:LЇ��Xfu�2u+[�'��ZKjz >��Y�(�%�����``E�\�y��p����\;}K4�M�p�E-�)���D2	:0:"e��F���B�;bc�XPժn>��3Q��^$�7���[�~F�C����j>A���v�����{�j2�o*���b�%`�
O��!��a6	�E�y ��.���}�U����e�-c:�-���ja�I��*bn����`k�#8m%"�p�脤�}}5�z3���?>�}�x�+ʔe!��%Vp�m�SL�5Y�ͭ5�L��{��ף��a�x�џ}R+���0wz�[�q�V�����d"̥`&�E5�y*�,�BM�J>9Q�O}����������0���� 8���v���O�����Vd�F�$�t�#z��I�nT���Ũ���b�2'�\��h�L�;�Xz}�qA#�V{[���`�@���͹鶙P�V��$9�����t�E��u� w�Cc(T$+�H�,��D��dW�=nv �.[�h,���E�Xô��e>�D@4�4U@u��ONQ>G�N��'�2R~Ӹ��pW�6�^����n`͘�@fV>{BT9�j��@���:x�Vʊ��Sb�Dt�i�j����6劏�1b?�P���;=��G�"d6sp�Y��V:F!�>�MN�bz�6F�`!������;�|ɖ��,�`h���?(��N;S�G�uC+�G��H 8�!Ti8�2�Vf�2�)uz-zi�&w���m+F�-�֦�Lf���9A�q ���A����4��e��T.�t��~���+��&=%h_LEq�Sse�{�$�S�M�l��O<㴒�P)�;��h����fd�%2b �e�pP�cs�H����㍿!1R!t��������A�e�̅0�U�Q��x�i��
'ږ��nU)���K7�$�����O��1Vf�{u���M�(�{YAz[��~�(�ƅ��~A�����χ�j�5d$9Hu�oN�i���J�m{ƜK��(�i��~�O�� �>#S�7F�[�,�}ve�]�-h~������3��&�X�.�G|Pġ��Jm��/)�迾�T�g�	�;&��b�V{��Ws�&�����I0����p��yw�W����_���Ν�nj��L2se5�G���(����R'T�,��=B^·/Ve��di&��z�����9�IH2a��pBl}4l�/��̾���h�z�ԧ#x?�)�^a����LWó&9U���j4���,F�*f��<.8�> X���k�<��cЫ�^��ޠ%�'��4M:�_$)�j�̱��$TWU�����Nz�{�3h�&fje��_�I��md�$��W�y�����+��>�i�dr�^L��f�����!4�&�۔�gd�!K���������'�R�)���%C����c`�'��}�-`/1�4����a��] �m{4�v#4�.^Ü���͢
���
��<��)n�s�P����b��I�Aldt�v렠H	n^���p1e���)Q�n��5��%B����2%S��P��	�¬Z�����Eܿ��-�k�6�s|�n�[3L$���7�D�MZ����O��Jd�{__��%������s� �hX��aD��;�8G��+��	�Iiú�4Y��,��+���@Sf��9r�a- �Vk��_�0[�/��(�����	�'W=c^�"a����/N�3I-�JnU1-1�$a�q��z���#��G�\ֆ>��&�a�(����V��~h��]R
�P��A5��BpҶWn�0�xǇ��Q��3����W������$��JrUf� ��m�<�;��2�p��jʽ�љR�pHo!vR���h�q���$K���z����)Ҫp7��qs��,̢�e&�Z���;�j��}�m�sߜ �J�	ә�p���T�8 ��{�:�!�w!�Y�����c@�rF�e4��0zDPˇ�-wC���
��\X�ءq����U"��9�6V��gQҜ��k�W�F�*�#E*B�
H�+ %%�ȸU�q2q�����д�ܟp������]?����L������WM����s_�^���ܨSHr �(�4F�Q�`�$�6�7��{�xb/]����^\�+�ÁB�$A0��~ʮΓhqg�����r�i|4�B3�^C��mJ�H�}uRI�zMb<�)��r�(����0 �o��F�Hŏ���!_�,�vߴIU$p�h\�ZĥvQv��&]0�*�f3�2�)*!��R`���3V���Tʢ*��pI�����Q.q�k�A`���מ���G#Y_�c���v��Xb��<"S//GɄ7�7$cb�(�ʣ5�|_��=�Il�1�2ndq���)��&�yV]���Ռ;n�Q���S�������\t/�.��D�r����pF�R~�G��B���a){��M?�t ����5l�E�_8"�K��5lg�$g�-K��q'��#ϼyu
#�y��Yz0�S>&�;�{(�ܽ]��������������z2t�}]Xc�__�ns���Ì���vSf���E�o�K�Z:e�
5��M���?<�2F:���Us���Xmy����U%�"oh��P�X������4GUg�l�8++r��-�@���HYN4�پ��\�W�x�C��dPj�eF���[<��Q)^A�?+�ɚn/Cٟw&ѭm�(Jǘ��-�d-�7/�B��A�$�Y�����2�+���zs��Є�Xvh+:��W[:R���T�-6��'c�;�n,d��_[�Y���#���~x�T��� ���AH����pN��H�GtS�y���Ƶ��m2��m��F.��h5�U ]u8K��v�%�dۀH�c�U��sP���mg���+_�4�: -6ݵy�m%?������)!LN�aկ�l�\	e���O��,gkAQX��Hw/����j�w�xh��3��x1� 1|��8��:O�0@���g�7\浟��t#�e��|Z�t�uU�euY���^(��CU�>6��D���ي;i��F[�l_}��ePE��*m�ޕ_���l�H����8��Xy�q|{I�Aw3�-͇��3ο����pQ�5i�1z:�Th2�!2��!D��5^Bj�I��Ho� �2�u閭#�+���	��e�B�g�0}���z]�N �Ʈͅ2��k�
��K�a�����;��<k�-�+�	�QO2�����p�7� �n�ow�]2ϯ{!������[j���v�����cD�kGN�/^�����U�}�7��̂��Մ�,u�;���t�Գ���N&���]��0���nğS��ƭ��^}ʙ�(I�����J�Z`4?��`h�9�����ذ*��nAn�0p�	����o��#>5dʎ>�����1.&�����D-�"�uB��G���E8�^W٣���o�K�,��G��wo�H�DC����k>�%��b�n�����D�
ɨ��TA���( 6�Ԩ���3WoMB�Se {��g���e��$4�kS`RK
�Cm�lY�]�G3Nk�Ԓ���3Q���(�Q�7"旦X�g�G���#� ؝M�r�,�L΂:�0)��93�dOg�.F��+m���B�7���|0ݜel}�H�h����ׂ՞��x���/`lq�̉O�2�Վx�d��s���בL�ͻ���wR�zjkcdT���HI}��lo/�	�H�?�z5�q&��H�-�$�$�Í~k˄�r4��Z��\%�������[>�t��O{��� s�5t�$��2�F-��� s��N+S�i$G��ۀ ޽�.�·N�����zN	�5c�lq#8�����OM��\��X�S�|�.w�M"�a��qz �1~-��VԔ�+��wcy�ӕ�T�:J��@a9`�� b)P9e�i8z��Տ}g�E�)��䫺�c2YbH"I���y'+�� �ž��[�X����e���{�����e������s��I���K���	�P�%c�� �G��<({�½O��JF�3��d|O����X�d鼶�#��?Tb0E��w�>�DhM�� �[�C���dŶ(�1-�¤�ј0e�|ț\a�m����_��H��=�g��2wN��>�z�)�����Xci.G�G�9b�Y����a��ξ4rA�f��e��UƘ>�f��z� �f�:Y��`�֥w�aY���dǼa��VCݍZ����(�0oQ,Ǚ�U?��wu�[F^K�YE�G:�pn*Qmt��\������,���Z���КL���
T*9g�E*�赥@�y=T2_�����0��[;<����&&��[��8j5��,����@S�s]�ڒX� 9�=b�~v�8������1,O`�r)�G�f�h{\A���?&����=��^�?m���D�5v��%����;ڂ��g=K���c��iњଣ\��&��5��l�(/w"����k�j�$0��Jj4Qp��e���V�D��/֟��~��G��)�R�*>|��ҩvg  ���~Q5�ֵ31���*Z�\f]���{ ��JS�sE���)e�Ő��
w�����O��bF8���Pn1#tOi��T�� �#���aZ��g1:?�/&�$���~M��S��R���$|���
����5D)���R���������X�&��X��K�f�+�,oy3��(�!j<��0j��?Vv������-u��۫*�6֟��V` i��E��	:ri��_GLr�5GJ O}�:bc�Ї�%�!�~�D��満促�,G�w�"�_&#v^�8k$�9:ǁ�:�}3�����'�r�Oi������#���T�'��5)MN���)p���nK���£���琔z����G��(�T�.��X���PJ��IL{}�vr����I#�ф@.�Iߔ�D5^A���ǘ�N�-_Pp�f25o�^
l�?��<h�.������R�M��y��k��݃�{�o��~$d�<G��\�ɉ!�7a�-�^�+������p��&������9��>��=#Cx�8q[��&��;3y�oa1C4��3�d����3M�L��!��5��)�<e���v�i��?�%��0�f��	���1T�նJ)W�
� ���ː�N������_��N2��HFP��<��S�>��I��-��9�QC5�����6|�	W�v�N�܏�lKM�u*�&-IG46^7W�l�0(�L]Bg�h���[��Z�
�NY��^y[C��&pߙ� S*��������	���.Kt^GhH�����f�o��L.O7�P���S���a��\4-uV�S3M�e�������ĭ�NL�!#K�5[��^��|�߀M�	*��!��y\,t@ӑ���2���T9��ҫ�E9��k����o�L��Ǔ���Ξ�&p}X���B����*��dؐ4���P�!Z����4�Y[1�!�1��T���I��c�A�� ��մ(�ˡ�Q�JH�6�mw��]�` =G�|����@`���p|%i�+�iy���E�d���YP�K�~�)ֺQ��O;���ޅK�r���,CDR �b�1 t^J$�>j
�M\x��H�'�����Vϵ �F�^֫8r��SK4�ɼ�շ|����g�0Q�J��a6B�de��Z	^�)NS��t�G#5v;M¶4���<���G����W?�F(���	l1�鎥5Z���I�TŚ�S�ȱ��<���l�o�t��8#�VE��:i���7}=!��F�+�R2!��a�\�n横֧�]����K��pr�m �tX��M,ɞN1h>)4�o,�B��������
��#,�}���>�tJ>�oS��(��{�����YP��)�.+�R_3Z}т���у<��I��P�h�؀E]���#f�!H�����g����}������/�)�1"#m'bL�%ZH�+��h(�z�����4)��L��[�H7	,	碻5����B���~{�C4��\�m//���|�B�
Ȕ�:��.qg�mKKc��`9ƒt	�79�T<f�H�g;��O!� �3�4;L��h�r(Y�؏�B�b��S�K��k%oo�����w.!}oΡ=�c��g���Z�\�-{n�k�不�mS7�A�X~����>����7�Հ�%�=��K0U��m(�w��������l�Vȹ���_�IX���߄)�KԀ� �����y,̭x�(���Ng�pZ�ַ�y]��]���eɀ[q�`8�%Y3�zlgq�=�V��umB*�� nq���b�`"�1Ľ��]ym�
���8�%��C���c~J��)['�a<cm�Ģ��r���P�3�;u F�����߀�K������56���y;��omB�m�͡�>	_b�8Ec�4�_��Y�C�����<��� )WM��b!`�+#ai�H��1[��'ݙÞ�b8f���Z�w��B2�o�u׻�vN�����#(�e�Q��8D�>�3�"��a׃�[�|�R/"���瑑e���O=��|^x��	Ź�n���ס�����+�K�R�uMIʩ�*f�yP�������s��)�+�m�"�r��;!���L2�:��A_L�i�J?�ӧt&����;[U|Y��d�����=^�㌳���
ۢg�%	�ݰO�Q�е	҇`yS1e�(M�7���`W�Y*��hO��|���\��Bw���b�j�Ƅ�-ת�����k��Sݖ&����#�Ud����^$j�<�M�fH.H�v����{���'�@���۷�*z�KQ��%Z8g���4r��V�1���
-Z'h�Ech�ӂ�ND�����ޣ���R�pq�	[(R����_�e�-H�_�+qf�OO�2J(�[ek�ZI��0�뉴8ʀ���5�P�Pw�=�v�D$�Nax��x�W#q?.�vu�V*�d�g3p�l�C�.L�+۵��/R� �ǆ�	����u�A��g"����ˆ4�EB7���rj]��{���5���F���k�?�/��!G�8���C$C�F��L�Kk89�L;�D����oZ��,4/k/Ə��4�s¥B]���h�MHo���F#m�g�;wl��Ax�/���������ű����X�T*�$>q�i����in���]�����H�'��$7.��'��v��r��s�.׻�{�cOW��RG�e�\��o��-���(�Y���wW�0P��C5���	��ůԪdhl"\���\B��Զ2��^(�ÿdC���|%�w0`q�����&` �e���zf�B���(O�&���;��^�AR7�"i�+�Z�-�qM ϸ+5И
��sWt����7����ߙp�2g�⎧�O=�b����i�pņ�7�����ɔt7^0.%S���{.�~�Չ1�JdY�r��y��V:�r���G9�z�:Q;�*�5Mw�
K��q��r+��h����^���v�twWR���"y����s���{�$y^����ps��4n��"1}�y�.t��7��_S:j�?X��j	Ty$�%��q��H#b���|N��x]��å�8�S�U��K~��[CW����t�}��-�~�dh�YoN��3�����X=�TأZ>F|)�us�I���%��fiPQ6��"�:C{&�Wl��{� ]������ج��j��Ztô�\���7O�3H!�0���2)S�+��	��]�|�;���y��u���O���ԟ��$#�w�S�=�����Ƽ5���OI���ݯތ`6,c�f`�yCD�_iN���5�N+R�c*�;����q�[�A�,��!ҭ�<b���8������v��c�2p��󛤓�>��%,����E�C�8kcZZ�f�zoY��ӧP���Υq�c$�nb#�1���X�����s<���� ��,�7�d`��/Aޒ����d�b�V�l�vA�lqe���J�ێ�Lө�P�Jk/3bJ��"w�R�y�w���8Ϡ'�	��$'����=6�H!��d�ܖ�%�'=�)���YK�C{���~qN�.Vl���D$��ã�o�)��x�.ǥ�\�螿�I�Pn��p���i��j�M��*�����7���{���zKVP!�8HY��{�d)ށ��\J��4N:�Qy���m���-b�}ץ��?t�cf��*:L��n]/����Y(�ox�
|�/T)�]A�U��ms �9A}����_�IF��4աq @~� l�a�����%�ގl����q*�?�,���Y(8�[��,�	^܀Ծo�l\i��s~�M4�$����C�r;9"6��&VH�;��O�Nif�UȦ��ޥ�[9Df%I�"�u���u�k�����q�5�M+�9c͞.(�X(!�e]�V��e�O�Y_︕0�����9�M+�
O�Nl z=�T��NMIQ�(������ݾ�
==2�O�|lU9�m�쌴�'>y�Q�,#8����P�� Iv�(��q�;M�")�@�E����� ���~�I��@���*�j�8{)&9h+^TE��=bܥ��C��T��
���R.�u�8���ZhR{�>��x�}7-;yn����p���B���=�����ɋ�`p���2S���LH����4�Ռ��l,U`\�9��@�]�G�'���'T�.��8К��3D駂�i�=Il2~�v�DK	��c���,wK�|�s�a6)}�����K�����#8@�L-)��&�f�1ň��]@LJXF���:P�����7}�+}��`ٴ� �Ҿ�Yǂ�y9�9AH7M������/U�A�@k�<�֞��葦�MY��w��/X�]0	c Ď[�_&���LλF&t�w�G�]��ZZDfi4�5��۲$��'r:�GGK�X�dM����V�/2\��d����<���'d�����̥}�0������X�9m$x5���ٸ�jjq	%h�ӿ��X�\�S�Ќ����c<P'�v���k�tq�����o�(Z���wo�����010mfi��� �,���[��~n�~��t��8l�9i��ě�T�ʩ�9
�PERW��Z޲F�	��z9:�@�2r�ؽ��ކ��ƕO���ړ�����D
4I59�ǁ� �.FVq�a7I�u�����p�8��f���}�ʿ������|=����8���ć����s�gX0�bǩ�K,�(]�L0�u�)�~��P����*�Kp.����%UD��(��$|pZ7+�H�
/⋫o�R�w��)�~��*�Ov��0}}��,��
�P��=�-K Fy4]MiM��~7�"��D�e����_��; ��ӵ-�!��&`�<u-׹?m�OB���ݑ0d�F5]�w���׏23�X�Lx�MY9T��Q�|r�I��#X�3�*�y>��}}P�f�f�����;O[����p�y�;�ޖ/����e!��U-���k`V���p�Y+Db�t��\������m�|��֧C0�\Y*��"�S�(��
�Xe��o�a9D��5ֵ5��x{e���� ߡ)s@�x~�G��N��"�ͻOOZ7��B���O 8=p˛_��\kE6�d(MJ;Jc���� ��n�J̩Ϳ��r�s���Fgԏ:79+	�2�0�6���>�5nt�ϣ�R��\�Z�<��8�Yh�cNG���W-�����|]�1R���<h�KI�fJ+S^�y��X�R�� 3�Ĕ��K} �9�wQ��?�!О��~x�vw��jJ���y�� )e�_�v�3��'�,����U�"��n���a�LWUƜ�	'~u�<�	���ni<9m�l� ��[!���Tm��
�-��[�?�5�)��q�*�]R}V*�s��O���$�rV�]XJ��X���V�Wϸ; �o�c������SuD@nsϪ:$�Z�˽�W��ƃ����&���`��xf6���L�8-���a��ԭu*���/����B��'<�lo��|�	���G(�(X}�����wO��Á�g���Lm��PmR��s@������^"<����v�1�2Z��Q�gӗ1$����u���h�I��r������e���8�\� A�����z�'؅D���s�&]������MP|)�������
����&�����B��>�b���x�� kC�u'E)��ιJM�4
�scY�M��[(�<бm�"�L��UDcF�)��pkۯ�n�ͻ������#]��n�GB��ې�+�����<�]4�0i']}�'5�.!�Ԍ��D���Ѫ�-I٘�y��\�B�4��,K,�V4��S���Keʀ���˧5��^7���Y�CyM�����g�~��T�Հ���,��G��i����?�v{5�7�Mu�/�Z�dy������DFɸ�Tz)0pj�#������G16N��}�۸����q�r�Ő�v��x�%�N+���?)�%�^ah�RD,�@M�$2]R;�/��3q���NG)X��}8�u��0\e�E>;Qg񱋨����[��-@��: ��@�*A�C�l�LU��-[{a��r�Iڐ�'�8FS�%��k �%��w�}q�-Cj�6�`���&��V]�-Rލ��۵WS���1�����=0��B���C�w'#&��kcNj��4�H�3
�6D�YW�jW�7����V��q�L��yq1Ϛ�-r<ɳ���s��׾˳��L ��W���_��@��0�~A-j~X��(�N]Ed8��uAy�ȭ�5
a�,���F����
���|M�v��O����[7YV�Q��@LAO�B�
���lw�i�ՏP�Eg�A�>,B�(X��*6���u6��^�=��}K���2<�rxk�7-˸?{�����}��8������W�C��ÞEܮ�9,�_����6��3Wg�X�3=���3�_8&hQT<��2V��i�Pܖ�7��� jϗ<��ʦEEj=萒HNIf�I7��၈��=��K��y�K!O����G�!Ο@�*ECb�5@�̛��ͅEbڣ���)2?g�	 \�mYUVk�kc�ٽ܆&�[�[�GM-�q�jT*3����h���7�+s>�*Q�t�����زnO���%�<����$h�V�r)(�Q��q��҇Ώ�����	%��C`�]�(�3�� ci���� _R/o��8�x�v���)���P�������ֳ��վ6{��(��c��~�@�?�� :ld��ֲ_N`���c8�-29f�bi�0�mM.���m\i-_�Q����s1�N�pr�c�02�D8�>L��8�NLU����܀NN���@#��;>�K�88���d�
��l0^Q�	�����&Bk!Y�B�e�3�Lp����Wo�c�n�9&�Ԝ�Gm��W20W2G�σ'�DY�6�"�9���.=]����kR+�݆��?E�3o�B�t�9z>�"b�x��F�r��nZ H���ѱ_b2{�x�	�I���˶˧�;���5������+f��`O�.qx���Q�Yb��+�߹�q�����6�d�3P���L��b����P��as�#0���e7⤏$����b-+��',��.+|w��2��8,)s?��(�^ap�.Tۖ)i^�+%��}S;50st��V%�F��h�OO6&����x�Qb��c��Q��4Pi��2W_�7��*��)u��kuӱ��	\���
s�iؠ���>P��ѯ���i�;�s~�p��B�,�F���������C�5��O��M��ԅQj�~�`t�9$���g	�ZL����5�|��IpE#��X@����X��s_���h���{�V�fm���̟��P|&\��x�}�V��bX��
�����EW 
#���٪�Yn�Ӧ�<x��8O���Gm��q��;�UNgx(ݒ����7��0���a'��׺����m:�ZF�;�\��n<�s������ꄼ��c�g�c�z3U	K���lıo,W#�j�ƳA�r�D� R�HQ�;���j�;
�1���$d�壢�#��Uע�?�/���c���M�%3��VbX�E����G���`��UK��0����o J����:��X2�t��Q��Md��� B&����l'��Td������V+���d�K�5���/��F ��Y2.�w����cY)�샽8&��9�n�v|	�V?&�fM�F'JT�]��Ii����>PƱ��s��̌)'^��g�H��j>� Gzr1�Y,��va�|b� �"o�_�Ϻ]=^��$���>��\���*ř�}u	Խ��|	~}ƹp�pR�7��B���;�E��-� �[��C��{���� I��q��VU�Z���-���_�,_��d}����K�Qۺh�)�� b�Mp��X���\+%	q�/g~�|N�U�*n�;���
�]�Q��3�k��,�y��,N�w�F/�yxR`c3������x���+�~
�{�r�@��D�oHWA�����v��[V
�����/�8��J�8�����|o��=��1\�d�i�J�H���!�x�z9���Vk%/�4}�;��Ja�$�[�5�B'(�C��q���%�JO'�&%���4���3�%ޤ��*y�d�n�#� ���v��u����P��I.� �E��Ⱥo������L��J�P�'"�����#�5�H�d[>�
5>��i���RhR����e|��l�l�2��
�)�3n�mK���	d��.0؛�+��#��b/H";��C��&�I�ʵ}�5���xTXl�� LTf��v�p�Ћ��o{���%I��j��n?���ÿ��͋ ��|&H,����ŞNz���oߨ��i����7��NH�R�j�v8!��\��3fN5A�%q��g���&��Ţ�	{� w
�4�D�Ms|=��G�I����z� ж5�<<�"��I�\�*x�yC�w�H��)uIq����ՁQ�xHY��=/�_�!���y�-�T	F��'�1\��s���c7r`Q���oXD�Yؙ�[��L� ��\�
[s aƼ8P_i�iq�R�υ�^�%�(��v�2����­#�20ޢhJE��\�n�RU���V�I���U�U����LJ����D�`e�S
#���HQ;%�1���^I�_���9�M�u�Ds�M�����^E��<tҊV�V�ÕS|��Pg\��T<UVD��L��=��t%���1���4��U���)��;�j��kq�%I����4��7�]��|'�9R/�L(X�#c3Q��H�;o���׀�������2���<*�z��BH��|N�ZpGD!�`��"�X�&���/c���w==��ɉ���\%��c�W�l�k�.�An
�&.�K���yp�cj]h3����Y�߬H�!S����Cw�_p��c�T�/��p�H^�3��Nc=�����~U�Γ$A�Pa��}(��!��<��,Ux�-�`���)�����>N/�
��d�5�Δn,H��	�c���j(Q��Q*f��H��Q{��z|�C>�%��{�m��]����)}�!��Os7�ᓇ&	^Tٙ�{ͽUh�E��o�ڀ�fvef�5*S\fB��]���1�6�3�S���g�'�������&�����AP��W�D�	� �#�?x�B3�ZҲ�������S�+5r��5�^���S�Z8���R�_��	њ��
i9�#���{r0�$r�v���� ^`��.�	)ä���v���ыCda�!pw˕=+�[A�F�0\���K��#hI�(�=D�ݸ����<�h*�W���-�=nJ��`�@A8��*gJ��8��'�v�ؒ�����@��Q��eƬk)�2sIi�T�6� ���̣��߱������h��,Vi��YO�i��I�=��e�M@�T)r7�Met�oå�v����h�����Uvв
�z�$��j^[����I�R���@����ԋ�����­�+�y�`�/�^�0�uߝ]��% �P$M�bDT��!���G�m*s��93�I��/F�4�NH]L#�A+}�Ł����OCž?�T�]�<�G�̾�r�.H/s)��%�]��yܰ]Sw��]��0¢�'ԷE$?1����wT�ևp��n��\�) ��	��߫�1���B�%9�m�aGG�^,���x�EH�5[>j0���r��6�Z��R�p�W�Jm���5��LuWP���@���@��Ԍ�J!�.�����9%�>[<���ûa�HQ���8%�5�������D�� �Ѝ(�q>a��'ɣfX<kA0��X��̛<.�����MpZ}G�+�[��&���[��w�=!����w��Q�J���iܺ����;�,���Z.����>��]��\���ite'�/Y��&�bD��j'=f���� ԚU9ˆ`�i���^䑰k���`���u���vm�+(��p�Y;;TB[��gp�f�n��������~7Υ�\�VkrB�c�}�|��d��}%�����/(҂�*��	�}����	�5RxP�v�jM�nwt���R��C�����͈K���5U���2��x���]&/&N^��@`����(*kKK9���>1�XS���}l���~%��Y��ϱ����x/k3��t���]8(I�(�;�|��;4.�D�!��-���q�\��5ٲ�z,�>�h�R���J
�wSu�2Z�m�����j�@��p�?D���;�ڐ�����}�w'U�=/�f�j�{��ʋ�{���?b��b��Nm����ue!�5��a�d���F�ُ�����,�_m�AkQ��t�-��[~�E<� :^�!�sX������X3m�6������5 �d��IZ¨K�Y����	��5������Dx�b�J��ioC������,�ƚX'�'i�?��
����~�K��5���x�m��"�����8�矴��j�h֎�MVg��t&�J"���ϔ����N��R���ҥQH,]�8����F��g�O�V���3��bG�y�$!^���"��"�&_v1_Bw!�s)�nRP��i�4��+�OAM��t��$�~��b.�?R��Y�qn!��Zs����F����^�Ѝ~p���Zv��w�����DI�d�C|ڴ�����Ԅ��z<
xE�����x�˃��P�E���\K���Z3��yfwҗB~�:��:	:�.=3�Kp���-�_(���z����NQ���c���Q�.��k�\��W7�o7ױ)�P��yo͌�7[�6>/��i�]	�&��.�WRҗ��>�p�=b܈��[���"Q�y�Le�}R�Ꝋ��t�c�w����iyE���k#4r=pޡ�t�I#�����a�z|1l?�H��' 4pcD�����@4��*g����h�3��s�w�'�Kl����/�k��*�ex��2y����P�����\�\�w>W��ܜ��	&uP�� E�?ܙ�������/�F9���Ɇ��&��J0nu-a�15�H����w�y��q�t��x�>%�(��u�O
S�oȟnݾ�4���"��c���8itAG��L�r"'���Ȱ�GK�L��ٙ���> ���?�臑Rw�����=����
���J�h	�VF@�؛ZWķ ���2Y0�ɠ?Ѿ�JJa��P���X[�mf�Z�ï�':�>��r���__���3_ů�a0zi%}s�󡀫dAIK[�0��u�=l	�p���4zfy� Sst,*a��nb�jx��
�Ug{�r�F�����B~S��}0�.�tQ�ˌ9G] ��O�R����F���b�D��9����q7K$�mh|� ��5��a!�Y����t��7CC�D,�|v�j5	�(��o3��������"P$��x9�~��滵�|x$��ϋZ#�[�:UY�dA��0҉�Ռ��������������7d�`��y������fG����Dps�/�`������u�'w�m����%���]G7�ӂJ�f>"|I�U��gj[&�U/Ъ��	m~$ٵ�y�QI�wwa%<��˃X��'tr��_��ܴ�cL���W&�go�}��B��?TO�&�֭�`�%qK�mv.����>��V;P�(Q�SU����%{sHB��e1��}�>���'С�x��N�)5/�ˬtr���E%��PۂР�u�$����̅ó��mG:CL�sL@_#_o�"T"��ehR��2|��|��f���hw(`װ?u�8�AV8]�M���y�!!�Ir�8�)�}#�
Zg���/��x9�n��j�7c�>l���@J�+�i������ɔN�U0Up��i���ߴ\���a�K-�wN�M}2�-Ĝ���P�8X
�rl��� �y�c�����]ZX梇R_X��f0�5H�ű����NE2����q���Ӣs�,�z&�b�B9^E��/*vY�Z��<f�L;t��6�X��~�����ćL�{vཷd%OL=�29�u�4��!P��~��6�"�u���禁 �K�B�'J���_F	��1?��K�νΖ|�L�"~�	��4,��' �3(MRj_L������CG��	H�	_L�yW���Zۜ�]ߔ��C��zG/�&a�K���(�!ه6�/Uͩ��Ͽ.�P���&8���ϝ
��f��{x�{!��Ee?�g��xw^��]"���>!C����LoI(�x���)�-��ȧ<c�=�q�t�C��℘@��&t��_f���<Ed���3��ދL��tv����不�L�f�1����y)Q�FB%�`�W�'�Y��ǥ���<J-d5`�P� 3n�.c��Ya񘃈�"�rIh%��<�Oqx��F�����1qfB�n0��2}ee:<,G��7��J�1�Y8�CÀ��vH\���r�M�f��v�op�h�� ���e��,%��p����w�[����//U���>E%�M�����RG��g��6n�������
�s��$�d����]�o�{�w�3r+M 4��+e�M%
���|�Y�˦�����V1����������DK�����b���2�;tz$ц��l囉�bp=��V��w���tD�.u��"��l��e�� ݹK�-��)~��J���z�a�ث�"�T�-��6���Y-�lh3MtpoQ}��E��l��pv*\g�@�F��"�#���_|=A����+�%t<Wm�璴�2�uHt���0��Q���)6�S<�z��|�\(YR��/e�I !7���1R�ʷ*t�t�mZ��p�V\&�wa��@�%�٘Z�ۗonXӽ���BS��M������B��&�Az�c��9���sas'�Q��o�P�aY�AF�m��ܭ��.��
+����*��ګ��}�ئ��ȏ��n���Y��h`�d���i�������x�6�
X&���jJaW��iͬ�F�ӏ�+b��J���D��^��N�
����V(e��=�+#������d��TBp�q���(5
+,ɓ��=�%�l2�-�1<��Qi��^�W���RU�׋N4,$g��?�����س��bG@u�Ax��?�ͲT]��C��I{9ɨ�/D�Jx�g�i'����yϪ��4����M�x� �Xkwo{$�fa���ĭ�Ha�!�&�
V_x-ӈ�?���8��s58n��_{O�P^j�S5T�����0�HW���[��4�����|��z�FK���D;{1�	j�:�W��w��i�5J��R&����|_��y���Q�Q�
�\2r�!ӟD�%��]��_x�c0�-�Rе�)�9\?ԁ�r�?�j1wq�W�F#�Qh��ʯP#��]=ΡMD��l�Z ���Σ�ʉك�i/}x�����V�#K��k����UJ~�����"0�Dc}���Q&����n�W�|p��;1����+U��®���W���i�a6Ž6pv�Ѹ�✖o�2���ȴ��S�����-�'BA����v�`r�޺0�'�RI9�PK^���nLK����pG	$�Z��V�_��:.bS���= ǩ�*R�D��aNt!f�[���+	QV�mA%p"j�6��W]`�hC��j����e��d���<� � ��߯5���N���ڕ��Y����m�?�@?�Y#��?�ks��/���Z�D�Ԋ��KC��p�c�?RB�?��.>�Qo��9i
�M�U��b�	
i�#�"�U�!�l���B_6.5��Ұ*����O����+�ƧuU�!�}�5��i�D��
.Q�9�E�9/�2������ƛ-�'f�vd����c��؆;@DBOt���tA2>~H�G�M
�u5g��p^�2���z���2� 3>�V���]�J-��3B#NF?����c5��B߂0�o���<�>m�AM�0 ����uyy+�mV"��PؔO���8�
 ���WnB5���wNC�~pV2�?��tI.y���e�x�ai(~o�꒫�t�3���Q��e5�՗DOɖ�|�Y�u\�����oj�~�?l�`�^L��G���j��ߝ�	LV؝�F�k�G3�"���G􋱳+o59������R��,'�h��'�����-ble#A�5�kv��[[_T��ȓ���c�V],���-�;
��M)��O�x� �.��@5��ʠ�J�CL̏?��niӇty����Y�i ��*��ʢ���U
V@��W��G��fROd~V'�*�� �f� ��?H�P/^;g$0����K��fx�lq��[���1�^�CU�	x\�4a��r �箜�.��y�Q6XF��F�$�m�#3(����i��0>�\f�t��hӂ&h��F�Qd�����s'N�G�����v9R���F �\I��{�0+�d��%�)���O[�r6�xc�#�#	J���pΣS�x;i�|iZ���A¢��^�6�!�qÆ�񮮈�^�������.ղc���x׸Wc�F�<I����
骴�,*OE��g/:��d��=��ŝL��R���8�{�5iG�¸5�	g&a���F�y�f|4�Z[�}�s�hx,���M�4泼��:/��LN�U�ΘF�� ް��'��X��@#+� ��wpK,nƽ������@��(�i4���cv/���������O-<SO$k+9���Ze�gv�5{�N˗D�;��p�?9�z�SY���P!��Nꔶ��{�r,����NT_&�j�f���u�'W�:1��}@zI���Z�(�z�&c�I�{5�=ވf/Q���m��r'�v�=��e��t��*{K)�"�|�@�)4m	��
ĉs����+P~�[�P��JO���aU��X��!�+���|��\��Y+Q��$�@tt��y�J��79Vc}#��p�����;�uڸ0)��x�{������:B���c+�_����q]���|o�71��Rk;t �e~��Aރ��8�IRgI����Bi��P'.N����qG��Yq����[��[����"�f�IK���\�!��̆d����:�*�����4��sM��ZS�R������E��ukANV7S�1�$�U�Q�M��2����T��5�%H:#��P����X}��}��_�c�_F����UQ@��O���4�I�
O[?��5�d�m���l�V�y�ל���0�:Ȣ�C\�*��,8X$�֪c`��et�j���L;y&	��� ��G!�|f�G��[m�f�����B2�<n���i'����h��Q��2��\���p^��¯g�ڨ�l����K�;�A��t�F�Q�"h$Y)�o6Pc>���1�y1�Ȉ�Oxޣ�7)n�|�[l�GS�2��oD||�]��ߍ���J�4�YI&��$\��}��
{��,�.�.Pk��U�k�;Ûᇔy�?��X�(X�3�7�Oy�je�S��$f���,)�}vȢwQ�-YB"Y��������:'���'�G��;ީ��R%B�irA,S�/�Q.�P�I�S�D�r>�ߌ/ߞ��^�f69[%$���6/W#g�#��ӡ>ϙ�KO����������7U�5KǍ9[�Z����@>b[��ɩU��1�З�rE�V�x�vM��d�1�' �h�{L[���kgbQř�|�MD��	-��E��)�LxH�/5e���_��� ���Z>B��e	�;���|�ӝ����"V�%�f����պD��2}n�O8�����v_����+�d!���ʢ ��Y�Հ�00d����I�<�,Qt��t�":��R��U��|1i��O��ZEL�&��s���H��M�h����b�����v�|����K}����`2�N_Y�����Dm��A첝d?�5�3��RjL�}�8�Ճ��:G�����X'�T�$u+�$$�k@���ޠ��o��อ���>��שr�� ��^0�;�c0�����.�\�y	�w�췎G�`P�P׺R𵳖��{%!�Num۸�KnK�[A��2����s� �f3�ov�4����T�]�{#vz��J)�`�b�LL��1/=�����{����iY��@!k��QF[�ML2]��׶��X�X��!ޟ���sc�7U,x�6);?��<8�B���h:%�_�)`gk	h���'�`�qK~+�if[��X�B�e5~i�f�"i�X�#�P߹w��TL3�m�<�2Q��{l;�!���~p,�^��Hj�j���U_?� �p�wi"8"]�=���s�I�Im�!����f�bLՓvcssuY�Mg�8R�k�ĕ`���b&�{��u�R�ƍ�;+� �R�_��ңг�k��G�/����f�D��r�]�ő�E+�-H�xep�]�� �Ƀ�GO߇��d��֫P|���)ƛ]��Hл�����b޴�(�y.[a�l����g,���i+W�Ɋ�$7�5<DTg�T/�'<��{��*5HJ�ɟ��$��E�Cy} �x�=܅��܄�����27Wk�dk�6r�m7��9�K�PH;ȝV)@��\2)-͏�'�w�?m$[���YF�ڮ�UO����n�����r�Nv���Τ���GAi6��\˓W��n5��`$���̞�)x?g��'�%:e���y�� ��Ɓ+KxiR��{�Mv��K��g���4��`���8���'9�*D)��	|U�a9�]�QG�kr��)㈭eF��~FfAs	�����>�
+Z�)���,kc@�Z�x.3�ҝN�dv؟]e�x�0P%����m͗�|#��3�S�L�2[�����x�-_f�񊭤q	`�����y]Ki�^\�c3`�X_F�x�����^s#�}�q�̡�;`i��
�K.n��^�H﮵H��:��_�t�%���w=Bq֊�b�����VNx��@,��{R���?Wyc��Ekm �d�p��Ju��]��Tڄy�ЌCM��Y[�<�$k-�5թ5�K�.7�?*��ij��V����V��%�����|_� z%�Y������1����w!�0�Ob��N�\�%�"�;��+�1La0?_���G��i㈬�/R�}�z�z>��	�Tv��`x�v�e^x�� ��qE2\J�W�v���F� �[��@A��$��pb=������Z2lz���O�U%���	nMDr��g����d�M
z����T09��~��ci�Y�>��i�2V)��M�33m��D[^�Ǧ"���*-g�S|�H��1��)�7�J[Sn��}���a���'6��V���&?E3�6�Qwb鷦����
y%�O�z�e��.�N�vC`�LG�W����1Yqܗ]�%$LHo�������BS;A����{�C�q�FO���{�|_y=F�ג	u(-x��8dD��0P�����$��FL�
�-Ds��i!����kG
�#��0h�8;'w�m�+}^n�5� ��"1���a�T���L_%F�,mN�U���!\-� �`#����J�K�jr����L�v�Lk^'�KGC����H��7J���&׼����9�����K��_���-�$�g"�dg%�15:������6<�]�A�{4 X�Ǆ��
h�w�����9+4����M���xPNH��� ��(���_q�[-�5�{R�/N@t�h:�R[����}�wd[P�m	S�F����k�Lxm�-Q��,�b)ᇐ�MpI������ŵ?^�@��Ù�ŋ��[`C���_���s�^�M9|�<�Fl���Z��l��og�t�і����w����ni�q��b:��7H��p�����-̢�޴�?������	�_�X::3�A�vK�_���Ҙ=�h�!(I���x�ŕ8Vx�|! w�ɭ֜r]����D!H�ߌ�>����s�]�f������9g��}$o�c��i�hL�����yr�)�*;l
K��ͥ�nx���C喉1z��3�����jo���F�<k�YZT��9��(-�S��}�n�0��:V�tJ�A{�A����=�
��z&�%�����f��Ͳ-�����1*қ^զ��_�Of{A�����ʼg �UC���/��Rc�V��)n"��˴[���5�ک�uj��>��y4)#�@+8�_q�t��$�[yGh^+��^�~;"��y�Ao��B�ry��K�~޻e�H2
����@j��:��8D�
�Ӗ��b��~F<�$z�|���|q�o�IXmL�B-��R�
�b;Q�r�%�}��6I����.FuQ�����p�� ?�; ���w=�.�ow�մO" �K$0����a��O2.R����yJ��;m����#C�=�
��k��e~�����e��]
��C؁�';Fl�#طb�u���|/�c��&=ٹ:�:<���V:+�o�L�8�/n�u��m }4*�u�	g���hi~�0�i����H"�Dk�>>��[9vg���"�:�y��'�k/�i.�\V4|?�S�b��L9�Bl���$��F�B�K����l��
����1��~c��r��D?f��q�e�It!m�P���W <J�ƹi�岱����HU���;k�(�c��h�"�jW�/Ջ��e׺e�4��,��C:%y�M=D�ܮ�L�Uj���-xh}42�c�+`�J���/��J)�e$ j�f��Qဨ<��=���0p806�Z�ɚ=�qXkk���['_�E��)%��&Y�&X@c�R,�O�i��R�p�W ed執�Pb������;J@����5�o�������	ٸ(�-,�I����?2���b��3�DSW�c�!Ph!$<1+3;yk���t��B�/����6��W�����cG]Hh~��5��� ���Tj[M��c�����&Ṇ458�-�A�eC�"�	��D	o��r�;R�ha��^W���71Ci���D�>Q� QՑ=x���i��g�׌�%��gH[�_
��bL@޴Yk���
�q?S�̚�Y_��B�Pg���&֢)W{��H��b�N�O���0
�,�|"�OY3'�2�L�l�94�,�v��=k$-�*�����"�{h������������:����9���a��t8�����=� ��l�<e�t��8���C7��,!{Pa���aZ9�T��6�g�L��P����G���'�K,�w��c�:�C��<�RA)���5����`�:�g"�K���7�J�V�+�o��a����/J�e)����⿽�dU"�%7;�&�]�`C�:J����A��(��%*���Ϸ���͌���`��-\��j�l'J#����ڤ��c<6	���%�Dܤ���έ�*��
��kMD;d(a3Y�>����6���I)x�mA�-7�P%:�1��t�Z#���^s�!���1 ��C��'�!��L��G��������tc�AX������"у�A sp7�nS�؝7���f�+F)�`MC��bx�qgZ$��
DÓ+h�Et܌�uN�Jf�p�b��.��'�5�|Eۃz]y� �����������5y'm
��������[����7��d:r|M��T��&�0p��sM�yA�Ǝlo��mh�V�c�E@��zE�
vD*�����u��@�OV��H,n��]�]cj��sspl��;�_�p94��n�A,��s�����&(TTZ�j�4o	�b&�VT��~"��ѿ.z��@��� �O�M�tx|�o����5�$�A�[��\���}z)���2���}�<�;h�0�ST<rK�uV2]ADx(B�>���{�\�]�&��A��\����Z�h�-N�*I[���PgJ(���& gO�l7�3���q�bܮ��U 9��4Z�#g5��b���V�V~��s�����cT�:���EOH1����=5U�~���7((1��}	u�Ċ5�9.X$_��Ǚ�`�C���~j)�8: K0l��f�] \\)��!
8X��U,()���)�?��=Y��:2y�r���Z��=��g��f��U����	v)�bv	�!����[*a���������}6g�+���`��.ګ��aVPc���?Ӹ]	��G)])����+�ò<שr��$�T�EE�W3��ڔ;�,g��>^�2@T���
��F�,Jp֔�SwR�ĝ����FY�'$�|yf�yD��o��j;L�c�4�� �}���&e#YX1�S���p�u�=s$>���᡻�����ҵu�ڍ��/�n��̼@Y�.u�����L}w?��i�Z��9m���O�8� ��n�&w��Eo�����>BJf�ۭ\(��4�RY�ZM�-�/n0���iri�M\����opm�+A�*�kvаǟ�Vv�$\�;y	�A_ج,_��]TiI|%_,Ц�v�Z	P�B�h��]�i�+14'u67X��$�a"�v�'���s��Ruf�6�������(�;)^+�p�)�eUqճ�P�J���)kù+���_Ts�['`�?��ӑ��9����4SHEz�!}*!P���8V'N�?q"2�����`6"�{���(�%�,}�P�f�Uc�^��0�v�u�/��v�����0ȃ���Yw���.A��1M�!D�TV�=�Uh\U	�lޓ�WAUa�+1�83<�f)L���/R���TY�H���zi�<�J�Vj�P	���K\����Ó��O����B �>z���܀/{|}�z��}8$�����ٷ���h���ƇZ5���38�R���?�ʿd������Sq{����:���|*�z%�����Þ���0��AAa�E� �ֆ5���ȉ>=^�t�p@EK��)|��6��=(8�Ff|
r�}ͽ�~�#-X����c����Mz	����8y�*!��wD��	?]4���l���䌨UN��B��?�bc����Jxԧ2�JLa`�ټ�.�6D��} |�`76�<�?�6qP�A��E%(�@�>�Q���a:̩?�7)�_Ju�cO���00��f���Ӌ�Ԅ�q#]s���<tb&��v�6;�å��p�Ln��=�l��&$���>���8s��S�K�.�X�I�E<�&LT�3�������⸿�b�ˢխ���m����+����C�-��r4W�%��R���<��Ӭߠȯ���m5I�?�c8�Fl00�lE���ǜ���E��!�f|����ݞK����(�iJ.=\I��yQ�J�J���ٌzM��
I����LF>��o���!��0,H�f�>B�7��{yNŧ�_����D�@Q���T6�zhC-''���[��f.!ߓ��!J�C>��sN���8��S��I.�����έ�C��@���Y�H�x���$RC��+�kp��x�n��llVľ?������ O^�*P��Q� }��B(��&!M�{s'?�>j�k�(zXR	����9�����	N�SL��.�>_]������]��<��#1�Ӓx��Y����5g�KU�"*���*Q$om�'<�Μ�}�O��Ze������*x�Fn̳D��
�q1
���t�=᷁���<�J+�.�+B1';��$��b ��_&�GO)iM��v>J|f��{�_HqGc��h�Ȅ�+��N�Y6����#t��G�\�}�?SMPs�Lp�{��;�Z��.����O\�1#�'I��~|�>k�f�+��J0�P/�̭��;S�HL���� ��d��ӿz�ܔ?�/��7���1�=[��^��R\�v����"����8k�x�42�}�G�jĶ���l��h��M3�{�w�-#=�:�0���/M&�Ĳ�x�/��b����Nk��~'Jn�����e4-��I��j��]�.TP�1���w���	w����@�|K�(f�t,U�����gr.��S�1�_��xH���+����+�3�&��r="p��R �D� ��\����Q�q�s��������6��	�_��>ݍ ��d��ύqs�gI��x'@}
O��5�gZJN+Ӈ�������{����1���G���/�`Ǆ�֥�N��jƔn� w�z��=�r�j]~1��-�!́��B��x\�8.��*l�ʪ�6�6(Nj?�h�LW�sM�#2I�yV��B����o<�/8�zq._�$��k��+�_�Ö��ȫ;zGS�g�2h,S����ʘ2y������r_������V�'e,��ʶ��sg��TN�\��v�l�����ЁAܘ�\ޟs!���a��Z- :�P�W�Z���"�8d�rF���V�ۨnG�_�}�boo��||�9f�lQ*;j���IŸ i�.Z�xό�WH�xU�b�r��A:�i��3�EiD,))���I�%8h�-N㻢A}t�|���Gi��s	o���~�\��jYd�3W�.hك���PwŞ����r(���+�K�WYy-�lS���M�l�b��(���j�&�A�yL��W5��^dq�]'L����3�)�.�y�*�KZ�#C��im��"�K2�G�v�-�я"�Q;���Gѻ49�i�� �[���6R��ck��dȑ�D�h��u粛p2H6�1���ny���h�^����+��hK�s��8���⸌�D	�L	r�̜P.����h3;�H�}��M�[�U�3���k��(m���=]%�G�<5�t�]�Y�>�j?L�[.�>�*��>��c7U$���]��#���7l�ӭ?y�����o��B����D	�@�΀2��g�C1��:��N��qP��;=�$j�\�b��7VFU_�?�9�+�����Z��v馡��7nGi4��._#�l�d`��T�}�-E�E�	�Ґ� b'�(���\��O���ܘ�iv��ִq����07��D*�k_~|~`|���i7V��0U�%��u=ۓw �?"�X\ï4krg�����Z����Uo��O�x����+�^��M�9�F �C���vS`Lk���h��=<5u�,��2ǐ��g%�c>���ע�d"�����F�m�
����;jx�ꕲfQ�����~[ͫ����y�4r�=����
��}����c���r�'o��_}k���?���^&N��R��]!���7�� �6��g��sZʃb��|������J��Qv���(��Q>j)��87�J���ް��EC�G���p��P�Y��N��s�	E��q���>S<Yy<�� �UV� ǡ��cj�f�U0.�쉗gG�T��&��%��h'б�t�v`��~��n16�&@����(����	 �����?S����Z��3#��Cܝ4�1o|0��v�5�������ֺ94'B�#�"B���9+�1q��V�r
�(M��J%5HN\�ͬp�����'È@و���Qj�؂��e�0ơ��N�պv>
vo�}H9�*?�m�D�j̒�o�����2�:ruǲǋ�I�B��VUvVu����09Fd�^tol�.��sN����q��tn����f s�P\2c�-�2������טvO�F�3�p]% ce�5۶��7Y���9[����mc���y<�^2�L�����(�jr^��������H<�#����y������ O����,x++y��Y��,��WM���qn�Vs��{�~�Z���WMG��פ�lH<��F�HS�d�b#
��q,)c������&�jX/5�ɐV�ݝ��r,�ξ�8ݘ,\� �N�&8	v輪���G����XqR��Ҥo���xP.`ٳ�@�gGE1�XM���ؔ��\�Rez��]O�'��]�s`��V�YLZL�w� >�"х�ˇx�V�gsA��S���)�wz���_�V���#�D����'4��oV���"�����=�VK@a���!^����I�Ab�J��nn��'���ݶ��"�V��`���N��6� �S�	w?bHo"����(Z_���C�^݄����.^-���F�X��פL�Ӏ�|����<���ď
ZM�B���� "KB��ܭ���Ɏo�@Šǌ�P޺�`��u�&U�C\b�u���Qde7�Z�.���r�AV�+�B�Q�;L�@��-&��"�&'�_ƅ� ��F�s�H�&*�8��Hq5�r;��U��Wܫ7��y&��	��걽n�0��5�ڋ�0�s�j�&�4�4{0[�G^$%W�Ͳ����~$�k$�����^�'$t���)%�8��/��x�������@����KL`��H����݆�e���b���kM";K�����@���-�r���������π��>��z_r����t��Y�i餲8�����g��j�I�5�������*D0��Q	@o���~�b��[4��vg����X����t0��Z�^������c+��*4n�^ni���6�Xx�����h�����V��{I[��
�#�ѭe:��|�kh�]٭�����y�]J1[r�(�~!-^�7�vF��[��1��PX���#K��w�(�l��Ш��A�S	Q0H.����[���-4�@��OH��E�����T#�&���*�)*7O��/��=�ɳa���������6��HB�b�y�+�O{
���z�Vd���E�9��VA�m�󘔊�N� w�n�/�^��ǡ�1�k� r�4���JQPz̾��z9`����J�h<p��o�7>�S@?�@�8��%]]\ӿ."�/�s�[�n�c(z%^�4��b͗�� ����"	9No�%�EYl��K����ѻ_�9�����������^fF^�籑G!~L�eV*���y5U��m����M����-.�:
�H�Գ�V/������K@����4Ĭ�L�T�>����AI�	!���Z>Fd�%^{Km\�~*���y���?Wy��?����ԭ���_j��Z=%$�a_S�X�H�����Ib��dud�*+�O47*�#�>�b���Y�:�o��h � =
.t��B�E��q�[�:��<-��K�)��"�jg�h�d�дi `M���������n�]��ݍ�Oi>�s)n�r[h4�(�3�����2j:��Hϔy���_����GIqv&�����Kֻ-a��O^)Rn���6��������]����ةI�`9���[-z&T&�����:����P�!���1���p�M�>.�3th6��t�&z��,RB�?{��0ƶ�n
�\�2��BrI��-)Y�{2̐]-U�R5lv18���O�f��ό�3�N�!kم{9/���w�DtD}���4�����NG���M�;)�V|����2!|BX}β@�TRH��Dȉ��E���4v��U�5lƢ��n�~�Dm^��w��d�a�dVqiF��-�I��x�`�(�v-<�gbq���Ӻ��v��{�$���	����7��A�n/0ƿ8���X�5b�q�<�^m9fZ����g{R��6g�F�?��ƍܚ<]ғ����ɕ��X1��z)��X"`�d��E�ie��JD25�;m����'!�\�A �f�l
������3�FRA^Y��vJZB�ra=�~Q�@ϖHֹ�h�u1���g��c�������j�Ք1��͵�R���&��,Jm2٦%�M՘��O�H�#fP�k����k��>�P�RH�-���4=��nrÏ�?�ߪ ��o���Ere_��c}B��v��Pː{;50n�9�,�Y��������Ԑ�r��v�� 0l�w�A`��8��������2�:��+ ��כ����O��nw���$��}4�i�j�`ur���cI�ahx2L'U5�v����l����[o	��� �0�Z1�}.ΟO���f�����C��f�'�mӦ�_�>wdɀ��Eg�L�6���,Z{�9C�דY_��1�N�D�	S4����$ݓ��Ձ}#ԔW��j���,���f�J������t�訌�-�ރ� 1���Y��T��4�~c�c:�_q�r��zօlY����:Ƞ��P�(.n������Uv`L��<��F4�ݚ�����\.��#��qA_(�L`{@�#�5NqÚTs����^:^SP���hi�w&/Иg!��T��m��DA�T)���?�5�"5,����h�����ǋc�a�2a�����"+��l�'�ɸ�\ C�D��^��_I����˜��j�AF)�*S
�����
�5�4�ƤZ_�N�F�F;�Lr���Q򩡏����j?�~ ��	�d-�m2���p�4�����P�(L�����Э0!���b
����X�X��I���O"ӟ�Q�-g��
-�PK��p'����yU5C���ɽ�,Z��*������lL�bY� �\ES��k�#�9Š��z2�$
��ݨ���A[�/WF�:��eX�b��rR�f�_�'^�:N�;����->�i'����IM�r?�?����|�"t�k���^��|��q���lb�#�e���R �ʴ������
9f�!Z�e
k;�uOO>��/Bk1װ���s��3�X�X@���#s����;D,-�y�^�h�E�h5��=za���b��A���4�����ឩ� �v<���E��Pg,�5~M�Q%ǟi�*h�jr��H�m�����}��ϋ�K�t�7���^�@q-��i; ��"��$nR��|Y���8c���g�4_���g�!�Z(׳R�H��XR����1�r�D���p8u��qt�D ��*s��P<�z ](d���nX)�j�I����6Qҩ��j����|_({�~p����޸��:@�'�J��/Up��p�܊ψ�"�s+�9jOZ����L�Xe��a�(�.�o����eգ�<�/K�չ�E��k�#��F;�4W�ˡ���k?)���S����wȂo�\4�r��u*�b�xQ8�JF��֔^<��u{ٴ	�`RW����U}���q@T_�V��T�ڔ�r.�ã G��|�&�B�*���Vi���Fz��,�L����YW.�GN>�P@: !�KY7ڡ�'N�I谡�6����:O��\(���xb@�1n�vn��1)B��d��_�.�� \�76�g�ΕOb}�'s��Y~�vP9 s���B�6 �i�������u͉hޥ�JﹶSe��� �m�:9s7�D_s|z"��_9gs��}�HhЉ���1�G�T����z�YF-�@i�Y3s�&�>�%-R���m?�ܹ"���S�6O!D�>�5�#2^a->N(�	ũ�� ���
��O!��.xls;6�B�W������|i�Lc/�DaӄDpi�7
�kw�`�Nn�x_o�E2۠R�	Oaf�	?�(j��ށ���d�e}�w,z���wl� ?<+�?Yhٜ��?G�ki:�5F��^Ax���+�g�c__5��k�ڽ?@qOw�nБ$���DAEM�r����E��oA�qIJ�Ȱ�`GK��Z�;7b���\�z����L�+����L��錿.E�\W���G�6���E����ƥ��P���\���6)��;��Q\�����:+���3|������:��0H`����]�Z��Ġ7��n�����%lVt;�r�橕M>���� �H
l��Ժ�S�ry N&����_�O����A�a�_h T.rEt���am�ت����I�旮p�ԇy�f�@m҄���+�Ykđ�nM8��(y�Be�Ւ�/c�ך��R De�K'Io ��|����U�G�A����Wz���2�[WϋE*�*�K/�ă�?��"j<F5=&O�R�j�D����,�p�D�d)���~Eق'�%%X��;��{��M�M�s8�g�����Kv�F�s 7e]�B�X#b��Ⰷ��i��V�:��a�鬤�SL��^�8&RJ�8�{�Ya�+Q�2����sq=�À��AӼfI۳U�B��d��������%&`pk%��U�p�9�'oE��O�ۛFy���*�O��OX(����3��Z� ��H�����@s�����5��P�I~�!��^^A��AN#��"�ȯ�����~��`�����$�� ����9$�q��l��5�MV7��vD�'XK�.z�aU-���y��u�B��R�rl������5(��J�ag"�ú	�i�ᯚ���>�Y�nBa3�:�F����2S��*�ht���;Qӟ(��X��]�4� N��D+S�k]�Pº��x������.����0��\���iM�g)��p�X��q��x���J.
��X�f�UN�t�68��ғ\�$��ƛ��*�l�*��(�6r�V�@-���~zs�x,�4'���o�ט����1;�����KOϸ&+Eb�x�,Vđ��զ�ހ���Ժ�����H�����es��!�"�t�ܳ9�2����L}�Q��8hp�g��X?;��8s�!k�/�;��*���1)jl.�ry<5�jF���%q�
�c[�0��PT�C�kE��7G�u�5��ty��1c�%E��a�5L2>�l�Y�M;�>�ar���/~S �D��4e��h�ɿ�-gb����E5��ܸ@\�!�z���l�ޯ�$���<*���h��� ذ���~���~���;Q�kR	���״k�:o�|�<)��:rw�G(����JG�L�"4g���n�љ榒�@��� TË�[[���,� h%��ܕ���#�ס'�c�����LtB7<�]M���/��b
�����Vs'����蝮6��a�7�_�l�"�Aԃ��h�O&�-������zf�hiD��f+F����M3%<�"mt�x)�IK��y�>�&�g��`i��k�m~��O��J�t��s'I,r����_t,��⸵9o[&l5���i g��j���S�&��~~d�*}��Fpb2Q��h2ñ*W�!�h��98]�fP��jO�7H6�W���a$�LrV�/c؜�+��F�7�F�jb��E&Ϋ͎%yB�I����D)=}��y7z�����3���Tu��%::[`�;pi|B����-�_�Ȉ� ����\��'�n����V�o)>�}��D�=��>�Y2ɞ_{�wo^@f@��������M���W��J���u��Ȯ��(qCy���7��Z���u&0���)�;.��3�0U8Б����jr����r*�LZ��1��أ$�!:M����'��H�1G�u>A����`�a��(�E�&�g?0���G���b�vZ����e�A��r	�2�h9�+�B�U�~�XV�����ǰ� G�H������hw�v1 `@aHЕ)a��u�ϊ�ҏ��H�,̨��d�Op@*/e3_��4!ɉJAU��!2BG�f�#�{\�dMe7���;̊FQ�ЗM�rrH��*]�q{�&�K���˧Gc1c\u�,�e�È�vq�
�?�+^J9c��Y�>�X�׉|\Ύ)v+`��Yp�����( G��!�����3��M���Sҍ��K��?��/ڍ� 7��o�xb��N��k�Z�9Z�XG	N�-��c�t��-;��_2<΀�=��f?���Ca�,�����;����P x����v����� ��qX�[����M
�$ʸ�\b��D4�HQ��X�L�*��;��$�ۛ}Ƃ��2r	��߷f���{��P�y� ����ܠ��zO`['�A��)���eQ�v$]�����ס��d�Rn�M��])F��2/*��w/&�D��G`J��V�n�� L�x�-WӜq�k���Va���t��.�&i���
�o��W��qXq����,�9!���B 6Aa۳���Ɍ  ׮M�qa�W�!?hwA>������q��DޕrO�K�@��ۣx@)���0Ɨ��Yuի��8p�#��d��nEێn�>�E��w��L��o����'h���wmuZGEh�>-5U��,_m� PB+U�����FgE%7�&�{1t�y��줮?�Ep�N���"�7ç�kFa�Z�%?�֓JK{��|k��$��/[ip��z���,m�(�<=�T��&�%
�FuA�(�T��C���d��D�� ��o9�`�8���7;G��Ei����"��/��<�$��y�J�Zg�����2��b)�c���p�[ ���^l����=��#I����Q�R˔>>��Ope��F�q���xFNSH*�h{�aE4]����h1@���VK�Fz���a%���b�޿j/��{б���"���Ěwx:����5�o��}AObG��""�!��+�t i���_��6B���ʤ��]H�^Z��&�-z���F�ҏ'��g���=I���#��p/[]'B7&'��C0/(��9^���=�����O��n:�<�[��������U��N?��%��)B~:�W�(��֥�cCvF�g�IڌZS\����U�0Z�>T����ėX�>��9�}��O���}¥G���B�+jd_m�����8Z�q��.R�4Nt׆��GB���4F���D��W�2&L����YCd�-U�Y��;���E������8�A��P��3��1*�{���7(b|'E.�M@T�>�k���k����tS�(�m����ӄ���V`��T�I^/����m|J�I���k�0ӻ%E�)�1�|�R��5()s̊-�X���_���&8Fn��4�}���t��8��P���U�E.,)�ǥ�/�vGl_%����<OQ,���S���7��&���Nn����Ԡ���b��바����n�qk<sF�&}�k���������-`���L�H1��6�5c�
�l~���������x1��R�|5o�.��oc�f�3X�:�|��qل�S���h'γ���)3?�تq��J�;r�^GĖx�H�BA���]_�Hи�ưbd@��c>�&��З-1�m�I�t��a+Z��|2� �Ǳ��Sd�%�Z��I'�`��������GY�d�qި���}|H��Z�aZ��O҈�^R�t�R	����|jT+�V]�(p��kT�m=S��Y}gs �ߢS=��}�u��R5�6Z���3(�@y�-&���V�pć��F�uʼ��:M�8��P:.���A|>�أ�s֎D� t�|�n$�d�?���܁�q�#�H�I`Lt�����������+��e�%-j���u�`�.�{��ۖYK�h���O*��a�A�~�B�%	������[9����)Zzr�g[����	�����Y�"����n���1�0��<�~͝����D,/�w�i���ԏ��[g�s�I�/��л�hH{��r���341Ќ�(��3f!Ǌ��6RO^��1�/g�%Ҽ�x�HťHe�\�e+�h��4t[�uL^L��K���)�Nd���V�m��ҕ:]��P̆T6���4���X� �W��,LQ?�p�E^W&H�6�Tb���ν�|08%	��{,Bc�1<N�b�voA���S��lL��5i�Z<�XH�L��>�U�E<� %U��b�a�j�����^s���̀��cx�&O��{>����g��a��B�d��(r�y�ROV�X��Q��]�R�=ٺ�%R�wob��{�������Z�ܻ�s� ꃔ�z�*�tt ���(I����df��c�7y�Cb�z ���;��<tU-��١����TљZ�򡄙��C�BS�JHjy�8������n"�f�soi;|��3�X~��z��ֻJ$�\�Y���{ԹZ#RN��h����R|�ɴЇ��T���R�"������Ǡ��O���־�$�+�Pۡm��vDX@Uy8��ӣ�+?8�y��P�g'�c��7i��"s�6.g��Ȣ&i�
F�X_y�8Q1������S�sq���1��c�C`�]Τ����$ÆY,����F(N�oS����SY���d˒]���G%�C��X�%XR9G�ɠ䙓S���E<W�e���x`��[2JeǍ�� ��R$J85\�f�����P���#�L��e�^=s5�ʈ`�c��W0�Y'o�"�\N��O�唇��#V��l�GG�N��(��3]l�@
	~o-%� 2�%%�S��&��ʨ�>l�����tS���Q�.�{��"U��}Z�&ddX8�,���F��N[V�N��b�(�G�\�b��8%�K�d2����؄�g���G��˺V��]�]�p*�K�%ۈ�Al���~�C��Fr@r.\�wcI�^v�}��|���!��]_׋(��'�����g�@��Y���d��0��#{�[�L{�a����� �U{�܀��Ɱ���H#^�1P7�[��p�Un�RQ�l��B����5!��~�*�������<�T���%�1<��狱2&l���2K���Ni]���e pA��r:=Y�+&:'�̉<����n5��M�9��ȫ�A4�~���mv-�����~a�K��crttO��za��t���,}�_'�%����(Wb�N�����	o�f�#��.����8{'5���9xl'V�	��\�^r5��J� �u��c�vǨl"a��s�5��e�T<xm�մ��;�������Ct��m1.|����YNx3"я��Dz%>oT\
Q����ܘg��q�X6�"����C�@O�rDS�h�R��6�Ü�(���o����Ș�l�����]a��?C=���N��MU�$�羽�ä{��[�o�j��X�rU�?݁u\ǿ���3(�F����0��-�7J���+�+G˃�AJ��njB�`���6��9�靮@!|#y�������&���o�۷��h��&1R$��8��Y�N��p+�a~Z���xrS��7�hK���+���K�V�ۑ t�A�	��F;�,���6�����-�ɇuR�4�"���exѿ����W�8�x���ʟW�z7�Ir�6�oYL_���-
K*�>����=���#��2#]ڢ���t>��Ƕb���@8��[Gp�`��@�s�8�n��_r��k,.�k�+� |�:6����R�V��0}��TS�Qj��J�도�	�j��	���2���N*l����6@9��f�0þ+��gf��&���͂�@B3�o�~	y�	�ƣ�8�uUW5�׾�VC_����xc�a×�҆$J���U�\$}7�w�yX���:�*g�C�I~ܝx�t�`o����]Q&�S�?�/>��_"dR�`�� ��p�D&�.�^L%X��v�3�Z��@�=�̋�.#o�j�x�k-�.�N4���C/n�@'l����(�kn��X���lh�q����C��?��/�ikXEx�"Y�]˹�9>�/'�E?����tt�,KK��6w���i8�).a�o�Ic��*�U�*�D����l�~�w��q<������ɽ�N�^:S�L䘮}�U�M8��}U��3�]
��FGw�?�#.��/��0d�ŨJ����o���b�o$����2{ͤ�����W�*������@� \Ŝ9��;8h�&o؛��.�_W��Zr`��H�}�<��g�Rp�����R8l���a�� ����-A��D��hi�\[��$vEg�?��d�T��`������'�����ف�+ӳf�rY)������H�PpX�Ǽ�6��p��b��7��]�Osۇ?�J��b��{�ѧ�c���	@��8��uZ����������ϞyÏv�}!����<���_�}����#�1/��w��h��M9r���E�bE�BY����Z$w&b� ��XX���H�K<���4�׳�$����/=U������zf��Ya�q�2U,�M�ou��?5�?"�u=���`��I�� ��&�����G�lʪ%Yw����)D�j'�4\t1K/���[E�����<�'g���hA��K�W�Q\S��2�TTӾ�'KKVc2�8�0��\[���K(���G�-�]�Y��q���q�#Gú/.��n�v˸S^G�:�A"𶲀 "H��L8f�j�)���WV�k5����:����(5-/o��lc�9�A�3�0v�A��q�IC����=��G+6d�JS\�)�f�)�~�}���؞�C�j��?�#��AT�w�٦�X�*V���Ak38t?ol�0m��E+ȥ�>D��:4�&��xs���T���/��D�\uh�o)�f���f�vЊ�oM�U�0sn^��/ B��e	]?��(��jG�.u�:m�divӆ�mx����HO��b��d��,wjkp�ut���s~�����+I;6-��?ArG��Ⴃ-�_�6�.ܯ#ixa�"��\� EÖ����RS��y�g�b���A+�D�Enq���o�MJ��=���*�� ��O��,?�e�B��Є��=#G`�i�3��>dL���^�#��"-c��Ѕ��|�3�G?���f�|=!tcR�e+{����CU���M�����Q:C�:�Yض��ڟ>ђS�d5�<�nU$��jo�����߿nbC�����	ѿĿ��L��kb�ޝ���C�����g�$$�ԇS���'A���s���p.�K�b�o�Rw�13�����@x��̌D�Ԛ^g=�)��ȿÈ���F��b0�70�j�	�]
�S�XVj�ʫ�����
p�o��TU%y_�g�Ǩ����Y_a٫]K��������K.�d��G��}6�A��D��� �*j��O�aR{p�؛i�c>�9(M�w�T^�<@��9��e|�F>	,s���P�W��Q�o�[�7R
.�FZ#ł~�,�'F�h�i�U�Z�<�E�PuS,S�15G,����i뢁�����I�J�B	�␃a��ɚlK��*�^RTOl��K(�Y��TA��`��A7�Z�t0�G�s��+��b��.�)��E�H�ؿ�ۛKB;:i����l�L�t��1?{�wXw�m�S�x�2�e��X���4n~�CUPͽ̛s/z��M��6VK������|��3�>:P8�ꏳ�	h�)v�D h#!�� e(A��(�AD���Oct) 5�G�/-��eI��ț�g?��H����|iK1��5F;�mMo�Msu?���=��jt4�#�6�F�4���-��t?�D����ky�>��ϨO '-�.�8<~�.λSk:�Z�����}�`���R��,Ha���ן�b�^��Τ�xK��6���g�;�ݘ�]�)�O[l�2C�_OO�BEx�rRe�c-Zl�ҝ� ��V4`�o�7^k��^�,_��F�r�2�=������R��\�HL���L�Q�y�$5}�Fu��E�����;5�#V��x�=UU�����惑�:iz�(��6B>�e��D�v���sB���/�'��KW�8���dp�L�����_�Ѩ{?��]��R��v��9��xu��V�H{�׺8�&m����gb(1��T��<����� NB<Z�po�U�hzh����Z1�%p�2��DD��b�L|����U�v�c݉�uJ�	��<�m����{���,���<Gt�P5*Cv�@x��{�R!G��Vhr�t3w q��3�4$�eAm]�v@������ww��ԛ�-5���r�`1 >�]Cܴ4{ѝ�?��~N!��u"Ŷ�KN|����1ag`��Y}��4�/�~��aN���5�rNO�v8o��K5 ~�P�7��J��6��׆�h:�t���y�"�)l����7=L����ж"ZW-�w���\ՌiMc��O��i�w��w쮀� �)i�_��J�l��NR`@v�{��Z�q*�ZӏSo�K=f,M��/c%.6�W�rҥ���(� <h�T��^7[�f��Y �(��7���`68kl�#~A�C�������sNA�,�"�G`�0���O�ƣ�3�(��\3I��#}/sb:�kUnط�c㿙��E=�0s98�p���_�V�0�J˯�9K�ۙ$�Z�tK(ne�*�����hh���1���h�7��ewm�8?z�YZ��7�$�kM�*�v�y\�Y�R����%�-��g�H����C���m���	6�Cp����2�b)���o����ъ'��Ӽ�6ڿc��!��Ջ�F���5�(^$��,�²�#��7�:�V�8����\��_����Ɗ!�5]��t��7�:h���q�_<����M�^��2����^�4�G6�ڐ���/ iQ�֟����?`@�3v-
=��~�TA�{zIWԗ�����r���[y&1�_���3�B�!.L��@���ϧU3���K} {=@�@���7�7YW�m}v�\�0C���O^j��y[�QՍ�)}���*���(�˄�Ix;�Bu�X�yl�-k���=񃨧�������)�����)�Gخ�`� �${4a�w�h9�����;]���L~���ԇ5�u*�vͦ[�< H^ҽ��R���y���f�dg�j�u��f�PF>�"U^?=h���������v�VŞ��ݹ:��~��Rl7��wWq0��o�o��=��0V���Р�X��2�����w(��Ts�un���n>L��f�}�N!O#�ʺ_� ���K����;jcU#s����X<���_huHK�m(h����nES��`��$zM��S�8��Q-��aRg����ǐ"%*���g�ƻ���M���6�$�" z�16�$���	b'�{�ҁ��@k#�RA�>���y�h(��GW�}0"N��Gw���W[�~䷞5��ӄ�lÊXv���Y��@,����)V4Z�>�-��a�A+9.0�-��B?�ߔ�ޖ�S'�3,Q_*���&��������كS�$�Z��l���J.��z?�I3��=�o��H�,?%d��3,�9�����}Ţo����ޢ���Wʟ!�Ӕ\�y��NR �!N���d4FE�3����(����[�!Q��ـ�ג |5t�C�;H�*2+��T,O����op=�׏
��L?/��҆y?j�՗P�>�	z}�Dq?ǿ�|2�m�`!F�DTX;�ÍY>�����~����Q9��wL?�v�7I���d_ �j��@�J&V�{��C���]e���?P�ͶOIᐬ/�q�I��Ǘ�b����T���.~w�69y)8e���[�S��)���^D}���t��D���}���
�G}�C�n(KȚA���Ua�
���}�8�����%+��|56�P �qw_�(݌m���qy`Ӓ1N�����`���Z�J�A��$�#��<rV��}̝��]�^�  �E�S�I�Ҕ�%}�\����T�學+��SB�q=S��CcD��vrʋQ���ĮR����Z�j�]�qba݉�v���z� -���f{����@O!�ҽ�~����ԟ�|��tJK���Tƽ������$�`�D��ta��:�N� 3/:?���tз��0���L� ��b�����	8�F�uُ*q��.~�f�-��ʰ�QM�ޖbV����t�ܶW
��'%;h�p7s�FS��ȾB���!I�;ӫǗY���N8#CB��K��W[���[�P �5�}�*�6~X <�sZ@��\���@1�NAi�y �!��Aq��X*�?i8Tn��S�� ~���$�Q"��3m\ߚP ���y@��d9v��kJ��9 �q�\n@��D��5�'J��˺����p�ĵ�|�5$,��$ϐ�Z�.j1q�B�ũ��7`�ߞ�ф|;������{�v�>�=��e�y�.��Å~����M��������k�	/ih[j��"�����ƅ��a9�غ��<u*:0x�r���b�����1�]�!g�t��(��� �E�t�&9�,5����/gx��CrlL�lr�9��8g�����y��L�:ن�H���%/lU����H���Ә��A2��Ƈ�ע��(E)Q���P�ɱ�A�J�,.kځ���`?���mYنa�9�+_�����;������k�b.[��n5��3�9��y	e�7��4�s:��v:��n�s(Յ9Em����McP����_y�3��M�t���� ��FB�߀�G�_W�w��U�k����{ӏJ�F�BJ2�9{�/����6G5Hq��=�TA_��w����"�tT�$kM7Ѿx��F�T�[A�m�~�����T�� A�UT7X>}#��n�+�\�[�oѮ�e��>�	�Te������9����t��Ҹ<��˙��@E�-$�ث�}HD�t27Z�C#�Pl>Em�K{�>���V)t]�����.���U>cU�"�vQ�%uz��a=���,��R��v�W�z�{b}��{�4��1S̺�4��Ӭ�E���@�/�����0�t9�nmC��3� B(��lq7�j(�����zcg���VK(�9��|JJ �C&�7a'�~ȗ޷`�֚#�ɔ��5�ٸ�cX����x+���o eqq�`�+[�q��������Ϟ��w� ��~��&�
�W?���8?�0��
͠�5E�,aR���O����Yew��$[bi}��@K��<�!�(�Մ�:6���-> <p����sWc��S�u��/c�A�GO
�g����%\udnX��YT+��t+Cb̨~���텖9����3B���}����lah���>yd��䭘�;���;}�<)y(�mZ�Ǹ*�>������(�+���0몦A�4����?���6���³x�:L|�éX
[,�?��Y�HN��E�j�陭!s&Oj�-s����p�jh���$bK3�o�&y�&�;�A��UǼ%`��@�ƲC���j���ݣ�X���n�+��6�m�:�X�Ju���dg(� ką]_�)���H�I%4��@r�JH��E���8�>C�Z(�'r;[c(@��?�x5zu�uc��6�R�|��?w2��h��{Ɉ'/`뢤Q[��^RөLX�d���u�(O�.�_M�p꼠�K�S?����7ݒ����gn�9�9���&t�ˬ����zs�Qs"�ǩ8�X]N��m�^��uYV����9�ݝ��T��)tmZ�x�S�˺Ax��)�eAˀ�LR�Bl�T��-���a��|��Y��ѫֿ��=��߀@����H�h�*;Ƃ��댴�SZ�mj�λ<[��=�fk>�!�-h�
�܈tڞ�$	��E~���;�>H���x���e��B8ɣZ�J�,x$7j�6����/�i\��b�?���W���A�o��(���^!$M> �e�F|�X�?[���K�gw���]��!
�y�2jo���:.�p]��W'�e��}�o�K!��׺�*3gYRc�G87� s��7֕%���N�<׏�����:}�Bl\#�x�e�7	��^�b���;�=�����G�^Hx��M�����#a|!2�C���g|eۻ��?k�j��&y50&W�8���Vں٭!�=�q�Ftpw�^�z�q|���{8��Q��h(��������L�zq�l�vu�U��e_Z����b����6��O�5�g����5����ty�B��UۏE�8��U���&Z*kC�X(]@��끶qz�%�������ϱ��O;�U!s%pΟl�$�2Q�g�H��I#��,p�-$��7��c9��b���|�;LY���2����]$�Zڼ'��
QU���]C���|�Uɟ{6*7����}m61��M'�����W��U��4߫�eL~i��a���0B�
Rp(�ͅ �~G�K������2z��xW��84�=�n4��Y��類����`����m�S��s�3�����nvi�u�7R�r���i(=�)�@��^���A���Q���?�rg9C=��ę`;WT�zb�ٛ��o�\0�z�T�#����Ď6C\qkJ0�V�⌑giӑj�Ϻm�q�'��?A�Mc�5ט�'��=f��f�`g����c�������G>�4~t��9L �=�M�+G�߉vGN�	�HYh�[k���͛E� ��1<��i�����c�b��&�:��|�b'�ƃD�irR�?$�� ���_u4��ADn�U7%�i�PK��mR��Nj��c���쯄ך*�	�.���47�ǡ
 �o7�:��E]����<�3<��I�?�gh��g�M\t�1ZY���F)�P��� +� ���Q��pj(�u|�AwH��j �L��ǃ��T%�Ƣ{�m��͚K?/@�8���շ��2����=ȹ���B��1<ĥN��,�(��"�f5� 2gX��[�w����Di�@��y��'p��ضe�h*Y99G=�)쮖Qp}��'E>��Ԁ^�;#}��H�*ג�lYܶ{�N�ؼ����_JQn��+A�I�ޤ7� ��^�5���0>ɑ^@��w�. ����j�q�����e�=�M﯁����<��$N��)r*g������R��9�F�_��}�Sja�m@�;i���X߃Ć[zw3ނZ��hA�;��ݻ�t�v3�,"q�(Ur�U�:���5���8*iU��4��)�_z~�ύX-B����
�}~��ϐnF�>���t8�=Qwi+��Nn��^.�d�%�j���C4SH����NM[��5P�)e�~�a�@���	���{&&#��}��ը'���\������"-�zi�Ȫg	�(#(�:�?�ez��r�ǥb�&3��˖�IЬtTJ+��~��tă ��n��me)�V��Xީ��Y�yw���4� �+6��)��;�N��#�����[)Szj�W�e�Z��=ԛ#w�NF*���ͫ@mM_�QJ�z~�Jڹ\0�H�J��)�4�<�׎Fq��
^#���[�p:u����%�V�f7�
�NA��-�R��wz���C�$NS����۹�A�.��u>М;cC�r?/��b�,�k�g�?z 9h�Z'�c~Is�?q��G�2��
^�@�[��Q^5$X��b�9����ϛ��'3M��?c�ZB���a�M�q�)��#� �������.���DRV)�Of��2�	sW�Pv^�Dڸ��(�yk��h\�U� 
~�w|�ao�E�.�>�F����u֒�*~�J ��q��C�;�3լ^���a�\�D����)1���貒�2'��{%�=�,�h��X�������Q��TZ��ȧ�7 �_�7	B�D����;G����0*?��<��&���I�wA��: !��G���z�D��-J�c����� �xs��^N�<�������b'�ʭLC�,�}���?�$�?6H��x�u��?�Y+O�9��k�G�B�!��.��7���@q8�C��<wk_��(ӟL���_�9�s��:��|.�)q�`B?[�@2X�4�"(-�����$C
�p�e 9�:OZ>�~ߍ���o[�wvU8%&����+�s��6��Y�ep�$�YK/j-H�f.�NUz�EX��_��K��X�	\9;Z$�)/��6��+�&#񆇩1�=��ߩ��g���î�o�YbI�0�z��U��֘=g"�Gw������~q3��	�\��'M�r��[�Ӛ�q�����6(��JBX�w��Ԧd߼����q�8})"�����lv�^���9�kG6(��T�b�e/\���Y��e @���X�l2ËM�LɳJW����Үg�����.����d��y�q��	��cʅ$,'p ���� ���A{�D��äD�A,�TN=�s��[��Dk�y�d�]0���3���QͭN�w��3�gM�Bt��;�#�6��Y8��?V�D�q[=�����,e0��^|�����)�Oˁ ?�<\�u`q[�/�n���I?��e����Q�Z��N�'�?љ��L����E5GON%Ԟ��&�Uk!�����M�O������6�V�K�V\u�86ӊ,仗uA
}G�HUB��x-9N�3�R��d�#5��ݣM�e=c�}z�����F�ci�<�&���՚���ڑ�F�����a�d���F;�����Jx�niJ`���*��,�x�-�+J�z��d%�PU��4�p�;�iN�F�I��O7V X�3s��X��#��Q�cJh��L���݀�J>�����Ŕ�g(��T���ۢ�iT���n�BJ�K�2�����r��~�����6��u
�Qs4����Bl�p�,K{��"�!1?v��7�:}���t��֠��#L@l�������}h�|��rN��m)Nǈ������Fl[=l��J����k����׉��, �m<*"�}^�d��5��%׹�@���T��e�ܩ�8�����c@�)A5eO}�Zi5�rN�����a/q=�YF�ՠVBQZOP/q��f�Q�<�����y�]֚���y�a*�vQCұ��yuK�^;���23���+�������L��~����.� h���� M�G�Yb���`�A����Ju%3RJ!��M�.cE���ؒ�19�tJs��߁K8~��S�fѷf?���A(��&� ���)�bv<l��-DGi������ӝ����ֳM�޴�d�{w<Ƹ[OO&N�}v(|C����o���Vp�7\�닅c�����c3��:N��n��_>Y&���s����� ��8�L���O�;���o���#ĩD-A?��iR����;�ޣ��_��'s@�?� ����?�M�9_Fa]D��;�8$���G�D��΋�
i���h��[)�B��a0��~���êu�����^iV3�ۈ��r��bZ�X��%�{�0>;�w�^&����\I>��f�5^s��B�p������Ե���u�QRV�c�t��?����d�'��"�N�<i�������'_�+_�b�2u�������5r�E�+烜�y�M������A6W���>��K��\�ή�v�n	Y�̪@c8��+��A��μ���U��b	\��t�1��7�$6�pJ����
O���H����Z&-(6	\!��pk��Q� �%�~E&ޛ��>X�O���?�d$�� <N�č[CN����fm��D�a�����_�)�U-c�S���������,��c�2�ܓ\Eؒ�b5�#	� E����0�z_�d[U�:#�!G�-���W)z1���\�N�|h֙w�^���d1�6�u0�
�RD���V���YI��,���7�&�)��$W{�FdbIn�6�:p�]���^�h�C�[0~br�LCI���8j�������D=6�F�ݘQ�a!�j��BD@�r���+� �{�ޗ�a���X��Ǒ�X�q�h����3�L�$�@�F,�X��N�;�8�q��4�/(F[�<�����Y�S��{:�G��&�Y���C"hr"���q���P�����p�5���+v����8p���D���TfŽ��zP���k�P��{2�
L�)�׭ڀ4���P�Џ/4�DVu����

�V�L2pֵܼ��,-����&�B�K߽k,��%n�S�_e��q��!ask�!�=素+�ڗ���K�ʝK��W�̣�&"x�"���2�#�DY�eF��̞���m|��d����>��A��Xx��&�k\�3�RGӫ�ۏf��i42i⇕�"հ*/m�ǹ�ڻ��&+���_�$+�	HB?�A�I@���}·�B�"-��o^�j��ē��b�eV�;�Á1��݄*�U)J����GA��,�l@P޶����C�޶#`�-��n�GX.X'Z+�`�����X��La������y�>ֹ-ו���TD������H�"PR>0����t;#I��1�q��tQ��q"�����Wޛ��{�>Q:N�a+8�L]�t'Z��5E}�=�vT�V:)�����~�� 7���v����EoX&��h�.k�_]���V���ǝ��|�O�����]�F�;�-j�ҸQ��I�y��h޻���߀�p?;��5$u)��Y�;�������L�Rt_���
'"I�H���E4冟�Le�7'ja�X�x��Pt�����`�����:}�C��v�?Hqr����dYkc������pap�-��QM_ ��`��֦�l�aЧ�m��!��{�͹�-3��:wmZCpy�㩫��x�;�ͼc��G�ޱ�8�}ד�~���/�)I����M�B#Z?��Z1����C61��jߤOh0���"$��bOZ*k���DQ�����f��R�~��j�,��?,���rym��l^䫷�[!	�W�ƣW�D6�?�~���B�vLY s^� ���[>1�o*�.��[m��'K�Q�Ą�d���Ѵ5��*�;N����U/����zm�2i���	T |��Igix�r{@��0�튭�,%w]���4I.;�؞��i�W��������*^� ���[�&���֠@XH6?��?x��HG�(�bPS�Gv���9f�%��!{���vec�j��CU1-��S�p�~��
_���d��el�u�?)���o��*}'����L{%0�������x6�����d�jIdn������eT&(���3�>Cޏ��	 #N�L�B`	rt%׾,e�}�yӐH���*q��t�O������;� ]���c��@S�br��z�(x+�/��ј�J������¬m�&0�;5���sS�@�?��$v��IfOo����"����he�L�`/ͷZsI��1^���L�4���������yU��_�A�,D��g��P�A��"����uލmO��"\�7�;�p���)B��9�����ī�4�&��$c�V�)� K��%T�>Vy�l����6�Ė�)18��I*J���w��'�Z�n��/�%��*]%_;D��P�!t ����ad>Q��wgx���Ռ�[���w�sfdt�B�U<�*�|"_#�����+&�H�Uy�# ^*1�j�W��m�4Ÿ��#l}qdH����c EGk�EDk��6Q�`��Fբ���v����sf��=F��(�-��k9�5`Ҋ�G��gp/���"���}�ݜ�@]�%������f"�R:�)Af*�`�ɻu}B���y�*F�*?k�bsM&w�;���$�
��뎐Ere���ףQ�����t�� k��+�
�o�dК|�Q��] 	�j�|��~�=�튶��m�fP�I�����eg��p�����>w��/!3R�p��.�pܭH7�-Q��,��(gFGJ}CG��-�R�%=VR�E���)�ꩪj<�A)���pX� �a��3� �MYn���	&�a�l�T�旒����>8,��Ku�`�%�yh5�;D�7��jw�0�o{]�4hU�ǥNy#+��w#"�s��)!���}='i�R,���R�j�EYk���P�<F:�a�2���?aZ�S*��6�����ԋ*�ߨ}f��6�����f4.������At��xMv��L��
��-�C��&=GO-����?��ۙ��ڼ	�EpM��;>$ܪ�Ve����#t�(#p�c����*�b�����bfpp����Z]��L�p4�@����d�|	����Zn�/��_��Etgkc�~W��D)�'J_
��b�n�ìK
�ye���9o-�Y��I����هr��V����+���`>����h˷�E�"�^uN����ϡ��sq0�כ7
իO������mݍ�%Q?��ͦT[*N2�!TfC�̵���x_%޶���X����A:��]|�Xp����^>	2��K��ĝ�������-�Y�:�ƻn����C��]$(�H�F�D�H�
��W�*�N0-(M����DD�|���<DR+��?6r����
IQ4XE��+��=� ��W�xhu�!���� ������Cb2^c�.��0� [t�wh�-��>7�OG�fڃȥ��;O��暰iץ{E�A���>���"w�]r(�?�W+��=�[�P�FSv�
�փ�Eh8������a��!�|I|L�?�aPI'��g�3�>�k��<�3Cvn��k=ֲ��܈����R^%f��~gS�yy9��Ȱ�4�r-���D&Ktetl7�P�,k12�0%uϗ�V6�1���ݵO�E[vu6GnPP�Hb�>�_�k(��ū��ti��"]�/��f�q�.A��B�Pq-��@�?"�dV�3?)��_-\��Hg�٫ǋ����}E�$$����]����?�Fg�u�7�dBˋ)g����?�E��	l}*ڗTr�t����/�����O��Me�!���L�H#��H]�R7 ժ���l!`���./"b?��ħ�S����"�o�M���z��k�S�2� ���Jq�J7�z�`ia�3>��Ð<� ��-k��ag|�K(o*/��a��f%���9}zu��@�ح'��]�2��UHCF��v�B&�;����\̰������S�q6��e
^S/�����Ɏ����mK��MAq1��V�6�֖K�6A,���/����zKޯ���������� ]�=�e�$"�^oBH�<G������3�5�>^~�.��%�y8�}��(���x��y��Kn�i��SCr��[�4�,�A �M۔���#7���H5�[�A����j؇�K���Hը��s<�9��mS5 �gX[D��H㺮�2P��OO���*��w�R*�1�=��|�&e�� U܄�S@��Q�-U^���D����u�a�+&wA����e��U�	D(}nćk,5���{�n����q�ߴ��}݌�T[�K}�p�׮w���K��D�|˱��VKؗ�u���6T��WC(��/�� 0� ��*l9�������o����m����}��g�E���r�T�Z�(�=� �]�-x���a��y�K�	\&6>)���k��Ѕ��m1#�8�!��+��^}������Ll��$�S�(�o?Ƨ�ݩL=��/m��ĻR��yH��M��0���Iw�ͪ6 p)���6x�VeB�u@oo���8�=�澙.��Lpe���qFW�(����ş���|����AEL���	���g�xd+�I��cz7Wئ�R���
o��Z?֢H�QJ} =�$��T_�f�bv����� pS�m��"Q��k4�1E񿧏T�A����o�MG7K��]�?m�$g����(�^j�#����@�w��,S�����⻉A���M���
� y��v@���]�uR�^�3��֏�I�G~��$c%~s�]d������
{�t:a������tȽi��Q�L���I�ЅAG�:�s�b�	��Y����F�`�»��H��Q+U� #��G��Z,��=!p]��.�%������(?>���S�S��p�|K�$Q�&	�����:�Q�׺����T�x�m���8�鑭 �5&���U,�P��//�LIӟ%�_%�������i*�EI��>��g%S��>icѺ ����1��%.F.N��0i��w�Q`�e���O�:0�Y1��_!���I��|��3����?FM� �\���s��\�j:x��<���p�;�A�д�7u���tt�����:������ßKn�9d�:��ٱ����/t1et�n���q������,��Z�? �.d���:�\��Rރ���1^N��d�g43�N���0!?5X!�̰lE��Q@~�j�_����L��T��Z�<���b��ۻ��O�Od��bmp���>�uG}u��FCo�X���*�N(�e%$���^O6�����DGJ�ؗ��(�)�Ǭ��O%#3tbh_@���(��VR1ǅa�˥�;�Z
z(2E��2�^p�=�V\'PZޗO�ⓞ�?�wg�����3����0!���1�3��܈�¨i��J��?I��;���Ga?�3-x�';�dʦ�l�"��
��%9�3oF">%��y%�E�yŬi���$�x�����a����[��?+�KZ*����F=�o8����Ҧ��ّX��A�l
ޣ�`�g��y�̵g>����u5�Bl(��@3�
���j,���ǡ�Iƽ���vʼ8��z��H���P��[��	,���\�D�Zұ���T~��ތ��A��Xm��=�[2܁�?r!�#QG�|=��6���9ʾ�(Q�W�Q�wD�����u	ּ�ZZ�� w,��,��M`@�p���TW~i+�}�܀~o�L�F&]q�^�zh�"P�V׹�6!���O��T�������D�_�=8_�pG��0X��c��Sq��M��<b39g��>)��'�:5A�U��M��LYi~GKC��EM�<i��U^��|�żk��1��T�8	����x]\$!�#'̀q�+3R<���ٜm�;��p�2#>����}���,���k��>tԸr�}wB��jCb=�,[�]<+S�шy���Y�_���e)�$R3�$��v2�������*H���v?�t�쩋[to����¡<_��-R�v����<�R�;v\�Xό� +(al�gaƭL�O�Z	mPw­�4�X��f�g���p����	�D%�����{l��R����0��+��$�RөW���C��N̔�ĖpӴ��rV�v���0^��'ш8�g �mqرk,���"��!�����}p�I5�o����3��D��%:얈�]3��Ѵ@��9X���`�i�����~��EZrj?C@�BN���¾�����I�$��s���[Y�0���[���k��y ���۩v��U�A�� v`��A�[>�,A�,X��0�%-�^\H��$�\;��	hMgd�Ay�/�c�ɾ2P_�yT�Rz��j2���R�����3����eQ��b�߅b+�`~~Ϯ�������?��!�^Y�` �w�Ht����N7z�?�"we�����\s�K��������W�犴� Z)T�����	E#��n(I�-f7A��&`ȵ����;��(?<E�ҍU	��o����-�:*�eAn7 ��&v�Q�����z6�G�@�c�K �A�4�}n@k[�4�\7��ʯH�Y���ʏA��b��t�x?�ч0Yܷ팽#L^Ή�L�E�k��Q�;�]1U ŧi)r|���F-�Z��:|J�A�ZeF���1�9����N�۫"�A�yD��!$�t4�"�0�E}���ԎD��e7D����x�뤇������AD{rSF� ����-\��?Y5h����x�L�ט5;���R)��8�}��B��8�k����y�U=)AP�b�$БW���L<C[ʉ:�Qdg����w����<5�f��U��,~s�r֩~/�1r���"{��$�����h/���/�	;�v)���L�?nU�%�ć��tO)cP�*Uw�Z�Ύ7� .(\�L�l��ƢqS3�t#��(�!{�Eo)�Ӄ���-��S�� �B���N]3#��o�*H��JYc}��%��X�e#���F���!�;@x7`(�,�!�\��I����2\HR��i���荄��r�����]�'����˲�[T�M��4x
��5vu��$�cY�`�6�10����&�4��^+r�iS#���@*�[o�9K��:@&0��Xq[XXJ3��*�?O�厜N�-K(뻡�e������� V�n���j��qH�E�K��B�h5�2?>�'OMnօ�9�,z�%��HA��j!�?�J�Y�
V�i�ǯ;�����U%9��뻸��yہ����,�.�)F6q��2�@��"�`]�j��"�|u��7e@Y�k�ܥ�X/Q�o�Oh&���SM9|����J����:E�<=o^Y��k��������fΊp�e�Г�+���&av޺��N�%.%���P{3s!8���ǌS�8�͑�3S��B���c�#��0�sCoّ�nB � ���2��z���IF����V�w-��)
E��,N^���R�W7��t��)/BɆ�E��k��ٳ�����/����>r�@��ox	 �����H����"D���DL-�VN<0jq�l�����z�[@��I��A�{̩Ys�X(T�XɃ9��^�u ���FK˟5���N��T���HZP�q�3�x����6�4��ŉ*u�[���4����������A��.�O�I͇#)v"����RW4�U�t��W��U��/r�t&��+�DY4���SI��P9���dO@��K�@�"Z�7����'��<̧�^�Տ�FΊV<p%� +�$p,�3<�c*���ЈT������L�"�lu��}P�����Q�V#�8H�e�x�����i2�x��-�F�3w�9��I���� ${ۓ�4wzA$�nU�8R}F��c�����'�{f``,���(4�?&�UġI�~��9�_��|c#��k��U�
��Lz���k�9�WYq�.������4����9��t�s��n��D�K9�G����e������ѐX�.5oxfIΚ-�^y4}����>�{�*)e"6����Q�F�{ӄI/Isd�LC\l�E�NV����_��ç�$-
=��Gi�#��0\�k�Dy��K( ��b�_Q0- ��'^�H�_Ĺ�;� 6-]O��g�fJ���G���ŒG��9S.Q�8<��oQt�Fo���[�B�)U\��1����g7?��������0�����*M)��P�*�2�ΰ^���}�}�$���g���9$X�cV�rw�	�-����GQ}�b#���S���F�q=��tCpTLS�T��p�[�����X��bP��� ٢���j`���,?"��>��ƍ����_���gej�砝,Z��9'
l�M�<�}�W��>jf��T���'FBuh2t_LƼ�߀6��k��H �����f���"�4�l��b�E�F/Y<Џv��)N�0e9d�ʟT1;78S�P�+�K�$�����[�)�E.����F~J��G����𩼛�u�2���>��N��-0)C�j��M#0H,�|y�{)z5pН��%̼x��z��F�0�e)�& �ĭ|:�+� �(�誔���F����z� d�(^�	���'O���d#�O&��ZmXZ3�ӂ����E7��:����X"�|�X�f�V�D��M��5��-
fa�Ӿ�~$�������,�@2n$�����$ekd���p�Xȟh���Ik��]�����j� 7×<FK���4)&�!&>���9@�_Z�p����m�	�z�h��e��28�ӑʍ�<��E�X�m��<_���]6�|`���ߢ8�C�0Wa�22�-7�t1l/A^��O\�פV��6\q_u��g4Z����g벺�h4�u��_��K��U)&AY��Su/�r�l��ӰH�_Z�-E�Mw��Ht
��ڶ�Zs�$���'�}�jU�r
^�\/���XM��c0ka$�t��f!��P� ]��x��wژM�2�j����'*}Y�ж�8����,m؊������3LFq��a�jE�~�VǏH����o@8��щ7>u�V[��% ��DWj_i[���/�^W�?��c��$�t۸�Vf��4�j��p
�r�3[�d�*r�Q́��#|%N'̠ƔF5�X��r���f7�b���l�I��`^)}n^�E��&`�"	<��ҹ�
�6h֫�e0L�� 43���"�r��Xu��4�f��g��x���SF�P-W�g�Cl�XA����p�#�F`",��_���ǔp��X����'�{�F3�@���HJ�Ee�e�-��
�T�WcJ="�x�Fxj?�Q�/n�����s�/#r�����/,�章="R�A�F}�X���T=c�g���#���9����ԭ�.�Og��WPoܐ�*�!7��uP�P��j#�铿��!U�t�k�W�A���tْ�;{�L&��;�{S�C��'��Ks5|���z��(R�.��+X�/��4��\N50W��7XJ\ݿ���n�����v�|���=C��_�<�� $���%��wɪ;r�XX�����	m�>
���o���ԁJ�����a���Z�.�`��ڃ`4���:bضT�1���|���C�n�xZ^`F[�*�^u��짾�r�9ZS�6{YG����<w�q�8y��9�;͈�8�~>i��O�?e|�e�>h=��� �p2
p����i�^A����U���{�!DoPEp�몳79;.��^ݗK5�RN����zd5ke�$I��qn5.gK�n±q���V*�j3S�`�ˠ��j`�j��S=EOr���<,��Y��[].d�F'����_��]5n��R;m������t�KoG�����&���(c�e(�+�B9�]X4�O N���_"|O�����u�7�P����4�vn�����<��Ф�IQ���xw��+�>���`���TW;�K�6#�0[�f�f��
\3�֕�p%F%]z����e��ޟG�z�e�e�ǧD�Z5ym$cg!�nf���Poe�~uwf���ؚc>�1Ȩ�8�=�(m������(W�qzNnnoS�N��G�|WO��|	���%8���N�w�`^�'��D�+�˒��x��HW���������R(L�<i�=�BI(�����e�\���D��C�t����um˙�8���Ք�/`��<����
~4h���A���.��{���玦����z�,�����tM�?�%[�Ztc�[:��Q�R�kyU������ ��� +PE[*ޛʁ�};�\�����ŕ��	}P�#�vo�G�����BB^E��ƪ�l҉:�c������7\��u}�$~�������h�{��5�1��9�6:� ��\�E���q�X��*��Iж��4�Qk>r��y�+PS�H=[r��/���B�ұ�}�0:�R�|�]�];����DpN���7$cMj"�/��bZ!�Y�u}����<DD_~[Y�'m��<�׏v����4��O�`\<����
�7�N�Ѡ8t+us�B����U�N���[��>�GAD�i�ε�y�n�AV
:�u�m��!ϓ8����[ک���w���ٲ��
D�E�ɕu�w���f���#J۬��\��&�ر�hw���ӝ����q�[<P��Z��Bx��4��X�~^\��q36H���u`�N�i��owE`�r�{Ô�ck��\��<C$!� i���F`��v6��S=����F��C{ �Mv�c��&&��"+��h��
Ya0��Kj�A�Y�S�^�x)NY�7KHH�:��.	%��\�����φ�H#)j;�דLӎ[ue ��Q�e@���|1�!|���m]`��k�Bmv6�q�W:����zF��r��lI��NF��*��G�t}GA5�f�7xk
���DO��mS�t������K��
� :�0hx݉_��S9=���d�W��(JW;,vC&����`�`[�]�'ϤA�aC�&D�/>H�Bd�q�'%'!����S%f)�\��'��[en2���-��ma��E�(����T�.������l0j�TL�[�x��������$FxŇ7��\ٔ��c`(!�dY��䬡���s*�f࢑�C+&���^�b9��t��/�&˵�#��⍰���2�|��7x<h�n��s6S�V�`��"�X���]�1GF�c�|���n<ܒ�d<l�|Н1��S5"�Ml�� ;����1|�2�C�f6ko�+�Z��/~?i�o.�%670�!�l=��T�F���m�H1��J��E�b8�Q��w��5꡽.������઎n����n'u`���8_t�t�gyo�xu�S=��W�r d���)��	��x?�s�����FQ�y�%/�i"����:�쥠k�}?�Y�!�!�o�����G��Mw��d�x�M��)[u�����LI�����289)ёҵ�}���E���u�:^��4�P�y&���KM5;��0:�^bj�U��d?�/#;��Sf(�w3b�,��@~�!�nTu���^�H��O���c��T�/3�� ������v-�,����p D_~+ c��-�׻cU�s���H[�@ -��,e�\C�����*���; >k����2�؇�D�W[uZL��M��p������
e0Da�уJ�/p�9��z�)��	�Q�^��U^'!�b�O\�5�<�!'-Y�
��һGi�n�gu��d�~e��/�FfXz�W%���ͮ�;�C̈�'��09��_V��~|�{<j�T�"��Ћ>V��'�k�5�O�u �Y~OO!�7<�����W�{�[/R�ق������(����	7�!{c���jFN�p�F�{)ث��_�������J�̅E��_Z���}�X��$4]�r��Ġ��C���W���#(�~� "_�%���8@�c#����zn��D+>�%�w��>��[{���TӇ��B΁����:m���(�"��<@��hy����1���zmg��x����1���O��+p��T�]L��Ԛ��.ȷ��)M8)�/�6�F����k0�pޔ[!�XQ
��j��]���`8�:%��Մ����կ�JӝO�h
�J#�[腱���oo���E��XU!B	#��Y�K�s�l�J?2u줚�}9�<����oO����f�҉�@s}����M��!�dcC�C�����g3�8�4`��U�>��'�a �HP�/���Ub�˴���zE����`M���2$�%�k���� 'K褼��N/4+��Lz,����u_�N�����ǉ�(��h!�Rm��4�+b/5$��)��2.�Oc'(F��L;��'�\Id_C5X	�[Q����c������J�ƒg�,����iX����e���	C�9|zO�u}����~�J��j:˯#�����-�*�;f5�Np�:� %F��̘F�5dg�R�8�G�_�c杅�@�!{�Y�령 �:����_}qN�.�싴1<��B��Mnଯ�;�5�i��5���@.&��BO)qD^��c2��t��J���1˨/񚷻��9�l�����O�M���	�/�Rږ����p�֒Ю�M�H����u�#Fi��կ�"����'�����t�nG�7+�2���U�~�'�
#u���g��=HQ�jAB���T�T���规��c��
J�k$�W��D�_Rܕ�����R�o'�@!7��x�xh(%�M�3�0|�J���7�Q�XG�[�z}�h��Ro��1#+��Y��&�bb�繥C�R���ݬ���@
����f?;�<(� ��浂\��@mp�܂�]R�����T$��T�!�ً���g�-c�5C�t�OM]w� �hD�w��~8�g��zުr~�����dV�*i%p
����z/>�X��'E�Fo_��;P�I� ��ibl}!7@�GC.�"��	�N4uً����F��" l�+�􃵏��!J�?����p�)�F����B�˾s��i�ӎ�ʌ�"��|�N��9Eqb@�މ0��	Yhx%�9��`�m?�L��b��V�	 �as���X�M7C-W�2�S��警3pk����=x��m2ư��A��d�p�*u�7\~��������3�4+��/� &�_�a/�Rt�@f`H`�H�C!��lSu9�h�$����_Ȱ$�2�	uV*@� ~��4���V]B���=Oߺod����)}�Q[�@��?�>��V?2Cc"I%[�6�ۄuS���M����Sdm���w� `�ۻ2�o�X:*Qh���M�|���`�n���F5�f�����D��	-�M���"_Hc�[�	�:@�����p��OD�&�y=N��dr��{�868�X��r��s�	��<Z��#�d�k�/�M
��L`�4�@ż�n��	�4�,�!��;�D��e݅��P��e���/Û�)V9����x֔Z�}9AV<0�jk�qS_��e����|��i�2>��|�¼�:�����<��}�Z� ��2�y���=�sɏ",7^��/����?c�Owo&����3|��m�֛(:-M�]dU�=F�pX|�qQL)+������L&ȍ��-�p��^����~%6�3��Л���	�Wq�gB5��
&�7צ�̦��or�����>�"RCi(u�tΝ2�Y���:�A�8߷e��� �p��FOU�1աg͂d-����u�A/�#�vZW䍍�L���N8�K�VڄB���h�_��[�㉯m�I��mBn���b�jٲ*r����P&�7�'�ǔ4�ω�?�3�8��8(?:��5��6�i}�KmN�恚��)/�׻K|�u;���K��qsA�T+�_d��X�J�)E!��#n+���������8�%�sF	r/��(��
���|���N/A�?�'!,��*2�D��g9>Uc��h|���:.��u�!a�Ys����yG������s�j�;���PQ0�b\扮�'��0A9��T]՚�ϑ�b��6�ǰ'�`����z]��ի5�VЃ���߿���.]"��_�L��G������L�J�F,���RW_%v/�^w.�x~��k�$�+��5遫I�T�}�֢^<ML�O`��<���3��cG�,身H��<��s8_�<�E/�W fځ���p��}_M�qϜ��v���a��F�k6��1c�84w�'֫[HKv�m�K�н���?���9�-�s� �of�l���7 v{2�v�^ N��)�b4��U��x�d14�	�u��E-�u��bҺ��ɴ�^��;��}F�}�]uB{�Φg�퐲g;��܆��r�W�m���";�I@w��5���b;��3�M�1�F]�����I����'�Η��?ve��P������}�,˴5�0�������)��XC�Cp+�fr�M�`����}�&k!����Df~�H�n���-įg�ƫ�&���l���ed��D��h�˨ݫ�ȞM�x�x$}UF�NI�b�Qie�\�_�?
{�e�TZJ�i��R��lm���R�,�c��p�0�Z ��G�C�ȧV@s"b2b���<
��ck�qE�6���2Ik"lBv����A>�emG-�n4^����_�%��3U���|�,����%���)��I����=a2=2��+��=�������e�(uX���XN	��━9�����f��"<L�:[ܠ��#��(����sᧆ���(�7�x��gEw�{�f#!�IF��1�ɤ��	��E3*�-�-���!� RƔs��@FE��e��io��:>HX�8v��Z�j�z�i�bэ�oh�x]�n���9ς�%q�7�@s�5�B;y���	��%�P����$/�NQ�����!�Z	�伯,z���
�`0xꢭ7fT�HCo�P�3}��v_�9"F��UsC����ؙ������ʙG�V"��R�׫�y��bӄ{�v#)f��D�_wZc1^2��F7�$
����}a�x?,Z=��d!�_�h������(g�/���<�&�b-��U�Zt#�����h��)�\�R��ͺ�xi�~V�+���D�p����Fz�����^�u�.�"�isl8���)y�1�W��`}�G'��j�h�Y�?��٪�	�emt�HG���7�HR��(��a���
��\���;�Ys�W>t�r/*4ZJ�HC*�ahV�+#X�u2Tc��{5�`��^�c���$K���Bq	�\6C�Y�]�+
�5z�)�W�_0�lz�<��� �r�� }���~啖�.�m�u��+ƭ�K�	DΟʴB�@A��;����}?�E,ؙR����?\���y��Za�Wi.�~�d�����@wm>LJ5^������w��p��~h9�~ax!�ӔJ�E:6ǝ���%��@jV�Rɿ����g�g���w��|0��8X���
OBQJ���������}�
�V!�&ۙ�0U�B-`�aCs�ґ~�)����V�lE,��IJ�[Ş����ː�D�(�ތ�Nk76В��3�k�x��Q%��$`�A��g�1�m߻�������z�V����z�֢��� ����yo�6��>R�{e[�^	���6�����WH�Y$�7o�K�������ڗ�<��>�Y�b���NTRfi�!���K]���O,�s�dp`��/)#0��ݑ��U���q\Ph]���ărz�N�-R�!ٕT�������xe����H�ѡ�Aj� K��R}���O[�%Ĝ%	I��7ځ(�3e�x,- +��Ǳ)s%��0���Jrե�M� =o1L���S���*��.�nm�Aퟄ�Í��=h���K�����������+5��0��۱z��L!��.:�E�����L�D�V@���{s�)�Lοt���U�Th	���p��X�l��ec0(�)��Sb�zkğh��;���d�_��.��+D6?���t��I��ȴ�S�R��NKܩ������jp�&�e�����:L��C�|�p���L�����1�����s�q�R0+��E�"����
Y�5�٩^�i���b�w>�Y��b�q�q��8����^ZW��*~hA��{j�u�IL�ե��9���S)"%���i���vaoYpb�v˕��o���x����a�*�e�纯�CrL�;wJX/H�������	����AgdQbn�'7�Y|�*��~ތY4
e�a��1Y�� Ղ�Oډ-�(�7ڂXXB`�,��p���9B��kn��� Kr�lX�i����q���_TO�Fq���kr-.{s�WEAv�����t�q� PF)J�źE��c��LBR� �,����C�C�3��C�.��(�~CX칟2�U\�������H�7�`�뀐�<��v.J��W�t��8���� B
��~��ch<�8�nT-�>^!<�k�O?Iރ��a�fQ@gmyP��`�r�#�G��Cme�#^n/�����j��)�$d�)i����c^���~��P�$X�@i �pSyw>H\�P�E��	�!�}�'�rF��V����S�/�*��l#4̕aay��$�$�T���a����QpF�=ݧ���ʠsns���?�L��V�SL�A�W�5�{�����Ǖ`_�G5��)	�ͮ��]�z�U����Ϝv3@�(�R3`��J�����v��b�d4�ۮ��6x1�� c\M׃j�@8�hQ���T�_*fI'�Lʩ�H'�@!-�$���Vx���j���p�����9����?B8�7�/���)���Zg�?>1,���p#٧_�ˣr���O: 	Xe.8�N\�y�P�qH�ף#�6�L�c�]xiXlU'�}�Ds�A�,hP�@|໴�t��1	TϸE� J��x=�fg�V"c�ļ]�g9Z� ���W{�^����h�2�\Ʌ,��\����ޭ�C�X�s���1Z��6_J�"�t ��<2M��20�u0:��Y����ZY����r��ف���k�xUmsTV�f2½8E�:ؗ��
a�Hjd<��B�"�o&,����~i��\�/p��Hb��s~�é%��$D }�~������F^AR����PdI �`5��ϧl�KI�?l.-[zK�Ͼ����5���3_5hsإt�+��J6�{R����&A1(�1�|><�V*_��i�i��ĺ<3���uO�
�#!�ٳp8x ��͘�r,��w��W�ՠ��X�x����`j �jV�5yS��UѦ���a�kw_���e�p�W�-k��(��Al�������p]��(��U��\&4+�XE%^��,�E	�I��I�~�]�"��v���0RZs��F�ϛ������5� aq%��NnF��"3�� $?���w��P`��K��Fߜ%��My�ݛ�p��ic	��}�ZT��QY��&����^�4g�@�+ijI�h��
���Њ���.��4��lPyw��ZJ����ʙ�`*l�ۙL�S�k�o��;j4G��جc��Ϧ�����M}�������f�񳮧I��dq��I�V���c����\m��f����c�U�o�b'%�q�'s"Vb��e"������m�tOR��,�m���H�S���1#K<Ri�PN<eW'ƞ���"���ЩAJ���HF�\w��n�}���R��m�㝶1�1�f�酼�s	�}k��Y�cc �(G�
�|Edrp���H·j�o�ŧ��9�:�`�5���1|����A>DЀ@N�ĭ��|�!���X� �R �CG�m��7u��=#�h���.�S�.�x���0���{�?����	-'�j������.��8[j騮;֚R�|��az~6���L[�Ct����r X�w8�q�D�������C8�j������� �k��d5�3�t�Կ_q�&���{yM�fj�lv?�ɕ�h��|���}+�-���n��j�l�ؠ�X!��`�K�K���:�n��=�y*<�����~l;8�IrT�
��$�nx+�6ݸ��~����o�l��.�we�~
	zs-�o��0A�٧
s`i�Ëy
�
ޠ�"^,X �a-�,����Vf�8��&/���_��ql��ц� j0���HM�ȯYm:�ҷ�Z�W-H��Vts��9ԟtWY�YXM�a}x�, _i����G��
c-�����N���q�0���i��ﾇu8���r�肣L�u�<�жv-Ɣz1�>�� ��57L~g�M�b����|�\\T&q���8P��Kb��[\�!5�zd��)-����P��{C�K�=�̾q��`;�� �	:���ݚ1��Ts��n(��1��hI�����i�3�+n���jUcC/�A��fm��~!I��lL`yp�U��̀�^$>�b�?4^i㒖ɠ� Wt�����JN����*���.�a�Z~�6�T9s����طGB匕�߫4��)E�q,��^��pǘ"QoC�����0#�<\��e�\̥ ǢR�=�M<�y��;�R�~++���?�-�(���=l[9��֌v��������W�%8bo�����@��t0&�y���c,��BBʰX���Ӥ�xT�m9�ߠ����'p��*��*
lH�0��@���{P��<$|e��N~���4������U����4�*28=N� O#<8"<��*_��R�X4ԋs�1�����@*�u���W��J�b�K��؛����V��-���e���L��B"�K��}��4�L=N%��BX+D���i�ۍl�m���)w#�	k,L��"|h>�E�4d�|:6<2Ij�cA�YG��^'�sM��Ț��q�hF�����>��+��'GE)�)��L�O�!Av4/o�IP���lkXbrMK@�A��Y|�OE���'�?�fָ����k��b8�����DS{0\�O���Lo�b��ދ�+�$����d0��r��(2l~�l7�������3��7��o���f3gCykb�.μ;7�?��Eo�S$�UA^��2[�:YH� ;Z�$f�h���6��oFy��D��q�����wR�M:eV��+���^����.�r:^̚Ns��`�ԟ�(��MR�-�ݍ����p4ǢDC�Y��)ꊚ�̡:XL����Do��:Q+��뒤N��+���eqA�9~�>���m��SY��A�Ꝯ4���}}�L5�r�]�L�1�o`�{�`%��s����EF�1a͜BP��m!�;�l�I$0�m�2fb��r�K�^B1��-1���VZץbB�X���x�4`-��[��V�Yg�?2NĔ�w�6{Wѣ��f��Ǌ���SQr��w���c�.�׿���_�%���4$�Q�lehK�]d��$�ĄX�W�n��}^�,c/�����VA����ԉ �1:y.��X��-:��+�.�D!����
c4�\�L�`Q�w��O��v}БQ`,$���S>ui{���q���<NzR3c��6���_�2w5�;�M�.��E
��"���wx�RI۲Q[ D�ai
$
e�2}���D�;*��n���'j�0�M�G�zt��������2~f��o*X���̆يKZ��FK4� ��!n$�K���ꖇ`\F�M�$�
�E���w�[oN�N��$���9Z�!Λ[9���|tR9RY������s����-a�O��s�b.) r�_M��&HzK�I�'�M)�*�r_Hi��Q�t钕|�nX�~@�}8:|�N-`b�v��'j|*ݟcӠ�y'_�7�Ѱ���(�׻�y���҅[B�6��h��=q��s�P�ðx#�3��p�m|&�.|5�g�2��2~40��p	�^��8�<x�� =�ـ��!�9�?����ӊ1��Y�a}B�,��Ō��,��Y�E�$�W���P�P��jj��b�!+\�d����j�f��U."K�zA@/MN�,1��/�ä��s�Mw\ԯ"Wt���nh'z?&��b�hh£<���v��
m����L�A,��s,h���PL�\nT~�;>V��<�xu��PI1�5�tE)�J� ����A��6�?QF�c��PR U+e�%G?�/(Fi�`d�u2�w���45�I�k`������=��(~-9�Z��c;��-�v������7Ye`���b����n%;�"xI�
�����\G���N3Fž�n:]� �����WI���zL�*�4b�D��������o��1�����ǝA:>��H­?�מ�	�E"��qeP� Sj�]�7R�x��b�Y��!���
�h�b�Or���𥦝A�4�3>��m�@P�<���b��}�p��p��Kr�Q�i��[zg ~�ϴ	«Tr�!�}�H��y��:� Pջ_�͘W�뭧�}1�H
�#�:ak��s\��������S��2t���j%*�G��ueW�J4��������O��5ֽ�6��K��蒟�3#@��7��3���� ���1��0�۹��G����s���&�"�[�|@)��o=���MZq�Yd:3�f�����Ϧ5�n��H���Ŭ8�����
�ZN跾h���m���;8П��*�"�� �e�
��!�睐|
���wVJp>�hŮ��D�r�5�vsJ���ĭ�D.�Α��	�>��Kq�N��yE�ak�Єg^n_�$[;��:���g���<��n�ı�mCiL�=O���SP��]e�9��u�7S�A���l�A!{���)]�n����i�;�I�]XD��,3

GC��	ƺw�� �k�^�0F��xdv���;;e���O�ok��{�+|���Ҷ�G�p٪��,��6٧���k���ύ��H ��@R�O`�TrL*���v�W�� g�k��p��D�E(���:r�����j����#�[H?s�W�S�u6�=��*+�I�����ѯr{�����G�v��dr��������嫋�;��Y��[^�Qv3n[���A��*�xf! >���y�o��&����%�~0g�AT��b��v����l
	�#/Hs�o����fH��l���Ӭ��.{�cw��oo�3swC?�%�����Hֿ��-��w27 �hg7�(Ӕ���H��3b��^������=�Mi_��i*��� t��� �� �[;��a]��r���|�7S������OߴL����ޜy��t��1CEA�t��ؽ��%��!50�
!���z�V����<�����\�2��l ^��xS<p�DPNk�'7]��]���7�h�1�K�����x�����>��4ҭo�sJ�.�9�"|I�_y�g dmr���]����՚�����k9c"�2�Q�j`[��kZM/r�-J{ܝԤ��w��S[�qj�����Ŋ`�^�s�w�O4�,C�B��pv���8�0Ǭ��gw\�A��IT�u��9����̺WU�b�����,U��z�dy�CMy���R_�{Ƀ<U~n�/�������[�m�Ԩ���2P��z�F,�e��S�
�v9�%~�Z�a�&�3ϸ~���"��!
���<2�K"ؗ�Z.h �qe�(�\\�U���t]�q*�tw��4 ��?��6p| �aU���Wũ��w�|��[��ysyqjQ![�&���� �-|���~��Q�oW�­�R��e��M�rex����2�B+�c�LF?���F<���=H!���^���3�P�8u� ,�X�j+�C[5sP$�Og[I��9�$�c
������sM���͡8u�ǧG�䑍��~���>��y�żu�h�V����H	]ۉ����7�k���ѝ��ʾXL���VT���"�?�8*[ C%!�$�J�7�-d�9�ԁ��N��%��O�-=�fQ�P��~
����Nv���r	и�����t	�ॊ����������K =S��r��;?����n��ǖt��Nq�%z+��m*����L:�t�T��B�N2�1�K��L��G�ț.�=tM$L�|B��|e�'�����V��/���� �v�@8�c5/��0H�h��c� ��	r�w���^�"�����C��ԟC�Na_��y��=[C'��#���z�y�A~��Aʇ�*B=`�ا<�!��q,���7�9;�,0�~zʼ�)ka���'�<�:$�c��C���UV'S9�|��5����+2+Q�1q,�	������. ���X�E������[�[��.�|L�ܼ+?w�ڛ���9mI��[���Ő��.<����!/ ��l��ܰR4�^"�~@��zJY�3#�M��D��Kg�|K�����w.a���X$������[���^*�Hn���xS�T��f��m�,@��켮�uL��Th\=�R�A�r�o~ 3���nO�"D�-�0�+��V"���;�  ��Kc^+��*0M��/^K�Р���� ��Mԗ�[�����;0M4>`�+"_����ZL�%����6f���u΄ͩYe�������KCt�FE�r-�؅]���&�}�3��N;p}���*�M�"������+�mI:J:�v(��� }m�<d?B�Q���=��٘�t�r�P�$��1Tĳ�,Ē����[S��+N�]�����"-�I���d���LW����\���~$ѕi��yk��T}�v�R��W�4V��G�o�V$s9�+}pN�I�s��!�O���)߄"��_�\�%D4|�4D�����$!%@$!�����B�P?u���W�<�_Y-��oߪ�hԑ�@?45*���C�P�e"z�����p���c�;�S�V��,�$�ƑY����[���ş���urF��X��tv���<���p��+��?hC�.�춷{�a�x;��Gv�B�t]��u�:��jw��S�#N��z�����~_�"g�Y����쾧&E}�Q���Y�)��|N8��W��{;m-;�
>p�ܣ�>I��8LJF_�d}��s���@~�b��s�1NE;~|-떭���x����a{�r�{M�Z4tK%��)]7���߀z�ٔ�� ����`��m._�������;��(��X���������=CV��`>�@u�k�72ؚ��*�DMl�$>F�IOks��Q(��K��#c��h�?����J�ƫ�
)�{�/����Z�2��"3D����U�Q<G$hT�-���^��b4fĽ��\ ��P�þ��r@��M��-1���th����i��W��^��蕣HNyA��2��W����F�9�Y쇑����5*;pf�9�0/�.HHx\q��WY#v��]��o�mHѾ�ض`ten�7��qCl������WR��{���a�Qh��|�:�\��ú�ד�$������V,��HC��#�vMh��$�S�޼M
k-����Q�s�g%1nB��ǅ�0rW��][7��M���q�m0��%�z'lʛ9�#:G:[x�e�;�MX�}���*+���iܖT��և#���A]�N�n�m��_�if����P"�	s@�)9���G�a^$�a�x)���w�h-Щ��{�ă/�"Oh�-q;4���i*�3����(�Dcs	�����[M�*�!d����=��i՗_�DO�B�-��19f���[�oNE�[b2Gq���"m���\ѯ�Fd�a�f���a��?$�%SFd��j�W���,�L�m��Q�V��y�����_�ӬS�����_��cΐ5�ϴݲ-�+p���jbj�&���z�pg4��fV��|p$��ޡ���S���(m�߈�}J��<rE����1e�}v�����sLN^i!{�>�XF�%��iKV?+�.�R��R�.���>���2at[�/��M�m�sN����c��yP��`e�¡��`)�p���okcH2��tl��Ӓ����@�&�2i	�d�����|"����.�5�a�n���J :-����28���R��<��Ze�νV������&� L'�}b���+�y�Fu[�܈����	�Tp��Q)�oup+�*x)��aQ���+�4n�M�{gAo5J��E��-�Uw�h�o :$�����j	�%d�5c�d�NS3��4^��E�>�	=7��OQ�ε&�� �5��Pt�&Ҧ��Mw,�V6�����פ�Ojl�FOJR�CI��)��&J/{a~;�p{�x�����Ί'���uU���q���A�T����͟�nz�s�`�^�qP�v�Z�yt����~A��&����䋺��,�`�n��
����;��_�{c#���~u
j�r�̓{R�H���c�� h�� ��O7�Ӷ��z�,cM������iz�D�&�9@;L'B����I���3EUL(T�Y�8�s�7�K�k�s��|V����%˹�Qg��C����G�꫌��Q�D���L�6ڜ �r��v�,c^η�#l�؟crn�to�{�*��J�̳����4lnNI%a�|ˇ�(����7X�p
>��a���]v�4Q�&Hy捜-�~h��56�wksԢZ�����!5# >����u��m�����p&�:;�>dziU�%>SU0��.\��Y��(0Sv��c{33+�@�����}�SS�t�?R���4�����Ayj���>��74���Z�U�ďv�����<|�c_�K�$����R�Z��Q߷�C�6���x�M-��{��P�R�� #�D��`*�D_��������������^���>+Q���LC���b�U�"R�n�@�eH�����l���j�?�b�����{��඿!��H��/p�[w�ߋ!d�SN���-@��b3���\v��A���O�?r�t� �ē:�U�*>��w7K�����*U�(δ�*N�>��#͸~�2��qH�@�Ȗ�[�Kq�k�1G\#��}�xLA)F��m����#E�q��h噬'.Q>~�J��_���u̞�D�@��-Z�J�zA�6��ÔR�IqK��d��c�-ڭ�dOl5�,�*�{%	�8�Nύ5ߤ0�:]��ԓ�� y�.Z�j	S E=�n�]%���,���|� ��`�"�{�7�b��ѩ�Nb�B4�O��٧Px�f]��G��ހ��Q4��� �	>�n���n�^b�Ԯ����r��]-��v����9��6Qw���:e���
!)G@���|�-2�?�i0��'�p�ZP-�s�CQZ�@z��&E�_�1
���Y��N��ub9�%|	�0h_EP�T�,[�$�{h�Ϣq�N�bB;�ň'I9��8+&$H���?�C�_q��<Yj������S���:��
*ӡ�x���#
{��g�;�nmm�S=��6A5;��r�Kon�t�w_��%&��<�//��n��`'a��nr�5�c���T�Ǩ�ɖ��
�p��/Ot(���k�U�w��f����kIȑǄ%� ���C��6�2>ja�˸�@���uLBl�5��ژ��l&#�4��?2�`�Ϊ��+�\�����dra�i:��(VN��;�rSZ�,sOL7������<)��#�4�[ ��[�^v�4���i�Ďn�3�KX� �&��zZ�D�b�5�EF�(w�>�m\�Z ���P���﫲fSB~�N궏��5y-�A.S���m����<*HH7�����EeG	g;*�6KơgѸ��ʚY����79��p�!� s�&��	��d��]���}�����ܣw�7�['Ϯ�0�8=�c�igI�3�V��.���ĆC�bO���<�����%�����<#!Z[`��$Q���΀�qݟ6j(LÕe�e'������"  �,�0��q��{J��R��_|�┛�B��T�A��MCx���ԥM��osc�^gB2����b�-���&/���9��ȒZ#vñ�d��=��Q	k4lš!I����L<�Y�h����Ǭ�b[��퉾���u�<� K����G>�fM� !��S�[���&|�� �R�=��X�z�!
kH]/��Շ�Nm�ȧ�aom�M"w�x�k���=����Lt����hZ��}�S��q9�z�'��<�q�A�`�e��)��_��\�|�9������k�Q��1��z��$�V���N�9����x.Q
�_�k7W(%�w@Q7y46!XS�W%Z����)���O���ܺo٦}DX�p�|��-��y'>.'(k�m[/y[�@�[�[EOMs	ʊ5�s� 8ݾ�~���/�h͘�B}P�V�S�d.Z?��h�o���1&�G��σ��2��)�������|����iFC�C���۳+m��h�-��)�8�JE�g��+%BR�O��yu���b���מ��o�C�b��oPtkݼ��-  Y�K�3���E�j���Z�3IQrú�w�f:���F������ʖ��@�<����V[�pI����@ |!�Y=w6PZ~oKK}��ٟ���I`��B�3XC5ւM�ޯ�����&`�{�R:^���	K?�,����N�Q��� h��(�XS�_H�#�$�%#* z���k��t;2�����?��^�\�_�c���\�e~�������-���P�zN�oh���7D���צ�7�tSD�~�F�K���t�=���K�Sپ�n۰�`�="Q�s��s;���� �ݸu< ��Z|���(�<�v����S?X-uXW����6��ϓ'�p+��߮�	ތqa�sqa��$�P,W`2bB&��^(`~/�Uu4�|��@O�P|�l�]8�N���j0��?��<�y�%s�p�v�ZEsCz`tv� #3����CDƱ������eR3y]�&>t�_v�CkpK>ĺ_mȤ���Y��K�ٞ�(�E,n����Y�����W8�Z����Z7�&����Ҩ'ċ�hħ�c�k=|o;$XEsw���!k��ڥ.o���`��iӈ���M^-��YL���)��2�|�(��iloB�y�Q���8L)U�bd1Sʌ�n�l�qѧ�p�>S����4oa�ؖ<E�����r��>�Y�K��i�%=t���Yц-��1�ys����D��M���u�����<t�ѕ0\�r��^��fH]�K�Lؖb�p��øu��.�Z��Y��?�à}j �v��y��Z-?�n�xQʎ����&��
ɮ�����-p�'?�U�9oc��ˡ�VB���W���b4j����=�m��*�r g��l����;aY���e��CKޣ�}�����?f4��enXO;f�-�I��n'���Ä��̕�a�����]V�2��!n�n[��,�kAq�V�K�[���-��Ne��w��4�?g��Z�[���0�P�I�Nc �Y�U��AT{s��Y�9��5���+��My{/�HE���@K��3񻟬 �zǻn�/�~��O�0�֟���,�W�pp�[�VP�=4g�LA��g��bs�'.&���x~������0�c1h�����ϐ-��/�\?�Ղ��4�aY1�r�s��%����{]�c�ЇlQ"f|�ݍ��=|$�	)5e���?�-�b��wMX�6�����߫
� �
��`��c�����3�(oP&��/��1L9>u�|`��ZB������� �(���i��S��3�TW����:�>�!o��|~g�<-�����<�� �����0���t�S�u���|�r�W��P��G��U@�c��GA�X�#J�}�j2u��A"��/MN҃�G%jq�U�����T�w܌
M���Z��v����r�6�䟕~�4\��?~�c}`y�W!�^�5�Q���:_H�2���9�bf��r�FQWY�:�+�����`�54+�����6���`��/��[�[��3Y���O������KHtVE��~?�/[lY�!�	��B��]�(��RkD�0L�{�
Ղ#>�h�3P����"LE�QNK�P%��1��F���BGd�x�N7�t��B�_귳�0ZU��ֳn��AVFl�x4w2�.�����-�a�0���+�[i�O�Y(zd��-
ERGh��횒\ �w! ����E��0!�S���R"�l<�o<�����U��ٌ F�"�����g�Q��#(�c�1o�P@>�Г��!8ճ����@(���PHu��{T�Q	�­\�2#�C��84�x�o��o����ρ�j���ec;��ޏp�M�d�Wtj K��ͮV}��X��*���!��.a5��(��>ֈ�j����MI�qdM��.i�j�w���nvh��R�ڤ�A��Ϻ5�g!�����gR�mj��R���ܮ7���!;�r�B^���������|�0+�$����F�Y�&]����9i�Q`~�#����{6��K�PkJ�Ng>7�#> s#| a����Z5�f���U�5y+/ dm�2V���D�"/�W����Zt�/�&�@u(J�,����C���p���Ê��9i譞e-�9�RX����O1�3�P>���� /��T�$�L�U�.��зm�S�:�ǆ�9��J
?�a�T���d�(.'e��?�j���� o�oZ�����0��,�PR �Z��$�<-*��G�2M�I,��������wFx�`@ɳzϵu�d�H82NAt4N>,�dAR��;�B�P|�H�D� sT&]uH6�w�x�z!1��;p���ف�kb���m�ۖw W��'�2ɂv��¶[�~�������~��D�N�_ ��H���ͮ��Uy��#,n⋴x���l��7!?�#Q���!A��؛�)L:��JJ�
��2���+���f��^7�������}\I�'�ܙt$�AkH*�t��Ӎ+�wI��Rzl������]qNї�d�,%M�n�RU�I�C���;��l[�Z7�!�.Z%Yl!st3����?���W��>������<7JĨ�hb�}+Q"з���	 �58l�����$w����Tй�uL�%�̀�π�߃bwh�����E)�Â���?l )�l�]oBa�ݖL��te��rn�f!q�M��n)`G�|�=7m��C���@7hq{���Kp(E�P��鶏��&ϯ��L�a�u�.q/í5��y��Z)�Q����*c}=j�&͊��fH���6�-a�T�˾ܔr{[l?l��Z@�V��re�.OH.{ą���_���q�_��� %p:�}F�Ԯn:�y�1|��0w�T��]z����9齪��ٷ�k���bhSd"��o_�$!���"��VRlR4�0P\O˯q��(�� ;.Phb�ܷb�v�
�E*�_-O��R��أ�20r��#��(N�ĸ�+���q��o����_>�$��p*0�D����ѷ�y�o]�1Q>��c�e=��ۘ��0#�j��j�}~TV�Ͽ .���/� /���j���Ҍ{'׊F/k�
�a*M��S��Pd��lf�4�+d��v�C�'���P�F3)�C=�k�D�����V���ޏ�&j`
���\��V����ZT���]�6��l'-��m���b� �-E+��?WQ��/����Y�0�fW �ݏ֋$�g�א�1�4{^}������w����n$ ,id �w@,f����K���tr�Au�~�ٓO��N�T:�1:_�	����M��j��.~�c�<�h��qt�u�����mT��������ǂ�49�|��MQx�
p��QG�D4�
ADċ#�˭%���$�(���������\ߖ[�4��PZ� '���w��:/D����:-y�"4خq��,��-mN��(�$���c��;���|n��C\�|Kɫ�<���<����2bd�
�v�2-j�T��7�����S��Y�D�ӂ�����\���f�,ސ�0ǲV�۵Gs�����^WW���do��2�� B���6 !�|}V�T�4��x :EAU�qS����у��C�g�����S��bkq�2��U�4����2D4����OG��E�_8�����Z�A[:"{�A�{���W�_�z��o>�2�#BDJ��5DM�[G��!G�	��=���鏢4�L9Һ�Ϛ�t
(:�!�srՁxYP$�2	퍏��q'�Sԧ�	T]�dW�����@ΘY��{�z�NN;��.p�L�C!��0DԈ��5t��*obT�(�P?��J���N�������p�ýː©o��d�wO��;���aO�C�ܗG&8���x�s�.��ep� ��Q��j�,H���[E��ha/�"�&Q�l@9T���k0迥۬֠�Q�\|��?i �74a���V���,=���n-�>���l�[��q���T��Gca��fnrLw|c7�;�o`�,9�s���%��t�
"GXH��`����_�+����r��Ӱ$�r�Mf¸AOW�����^;Μk�M*�!S��A"g�B�i�,�#lS>��d=&�@/�r��zck��)�P�ŋ���M�
uѺ��3^$;�`�����v�l�����
x	���ʹH2��bmŴ�V|M��Ǘ�N;HkoT���܃��	�/r�\����&���������kss��usf�g>9��I-��Wh�,�S�M�cek��i-�E�%�r�$!�!��\�s��$u|��&��2bg�3k`�00�ZOX����ٳU����:�S�n��(�!���e �����I�m�#a���Gh�Yy{Q2�~�9.�p�����,�_�V��>1�����9�J*j<�7��PkO�~dl]��D�� &��N�#zU\�׉Ԓu0[Ҙ���\	��g��<�HP^�\�f�V�A�W�F(�-En[`��i'�>�]q�g@�U�퇾�P^�yh"=�R�rPù����uon�?6�sZ.� �ת�.J�/bvB�����fj=����y�Ďv�f�oJ��G$�-���#�$S�]u�2�GЅ��� Ӈg�^)܉���8�۱�����^Ֆ�O~�T��Mn������>�wTOۆ@��x�0��iT��Ԧ���հ��o��,�҇R���(j�M�%�~���&�;���JY��mS
0��H�	�b����/5����&�t�/u&�o#�E�eo����F�D��U��r?Ԏ���1`+Sn��3��������Fn�&����m����$nǞE��Z��$��.�$��p���s�'i��F����-|u�?�Q0��L΅��D���ϗ�^7�Q ��e�Ja^�6�x�z^�y6�����H�X��������7�A�)��RK�D�����}��*m==I5��r�[o&AC�;\84�kh��������n��jfu�Eq1���Bl;=�/%zV'�4>�D�2��p\�N&-��K�7*�����!�A�߼X�ar�"��q2ry�܃-����0�m�<�l������\�]�%���rc�`��7p� ez۩���[^P+�+`�IA��q��1�Ԍ:E�Ü2o��p^�@�3)�31���Ѡ}U�&ģ��
�i���,M����3�(n�	 �ɏ�~��>/��_0Z&�(��y
���FO����$�.�}�$g#��f�a.qI�Μ��=v	ᦦ���?���X�����U�
S���'���W#^�?'�WMc�M~s�# ��&���\�۶��ܤ��u����_+��m�������'�X�s�C�$]�!�N��&�?e[�b����0{�U�p׈;���׍�Ở��5�n��4v��iԮ�ҷ��ݟ�e��jȬ�u=�9=�lC���%���-P
�tܵ@��nxB<r���VX��~�i�'z�>���-�L�T�E���TFq��ܼU}ށh?0��YORܬ��C�P��tc��W�m�R���Xm� �u�u����,�ޝ>����H�38IK�Ѐ�c�� �w���(����|\B��}�탺)���P�&!����ل�����8>�Wd���"��E�_v��C�i*��&�
�&��Sv(���%��v3���m�!�x�+���T�t�P������̢�ü@k��"�>G��y��T�W�K����A��o8i�7�����.�;c�uU;�<b4ju����ڲ�H���,u�qs.&qZ�ƍ�%���{�/���P�$!�>�w%���F�ʿ�x�ilJ�ܔ��nSuC������� ���J���35�Ѣ,��#:2���hgp@�� g��=��ܙ+꩸R��_~ʌ�b��9/�&z���#j��ۢ����� i�Ű�+�O����0����HHo�n�������~�:��B���6r2e��a$��K��\��T�m��ԋ�L".�F�'؈q�N��\�9�З��Z�4�Q�m��c��Z��p��p�o�4_��i�Or�(0�{ߖz��h'9����U��ڒu��NU
"��4�T���u��|sE����c��%n�ķ��m�Ơ���]��8>�\ ^�e�턺�Ft�.��>e�X��!0t�S�#n.9���p�����Ϛ���l$�+�i�uj�Oh&�(/JeN7?��r����+�2����=c98�ItUX�w=�?�I�?Y~����F�))�c֌f�Pޱ#�y��_�� =Շ���@���:�D���	�ԋb�����5/5z�4�_��x�tt#��8���uڟ`����0^��?�QB�*��?&�>( �9;x��d:x��Ƥ��Á<�4���ɿ�$�I�w5�?��V���������^�I�5�*kIw.<�?��!O���<��=��I�!X)@}�מ�C�lT�D�A@�B�/<vT�"Ȓ�7)W�#��R�[����,UT�,��Gɰꬨ����V�3�ȷl8 �ee�R��p�H3� �g6�CE�+�����A��#(�5��wr�m�a|�y���k���+aV�*1�e��_l��G\����J�X�6
_U��7]���ڎA��0���NE��!�aEz1y�>�^��$b�}�2��?���L�F�3��r����Έ��	A��b�]��Ψ�8�A�el�����(��:���������}j{�gX�<�+R�%�[�
4=����=V��jkT�@)���$����x���8�A��Ȱyy�٬,V�Lqkyϔ�&.��F'��8lghߝ��)R��a]�J��f5Cw]�'N����1Z9�
�Ê�4�v�Zl[�IuD�!�`�=��L��z��#�x3�M-� ^�{�m��;|��� t=:�8	���aIk-1y�p�PD��Ū��e��x�d�a��� |� juB�7���"��x�<���N�
�|>B~Se��\W�Y�zW����p�{��-͍�|&͗w%����w��mi�*�D�R��TkT�����#�q���V1��I5O���O�)��ySEۯ���A��6�T��BQRj�Z�zbE�Iꅤ�>�Z�~��-,�!̖�T��:�~aMF~���ئ���_lH��O^�I9	�Ep�̐T�J��b*	�,(x|u�@�!�p��iۼ��r���_�U��ޔj�<��Fg�*��� �Ē>���Sؔ�C��ݣ��1��SG'л�G�?��o���0��_~:����;H�>�z��*) �D�
)�y�G$6i?;M�D�Ƅ6�̺�s��n��Zl: �����4?��QcR����w��g��ե�����v������,&�a�o�	�+���DV�]�ɖ̛�_&�Z��ʯ�-��;R��'�����*��Je&QX�} �(�Q�n1D�{iH�>�Ke#q���u���7�i�j�N}1�����S��%i>"���0�;�j��EgsT5��·�g�,�<a�:�^D Ǧɑ�����!���5,��Q� Iɔ���7���4$կ��o$��Jc���-1��	xq뒏�*~8�2��zMOO����F�C��ơ����`�HG\T����i9�(��b��8���	>��AGx���C���S�-ܦ�U���N���Y�Dk�D �7Y{�;��f�sF�&w��ZLE��C��v�b]���� _ X�����)����}FkEk¯��	M\��b�s�$�S��zKŶ�u������$?13(�"q��c�Jr��F � ���e1J���h���\�sJ���`���Sذ�l��,DTqta�l�4{8����y5�ā��G�0%5`N�C0T�ܶ*F�R���bK�VC���b�`����:/���o�P��ƲQ��ŞH9�jOF^t{�>.,��y�yDT=?(�k�x1]|XB4�GhS�t]��9D��S�@G�eI|��7�(yb]�?ag���q���f7�{�|g�?���ݬ��R\\c�9�P���n�8��[I���4.'F������2Q��1�бjgT���»z@x�Q�z�8E�F�z^���/�9R��O�"�w�Ͱ������)ݹmjn��I�à��9 k~��}�g��@�sUC�>��6�����i�I���}`���v�=���JP=�U��,�I���!��'�p?l�H���g�Ɖ_]k�2�M���x}��6��py��@�������S-��JnWZx������OO̹�����:�V�o_�)�y�������)|�P�ٶ�`O7�w��#)�ȫm���c4��B\o�b
IX�7a���}�[�]K0�亘29�g>r�?|�q�����Uܯ���	�Fo��JV2M����E{Y9�<�B�[��z䁅�OCҨ9Pd_�}��Ģ���p�>q���;3�{�t�?��U��N���vb>�I����?��神�A�]f�f�)ǳ�+�;��F#1x�� �̑/��Kk�<�~�A4�ް���
��bv��P��]��U@#]����Q�~L��7rI,���Q���y+@�s��zť{��V�s�ʯ�C�<���� t�ě�@���Y��	�*q��;u@Uzz���w|�a�-��MչI(�7��K�#�zZ���a[T�D�%��1#���Ԧk��ܽ�B=�B���S(���Jݥ�
<��*S�o<q��N\��g,�`!���~�֠����=�d�vi�MT�gf���2׬-�BQ6��9�A��H����jA�~5f�{&_&Q9,��W���� ��c�ght,�V�4_�c� :A�%F�\��8�:
��D]��ƿ�]/Ԃ���A�������sZ��i��������k{�.������/:�<G�K�Z}�m�;��N�R�WMV֥*"��Q��I.!��B��+�3�T�>�;�ss��BE��L�|?�Iw��c܏�a+��1}5��	��7"{�G/�D���"�qA!��1�����(6�p��fM�R[#E�n�Oy��`EIop<�_�D�4Ez�����M��Ն��"ݸ��'�疤'љ���Ϭz�6���&w�ߑ�О4=t�ms *����ˍ��K7�J` ��=Oe"�h��^@L���Ua��	t{������*d-� 
c#�׷-M�jj�N������f��O]-]spv��{�5a�d�@�����X+���٠�)x��m6'�/����-`��Ov�~���['����> ��pZ�7s"%3��PG%"Pl9M�!s�ehb\�G�Ww��Cr/b�IB��; "~U�Z}�c�@�Z�C�1̩<w�ٶzD��Ș �*TVe�б8�,��oph���8o����<jY}R�5�X�e��� �jbnbƋ;( �R/��z*\��z�������lC�E��	&�	���p!�Q��}{��?wPS&������!�iB�$���N{��/V�/�`�y;^ �$�`9�$O�k�t��}�Q]t�M�
�^�0�SI����jZq���qF��R����%-A�3M�*�M�Zt&,~��m/��6�������z��\�F}>.��d�P]Ӭ>T}e�9n���AYꤟ��l8M?��g����������y˗�j�����z��,��}��JL˦�k*9�`�0)���j?��w��H��.3x�D7�8p��5F��p)��]
������ȼ�t����<xo�'Ԃ��}P]2lh�`�J
$�����,�P�>�^�%듗�RQ���;�p^����e/\��-e6�\r��U|,/�|=nW���`��FH��<Z��/ɨ|��Ï^�����G���]|��8��5�_`& � m�%Y��F ��W&�X�bо�M�a��]�l"��n�f��6vx2h�ǚ���r����joY�&~���}�
`�ZP4��Y/>��-�Q��)P����h�r܊���?���F��*G�X�Y�����0��c��C��1`��
w?K�v���CK��X�P��R�)���m�̜�R���@%;��vb��D���@��P1�!eP�Δ�y����/�ʹ���c���^sp�W���K��ljQ��P�l��M�8���u�zm�֝T�8������s�
gD�=�1�T��v�����I�32�M�� XVf�/�s=Ϛ�>�ԯzFq�Q�ƿw��^�i���5~�Z�N���e)���X�9�a{�����Ln ���͌ԫ�Zݓ}gm_����p�z�
;-�
ZWV����`���=��X�-B^��oaWw�{ �Fr�������3[e�Q	>�{�޴�M;M��?IH�n�p� �>��䬐��C�'��'����#��cȣ	Tb������[X�j;��M��uB�d ������{N�l���^��{�]��}!�V$B�|[E�i^hZd���<�����ώ��S}�x ΋S��Za/wn&AA�8�S�q��1���w|��*�l��~��;���U�����/��*^�z�$׻��SJp�~��6�#��\�	����V�UE����d�N�Y���vE���8bXJTRh?L/=��C�|��v����\��z�w*��W�)� ��x�=��d�1�I>����I�.ࣰ�P�&eL!{I�	F��આ�[e��+��� Ni�,�����e��'��K��I��kWUz���}�#�>����vc��8I����B�+T���ym���6���f���ٹ��R<����i��TDZ����e�o��[�Y�|�$�2}.�h5�����$����-(�R̓.�ƽ�`{}��6r��U��#�nxDS2�di�%�-Bj����U(Ū�8����6	1��\�hu���1Oͨu�;K����-JI�d�Sۀ�1�\�y�5��-��2�(P�D����bL۸`+���C�*��Xo3c�b{#lw��q�4���X9cr��J�����MJ�$k�W<I���D*��ު"9�E_ �Pf����_������8C���D���d:6�̔6�W ?���0�����)�\��m�+�����`��^5f���_S'	rB��(�wz=�R��ڬ�v����nE;u�����S��>��3�mu����_ew��p�碜������1���,1�>X{Ҭ��H��h�!�}��"�z-�U�/2�N��L�;!�l�ΐ]+I�ύ�R�h�.�s��vZ��
g���R����j4D���������~l��ތs�<B�gW�>�FT?��	T��?�#_^��_��,�DN.|�f�$<���3��D'��B�NѾD{�~�+�Z<��Q:c��$�3��9T�NW64����ٲ��E�_l�l<H�=��켬�;�u��2)a����\.�Zq��j}�#�Z�W ˉ �['$�\PpwK╆�+�� ��G��E� ��¨{.��H��X���\�x8�7P��كW��S��c�q!��d���NL�G��F8 �S.�甐QOK���L?
~֣�������� S
��eP�A��J�C�=Ej����IU�Gw �P�{U�ؙT2jm��d����jR22�y�3�bP���Q�&�W�V�ާ�I�(4��=���P}������5�u�~ۙ�Ҍv����nY��=?�	�!���_$��e���:؏DYMc�y��@l0����xIGj���rP����;} �1��a�Jm��(^�[HffT�y��u�[>khEW�o!mgaD��āvX���7����o:G�vKϦZ,��XM�YEVкgR8�J��%���@p�$3g��)�^B����ï�<�j6��(u�Z���.V��<��n�W��B��� aۓD�ن�<
[��4�W(Į�\���B��
z��-1�Y��́԰������ܡJ#�F�O�6��t\�!�U���"��\"j�#�gMc���"�i��UEt �y���û�����Ռ�۰{1��[C�ڣ�	�ʗ~���Es�g���/�%�S�%�w���6��5�z�߷��r���C�d"�"dGmRŏ�x\h���
�
�3�,J<Kc-����.{��iH.�|��cR`F�����V����,~��G�$�ЃF��5��K/���s$V_�}���H�+�БH��!�JE��o��O�nБ�n�������2a(�U���I�MARאJԎ��?�s�.��n����u)��v�g�-�`&����3��0 9J��
2�SﰙO]��|Hd+W�`�C�H�ְ�`�-X�|��� ���%�Ē�F7������%z��4����;[a�_b�Y,�o��Ґ��!ۮ&f��1#���޿�/[�X\ ���D_5���<z# �dz���5.\��kPgW��"fє�I��?����Ch�)qa�8�p�ϊ5�.�C�Ց�� 8�V)5%麄0̊�y�^���eR7�> ��ֈΛ@��@ �0��W��kF���|�N�͂a^1�
y��4��j)���y�� �����`�)4~,��9w������Nʰ��ߗN��8i9m�kp��\��CK1��X, '��r��@��d��)B,�~Mڛ�	ʑt���c��e��l�n�}K)Y��&f�.�ݕ\:d�P�71���{J[S��9z���asR]\��R�w��k#��h���yʈ�"#E�%��Z ���)���:"�]l�2:��38c��)NbJ�j÷p"�ḳ���\;YW��`8;��37"�J�X�7
�+��{�W�mMS�8��p��Y�F8%�M�S�������鶛jJ���d,�ݧgDXk�Z��T�A��7O��6dDM�Y�4�g�Z,�w����'�6��~���5��� ׻(�`͊�!����~Yƶ�ȩ� ���!{�F��Q��������%���)O��ԕ���
Ry�ќ����:1I�׫<�1?��i��
uNkKP�F�g��O�e�D���F�;��\�������#i��䏌����|�\�:�����ԧ�:�oS��I?/�Kg�ʦ-~~؉�I�<�p%�M�Dk�|��"�o%P%l��,?�A=坈tD����W���yO2|�󻣔9����>ߟ�1C%V����2t�Bm�T������J��g�W��r� ��&�]n���odA�+����l���b����=�Z�9jX��QhI�+���[n��O'}��Wq�?X-����@��e[t�/RP��Kê�b	�k����f�5�I���8���o��s�F�־��.�;RT�o�����9fqli�N�-D�a:dV�[��ѱ\ �ٍ������_B,��K�oB��m��w�v#מ�,ŉH VQ �1=����9��ٿ�E�E�!Ѻ(HBG,{׮6�
;�Q:1$��EB��H$�n/�P����
=N�o��������7u��E���<t���ґ��:4���~N0/��zp	>���)�n�ͱbT� N~x���ӳ7ZN~H����W�6_�,5al�9y��,�o:/�yK9�nxF5��'lWw%��N?Ȟ{j�!��G�������3���D�*�
<�oYf���`�G~��߽��H�+<�Uns�/�W�̝yC?������S��2��{�(*t�=z��I"�!�t��}���9�����Tɒj�>{�El˗�\ގ���L���:�{t�����4� ���&9bG����Տ�>��^Dl'º���."�2�����'����C���_�g������_;��_��~rx2����T%����R����B>��*�sP_�ޑ�[es���I�'�����%Kڜ���s�Ym��_F9��}�1�W���Fa�K ��<�Q����u�GtjnM,�Ud8j��Wh�<}�h����2�l&D G2��60�-7�Ș�;�ch܏{5�1 Ĉ��)�w���8�Q-U�ZB�l�2�����Q.k9��m�1�NLH��P�2xĭ�.ED& .��B�FX�a�Ix��VSwm�R'��%�$A*��z�$�y��$��7��҉�����}� ��;��2�wE��q��ϼ����b����T��^S��:Ph��9Q�����s���exG��� 9$c�v�Ixj(�b��dW�0g��w,��׆Z��C�7����.�$�G,(�ᴌhpz{0ٷS4������I%?�$��m,I��$l)se	�zzd�l��Єm�ݶ5������b�0�s�;$�)پ��rou((]x���8���	��[]���=��l�R��C����5/��x*FB�o
���K%���p��~'���f֑�a�M���9�
@��^f�OGg������j���T�]�B��������9X��;��?���!��H�o09���6�s-�r��()~��Ǻex�&YI�@��-���%�_~�ClTΜ�ZULsf�e9�|�����و�t@���&n.����Qn��^�w*��fwPCآ��7�(�h��WZ��1@��p�\�B@�����J/n�A)����5>#��ʊ�S;�����Ӡ��x ����7 �8���̹�#_�Ş�t77��햞�hu�|2�
���P): ����1Q�re_)&V�:��abŔ��EN?w�d�J���f�Y�(?y�q!�^�� �`6��jL('�����+�r	�4����a�y���Pt�n���;[+6����b�����5�$F;q	��:�N�L�t=<Ʀ�����~��M�� �3�����G�M��0.�ܑ�2���s݈xF���&����|s�Z@8p/�jCy~%6��Td�ɣM����ˌ��Q��R�$w���{4h>�h`�Gj����&�D�T���.��-��w��Ӑ�H/{ ��HU7�>��gma8֊����� ��]d1�0Ss�tU:/��r ��!�m=M�����niy��ڊjg1�'݆^�%%�5:V?�e�]a#���_����d5>Kf<�g�8�����O�S�&s�,�|�0`�f<z�?�μT���i�o��6"bz�̼�>��|Y�=)�wD9x${Y{ ��߰r4j��d.��x^��u0ˀ�Vv� %�����ƭ�p�����^�=�<���x��zs�Hm�,�T�(:o����:%�%��i�N0( ;�4�_���P�5��%�B���)�J�q^������5�n�+4�+�ش���3^��|��1U�����Ȕs��X����*DD�4���j����x,�2�[��1�����n)R����X���h+��~WXCf�\�1"���g�b��@��+��*Ƿ7����S7��DN��V��l:�7%|p�þz������<p>H���Խ������M�� �,t�6Qg`��Jy{�2	؝mI/�xpu$aL@~m�!��6bɴ$>����EM4��N44�#%�Voϝ���V��
^��s���Q(r`h �� ���ݩ�֯>�Ko{[�S�L��$jTr1�"�5�l�
��]��3��~.&��/^�F_]k�nw	�(�9�����'V�2�.'H�'(�%��"M�Eӎ%6�r�؊k���b�C���u�tI��)�ʮ�;Y�V���R�Bj��5��\���g�o@��mU�}�FE��i�R˓���`�P��l��/�Y�-��$���rnէis^�穀�۰ˆ��T%�����7Y� �G%��E�r������+��t���]{	W.=���@x$���/����ǿz.�
�G�P�"JR�-k��7i�$ P�O!V�R��eR�v|B�M{x�fʫ���	#��9x���XD�N�EMϘ�iik�>NC|1�z?v	��Sz|��~���@p�eFE��Kv�C&fl3�g�t�EV�鎔�@���Gp�V�*r�ߑ��|?�02i3�|�@���B�F
���̟CLӱsKF���@�mb�����u��O��]��l�o&!<����3t��� �Y6�g&�Q:�֞7E('M.v�qP�˭V�E�>�p�%�x�|���fq�9�q5�m���I��� ������j��?����LG~,�H=5���<�A�$G��n2��x���b0L���!�*ɧ#�=���v.�����	.�����+\P�R�n�6��+�/�o��i3�iԴ��-W�ٟ�(��2��IsPd�_R��Pp���t�p�Ǖ�!U����r��R�iR�Cn4��Z2f(���Z��:�)��^����-x���op����}zS��F;8Y��,���i�����ʊг����	d�AӋWJc�n�l:G���F�n�a��f���б/�^±XƌU�(�֪����t5�2�umS���K� �'���e�t����]��:�y�Q\<5��P?|eb�r���7��^���L^�9r1��N+�1��&gF �ں�Zx�Ol����xٯ�ێ�����Qn"�|�&:��$�h��һ7=Y�l�v.V����+xrK����|�|��(puJ5
蘧8I�4���%��F �a��U𹒮����c"�\��&��]�>�/Y�E�����$�PW�c:$J~�a�:���!���,�Ӂ�%4��Q�u˃�Ӛ�P�+aF�)��d�T��f�>�fA)v�X��R�$��X��T���4@�\�<r�͵�ě�����?F������x']���k�ws˹��Ƭ�P����&�흫<�������$̦���Py�v��_ ,�h��"�B��H���1��n�ug�`�^�'͟^��O�}-%��Vu��_S�+c�u� ��`�ІAT�M��DX��0��$�O�����԰f,�����(l�X��-Xf������4-��<Ɣr0!Q�d�yLa�"`�������[G�7���PH/f���h9���G���= �^��}��9��K�ۼi)�?~/�`�M�X_��z)F�����frl�u���B�IyP2QRo��7��Se����?�]���v��`6l٩��1�te���,g\G}:l��,�q4 :�=���s��!"/4��y� ��4�x�@;�5��ɐ0���eS}�&%z�d�ҟ�˃��Ĕ�S�2�:H:�K��*�����	�L;@�|
�3}�H$��kL�<xrb�^�|=f��%���
`��������Xo������u�����A�b�ӽEBP�"�Q�?�dl�k�l�G���w�8��2i��_y��7�4{���q�g��4�ǒ �H�K�L~�����4Z��_>��g��e���E���q��;�M�h�p	/�����\e���ֺ�ߒV��3�a���O(��̟���e�.q�[R�Ot��\hm
r��,cXe�#�+�'_]�^�s���-D, )��+k�K��\�m��
(ӕ�rH/�q"�4�b�jM�e��������쫂Y{ RͶ9�gN��FÂ�b��#س�#���-�} ���LI����tr�)O/4�a��X��&w�;�L��V���/�@7j� �.��;��P���������D-n6F���]N?�O/z���U�G=)W
�W���0p�O39w����Ԕ��o��5r�S��x�*�&�mX���y�+\�~�M"�,#��t��CT}�Ҳ5.0�@V��g�s��n�Q&�^����	��GE'���fUp�>$X��e��[�+9g�8���* d���w?�8�
k��<���N� ��H��R]"΄��+;�!ЈE��k	�\�H0��A�s��kQ?%���\������r��ҙ�8!G����Z��M^$p��q��2���_I��\��2�1Q�q-���X��A��W{VRի[NҔ��>�x��ª�|��^N���w�#��u0�N�수���48��@`q����X�Dn��r�{�sZ a�+����J}p���]�!�Bf���4+ě˖�k�Q+,:6�=�6���X�8;�	T��օ5��4���j�>[���n[h�o��US�ɰ�Y��SIY����)���t�1��?h��Qs��J �����)��ڋ�c���Э16Y�K���灃KIqL�?�2�V�W��ge�]pY��^Vn�B�9ϰ�
%~�[����r��|?�ϑ������1�I�O���/tI�I� PD����7�c�\�e��o��3#*�OE�G8�ߐ�|!q�  8)�Q�n�z/nΠ�r���~�����)zb���b�O�{B�|ʁ�;��;�Lƅሖjj�GRjk�V*�0��j�᠜�e����E��j]K�3�3oм��C|���c�!46�[(�YWN1����0��"����7��>T��n����2�8fi��ջ� ���?��D��b��й�lG���_\�;���OS NT-/��>������.�=��P���#�k����0[�q/�JAzW�	F�lIQ������S\�Iǫ�1���8)�6C���������Rw�$����dmM�M��FǱ�%����gIFJ�;���e
�"'	#\�&�3;�x�V'�����h!��d�
�J%W�"��|�J�k��*��6,]�D�����	}I@�K�t�6a�Y,�������hk�;-\�$���Urr��9!k:ʑд�mq��|���S�4j>�I����������)���E�.sU�t�5��"���"�s;\혧򅥷_@����⌄�^�pM�ɕ�/����7]pE�;Wr�eC�� �<�������T��Ӹ��Z��A�
��֪�2���t�w(�~��&��U�87в�{{��Q�jq��v�*:��I�h�Ӟ`M�k�x#c=�VZe�o��ޗ���A2��l���e�n��=A�=��iDU�R���<P�����E����G>�QdJɱ-�yH�������1��2w���7ڴ��G���D�HSX<\�6Ě����<PO}�w��u6���M����O|��*[ԝ���tP��!>X%+;=�����R�C�A�?<�O-��3.��M;�,!1(U���Y�E(dN��A�7�M8�?��1걉�C��f��q����LA,S���]zt���H��)�$bպ0�S���K@�f���<=|3�mx�ѵQJJR��bF"uɨ��<Ùr���U�2������o��7������yG��s��2��U�QaS�L
�B-�t�0?��X����֐�(�pr=,7Cl���T�r��q}Oh!6 +j����Ai�1rXKY��
U\7��Q|�]��x��Ēx݆H�TQ�"���Y�׊Iv�����Jd�V�����$59��ϛo�����K럁���eƉ�/��t�g]q���	7�8�5��e&�[����Ho� �� -~���՘*�5�K 5Nj�)?hLS=�y���6֪�R�'3{����f�����9pC6��Q�}���
��q{�ۉ������v3��vǏ�D��e�Yq�ɺU��z���/�?�]k-X�� ͗W�Bд�tΈ����>���ZJO�Ǿ�W~2f��c�W\:õ��s�/��:�N1�]m��I(ߙ�r7\��&�{u���Ε}�'E���q�"&�s�� nFk�*��Hf%O&S�' m���J���QW�篅S8���2��jpO⻟��&�~E����tA	�\�Ҳ�%�=�f��|�+9!��Ci?ҬK9�EA�� ���?��V�ʳ��@`�ᯐ������s��!%��K�s�A�����	]��uhk'~i]��;h��m`ap��֓�Ɨ�1egCE˷��H�W)&}�xF�x�x��zp���qk@�5^�tc���z3Kzk����Z�cx%v�2E�G#T̓.�@�"Z�]��ҍBu��9!p6@�ٗ��Y ?!���_������މ����m9Ň ��κR���$�gl��ǿ�ڲ��xN^Ȱ�]*�0������/J��_Q+�3(�((��v�ɵٰm.S^����Ή�N�a^&HX�E[�����yY���cڥ�tji�͕K�T<e��y�+�{�
�E9�`��N�b[b�4��9��-iA¶�2M ��6���H��Qe�G��
���%��yf#!���y�y�Kz$<�@w�|6�* x�ްUkk"�g��s�L5sr8�DogI	�{y�量�~ܦ��}抳�l�p�S���:a�
�>Q{��N�����������ű,��iN4�}�w�O������� lm��ˣW*ƶ˹�&\�j���5�n%'Ƒr����[|�����d��� �r(����V*�V�5Ϧ@��c���q�"���f�e�GC��`1��0`����:X�p����0E���F�o\���������FkOV��$:ul�3�||&�9�L���ej�.�D3i�FL)\؟+�����k��=j�3��o^$N��i���%��H/mÕ}�a���i�D�y�3}�.�����&]W�mS�l���(�Ke:'-��Tﶘh�&��R?����(��kxB$͜��\X��m���^]�%��H�>D�J<P}�[dپ�ܴ7�`�p � �� ��j6ڏ��c����e�xPl/�B|2�ڗ�!�sA��'�*����14R"�%�
:��5,;�G��q��nx�s\��E�@~`���G��b��|-<nSv�p+���Cɀ�q'HEl�>.4�OTo+A��f����r�v&��eC,Ṫ'v���W̼��W�d�
�fS��@<����:�~���]�zQ�{]y�[�"��U��S�I��N!�=�ѣ5���JS�0��I(HZ ��Ÿ+�Z�%,�y�#�9�������@�e�O�Ax�
�^�r��/ZI�҃7{���������3T���a��Dr�N��Ėf&:�j/�"ŧ��,y'�h���~������ޝMb��"��{(�Rh,�N�<%�8����� &��2�]ʺ�����޶%�HG��c��J��"[B($<��u�&�Z��/��3|]cg4��W>w����Ws�l5��^S΄_3-�@��=q�f�;�%���a��F���e��a�l�06)�0�x�����q���θ�����7oZ`�׹�"����r�;@ms1a´�u��������l�lq�c9Z�;��I�d{O��qz�=!�R+'��~��L�@� xTέ��f��2u��K���ߪ�@�e%��茾�D�n*�@pY�(�"jU�Ur��,��k�U&�L��Q�x���z�����r���fk=�Hܤ�AZ��IZ'�4sK���z,��>+��������S�lk}5�ysڿ�`[�]�2�/ƙI��sP�$����B�ىd�:�-EM�Q��%ѡ֌�.�GK�3�:@�<�zv`k4�2:F��6�m�\�[`
=��5���Q�%mp���y�=&��
���š�{����	�Q�R��g��� |�����ek�+��S��H�m��:Wż��������+��VS%�.��F�P�c)�������y'�X����xu�ց�jL�T��&q���/hZn��k^�ֲ��a�TݒM�f|�۟��
�	a!k��G�K���X��sH�m>W���;6 ��ŻJN��\��'Yc|�����MA��y@��)rf8�v��>x�.�� _93�rP�/u���X�/�=k�9�"vYƩ=/�%�����ۥ|�3�EE�A������=������6�s/O���%vUN�zX�>���:�����di�jp�`O�դAx<�q�^�*6�?z��Z�x�z�
��#�`��WH�ۡ�oC�,���6�[7,8�|`^����| �=�g`����Up�Wf�>��(M��%M��]S�݅|�[b��Um7}���ɶ����ޠ���Tq�1���t����)�(��M� Iz�BjQ�-/ɓ/�/���3�|(������|��r@~���ܺ�W�r(��aB�T���ª���UfFqC��p*Ȫp(BN���/ZZY�?��z��<l k���$�7�~
2��m�Om�ex��:f0�$S]�xL��E/'+�K��JO���>24Á	8�#�s��Ҹ�+񪴩I@��4�K{���Є��$��#n��L���e��D�!L�v��>�L�����Y�l#�z���w�_����(=_	�#x7�gΪ��h�!��P~S��4{Ş�ѪH�:�R�jEEy�_7�knfR�p��cU�K�� I�wXl���3���?60���D�o'��hW<4a轵%蛼39�����d�o�����	>|o[�p%)OP-�@M ,fP+�M��w�=H@M���w|7�+ �
3G-��MY��_X���_C���[�/�N�������ռ~���T�z�d;�j3,�8��Hq�14Q����K8�+�\.F��Y��z�-���"���Mmh�g��s]i���}Onu��K�5��HL���WƟ�J�4;��s�dy���谕�S�%v}�����z^i�jo��Gq'1( r�+@Hw�y�΀*�0�ÃD�yī߻�ʯĥ���(ۈ,�W:�?>�퀳*/n6����1�ԇ�iO�|W+w����ɨ��v#��~7����t���+�<����>�3¬1���#�\�A��������pf4Z������"B��.'���@Z<杂צ��$�O��>q��3�)��<�W=h���K��,���6��~�. ��bC�VN�,�U�~,+]"�F���E��ژB[3�Q��j�{-�@�C�$0Z�DS7�{��f���"�{L��'^�EX�6�vEɐ9��(4% %t?(�;jK������0��T�E�)m�x*�ES�K7?��o�_�o�F�-�*İ^Uiq3����g�O��4�bG
	+X��gCE�����a�YQ��] �r��{����T��m[$ӫ�;�`̭��>r_^�j���� T��eIU6�9<I�[�����]0�J�_:���T�O�qH���]�YM�hӻ�f|���W�鰫j��S�����h[��1 ��U��6س��}�=��˔1�ֽn��!�B �[]��ϧۆ��_�������I(���d�y{8����ތ:�~>�ݗ{�X7�L�¢-xA��<;�����H�(R#'���҂Ő��g��톏p�g��+����>.1'���7��o���B�H�/�����?��,��D�$ܽΆ��ק��m��ڼ<)�7��A�I�o_l��S����-��WCE;���=��K	���R��>㸓�+=9���Q7qD���<?���	�]^8[s)ʫ/1c����!�95�͑���A��%��=�%���T��O�8��4�����7��Om)��G"'?Rr!~��qs��˗�j��W�D�L�΃�f��m�yh���+�,�Kn�%^�R��B�7§�mT�j��c�_(D�n��L��eD�v$����܋A{O˴��aD�N�bGs{g���
R�m��g��aT�Ș�� g�����V&��M�_{�o��>p С$�-���xB�3f�U����Zq(�P�D��?"��EE�]��:�I�=bq��{��U����־�t�ر	��ɐ��Ƞ��}N�F'��B�S��ǗlҩD�]O�
_�XB>e7-柏A5�HVv���4鸅�7���f��<����#L�6"K�&�Ro�	����:��K��vT|�Z�����Z�'ߴ��X�>Z��c���a���W%G��3[����ģۆ$����y6h��~-ڌ�X�a���t�uMv�Ȟ��Z�r��)�T�,]�8�F��T�~��;�JsjɄ���6�fEh�lR���cl�7g�0i]Ʌ�w��Hx~������D��	Q<�)Rf� ��y�'��"���(>�p݈=�'�g� �bP��Y~��&�W��m�Ҟ92�<��,R����ە�E..�0���(	̺$~F�H��O%����5o�vJ��r�����[�FE�����X�b���]��Wۺ전�WgH������ ,<��M\i�U!Ǝ�$)P��c���
)��9o� ���0�G���k`I��X�G��N�m�����/��`>n�^�Tڰߢ�S��2r�ŹՌ:GӁ!(�|JD|g� �v�]\��܍ᑅ��Z����-X1�t������@��#)Q�(m�B�
�U��]X�<Hɋ�O"��8yǎ��?lO9���}����Y��?
�+�|�ZA���ԡ�\��gk��7��C�����Vᨒ��>²k��E<�Α�o�CӮ�����y�ռ�j�;��,ޖh�*_Y%bO����D+���)S���n���<��գ mi�����RO��ۋq�6�[[@LXCH]�l��gb��2JAnD*����
���/"�q0� ���9�@�J�Ox�ڠ;lG�>�	�ݓ����>E�`��7�٭ki��f;��\��;~q��{!�S��>�U>�����=�F���e�Nj��
�U�^g�D�����%r���R݋�&QU�M�P*.�mS�<�V��@��f$��X\���h�<�����ߠ��5��ܢ�'���/�-�]���+�~k5f��b�O��_��
���J�a�=K�\#���'�\q]K���3&s���5��ig"��l�M��M� ��SJ���t�qHʨ���(ߤ:�ɦ�\Pp���u����e�{r�*/��E�3�P�R���ַ��z���a� C�փ3۸�-�(�5?���OФѫl�q�A�� �x�Y5��l[ێ �@s��(W �g�UM�ǐ��In"Ë�Է�ۛg\���� "Nn��ɰN�vJ��cޜ�~�4{L����p-�È���|cQ�D�I�y��X�btrj��㊨w��Z���gqG��Rg��Mr����m�����S����K�ǎ��+�<�_,BM�MV�b!��guRQ����|�(o��r��padZ�[�M�[L8��m|�O+��� M�`܊���yU�~2h#X�E*9Ɵ��	=rQ�Pg0��] ��K�\���v��MP����h�9���L�M�R�.����b�m�;�z�:!h�_���>bd��k���V¨��h�� c�*)�ҥFv�b`MF#z�'�)`'�(�/�7��:�Ҫ=��t
rz.Gv�<2Fp����aS��!���Ö�D�#���D���~�`n��P��
�1(\��I�֝]�`0p������o�[���8�%<��a���n���Y�d>r�����O��D+ݑMsF0�М�Ʌf:�ˣ�唉��[�"�P��7d捭�r.�Y'\��b���	7�?.�	��yr֝�ml��~���QƱJ6��gnx�TQ�#g�G�~�޶�Բ1�����Rg\DOw��F�ta���T�Ie��j���/b0&2R���q�����?/=/y�=7׹�n��G�	^@��Ɇ��U��|��h�yV����O�;��;��꿻�H��msM����[�lp���-���6ČP#��Xi��f]�W�ۯn���Nl7W5���x��mg�TG� ���߂**��)*�Z�|��Þo�`��E����`��(��/W��J�N�� �����,P4�5d^(k@�)�&�N=�Zּ��+�#z�����>võ-)=�Q|A$��b��K�O� �E�B 1����<�Ȯ�1����a_)|�d����m(���`:����cL7�ƾ�lf����BO� il��'�l��oJH2��r�g��^�JA1U�m�>d���k��O%�3ٍ�_����i�����c�
�ฌ~���� ���f��./�'H`<��׼˒���"� ����tb���%ޙX�j8�� ��)J���M���<W���e�޲њ�y�q�V�K5���vr�3mNT��m,e�D��1��̓�^��P%�6��ū�4��E�nH�zגQt�y7����0P���K;f���i)�%M��0�-#�!R���yj��Q�u .:�*%K���T��Ŭ�eIŕI��Oܺk�� ��ax���l@�6̜���	�UFP�oa�/�oV�/$�Z�k�Es?��q��.��߱R~���O�#q3}+塋{ƅ��o4^���mrK�Gε�v�{��w���uϙp�=�X�����d�k�(���[��h%Հ�l!{4D������8�C�(���(/�QЪ�d��k���e��l�d��WN��ar����!ʢP<1	�ʎ�<�u�F�T"n/��4��D�5C�������)��#l��<�r.z3�����l^D)S݁��g�	E	sH������ W�޻C�B�=m�]׏[�J�\�1cVJ�k�� �+�����Z^E�EU��Y8EI����(�b���/�EY�ʩ�l<���P��`e;hF��,�Rm+����7طq� �Nn��;+�Y��=�
���ZV�6 ��^�#w�`ݥ߽-��	$��\��'����;K�]:�qI
���w1�Fi��3yg���z�_^@�OPh�Wa=�t܅���}���^�"ȝ,{U�I�˞ZlO�_S�d���HF�H���	��o#��hH�;
iK�� ����x^�t�O�؊2�U�L߂��y��;�f�k9��f܎
+&�D�AD�I�d�?�og�~@B�T.�;��z���=��EQ�n� =8w�y����X�b8��;�Ζ��X&����n0�'��'�受�W�/�&o�!x���
�^*��MU�g�uS�G�mP2;���.,I�iC��B`�\�5�Q�&�!�����$�X��\$e	k���UB$Q�#_�X�f8�X�7�Q�׿�pH�bBQ��̚C"&�#�&���O��ZnK�.8wF'���珊I��T��I�>�ƻ.��iK��~��y���q8r�N(�-�/,풾�T�Xnd�"'Eδ�&��& �7�~��3Ȳ3�I��G�v� ,���o�;Ѐ�C���_@ϑ�<��c�xW�Bol���t�w��ޠ�]��W�	��eY�؜�H�"(��&�!�<m�D߿}�� �n��+~��fOe�	��D1�����mĮU|O,�X������cq���	����v��!�V����+j���Yq�����H8�ɤ/��^�d�p;W�S�'�p�S��q!�/g0(��4��w��{���x�d�	j���ų���_��+l^���P��0���G�o�x1�a�n?���[ъi�0�����wE�}������|�kelSs{S���$�7݄nSq�'���b:hۅ�3ډ/� �ެ[�A� 	._R�������{�/ȱ�ܜ��"5��&��y<Ε�s7�r���D�%Q�Yw���x�%1�3e��9�<KY�t9����G�@�{x��{Z���%��Q��(��o�F��U��+f�Y�X&Q~ �ݘ��Z���Eo��.�3�D�4�^�L�v#�Lm��j��>��Q�6��|V��9�^s�i](�O�	��
��oD�O~P�T�(f��~�f�,7�����bgVf�����}
6|W�ۺ����r:e�����Y�#��1w���&�;��n�E�s퀼a�<�]��Ӎ�ѷ�@┐Y�}��G ���#|�l��Z���A�A_a���ﬦ[#uWS��{��d�]twW"i�<ï��h����E�t��:Z/���10� <qY����ۮ�o��!#Ϊf���,�3H�'��t��maB��3ըaM2}O��F�r�U���.�7Ⱦ,�������7H��A���I�U`��e]����ӗ[s����ЏUSF���
E���ߦ�M���l�q�K`� �s�ωQ������?�'���qg��G���t�Xߙ֨&���EY�|���p�%*n;��쀪����,���b��=���U'#_r$��	�$ �Ă���s2[)�x�H܆�"�ܴ}r`�/��ё�q�/���y�[��jeNǹ3f�)���i���<>*\��%m\�@��xYμ���<����s�	y"R�|�&5����li�EE���C)��]�:���!����3��Hh��1��-z��d)������D������?M��E"�y�/����G���wZL��_�	����g�1�7+���\�LC~��Âޚ��*�[��g_hL�-�6�ڌh#�^]����"{���׼q�pH�
���C�z�<C�O��٨���mHvφ���:���Q���O��|7����扳_J��d2é��ha�@�"v\
�?�r?I	����1�|�5��wßG/q0&��'�e�6��`���!;=�\�C����|��8��0�����"Ѡ{�<��WѨ|
f��;�PK�?��Mɓ#JL)}XVC�zU�I��*�]m1y�I��ʯ�q���H����^�\�Z�'}�}W�>B��cpG>��a�jj���-f�%��G��v����bu�?��E'P�y`cH�s�n>��ݖ��g�`kJ�Y
Of��V�(�ʸ�(^�,�`�q�����/�����f�*	ԧVH�@�E��z��f���tD�+�-����g��Be8FP�Z���T�9縥ʾ�h�̓��d�oX�B?���抡�[,���w�Cm�E�$���1	m��"����A�YS�9qVV���=K!W>��:ǋ��2�g�f�0q�r���P��H��^���\�Z��,*�	 B��K���-!��FnB���i��i�#�{ٺ�i�nw#?�u_E+�zF �tq?�a�%�v�	� �A�ׁNڨ�y~�C���l�C�3S����'�L�x�	��gñ,*�Q�����%�hx�	�0��e����X0�Rp��_ĦRS�B�J�w?1�uk%��hR������ � ��V��3g�T����r%�� �9���0J#���A+iݣ�oBa_%�O�PKPy9��jc<�[I����+��CΞ�0X�)�t� ����`��9�P��3����(vI���N�|�Ǌ�&����[��R���R��бBLj��} q�N�g���aa����/�{�&�L,��"�x��̥X�6��R�Q�DsX{}�H���Z����)�fwc�C���~|��<(����<�{ ��}��=��uH��u�4���$�'�
�h>Td�Bh��0�����P��m?Y���|R٩g;]�]
�_��V`z��2�R!���\,Jl��X���4:�7u�J:��&�G�`�1�E�]%��i��fBdI<b�U�&���ۄaL����T��y��?Ձ�~�]�7`H-���Q��� �g;�jG}%.5�,n�0Po�D?Fd���H��L��<H��͒�h�V�w)�W�)>���ў�[��\t��Z��֙2* 6��=���`I�z8jv���mz��h�P6��^H\�0��6�G��4�.5�VS��#f흑Lf���ۻ�X�D��f����:R2�t{Ip"@�
�>�6���Yva)�6��>z-.������<���[�>: E�gF��G�&�*Һ�M㔓+��|��_�_�)��J�Dh��H�ı�d�m�B�!�R�ԭ��l1FJ��9�g�Qx���f��^u�G+$�[����C��[�i�(�'���c��b���������RcA�^h����	�O��S�hz�"\�n�g4�i	T��:���~�bs^ߌoϘg����Q~��� �%,��J@�F���k8�i��/��h8e�^�^�zt�0K[1�QQ$<:�z�h�(¯���;8�Z��/����+�D�����kP����(�D�����M9�s�u��ˡ��-��_Q#p#��q<�<�X��q�m{`�9�#��@QO�CA�9b���*z`���h׹+o0:
:�	�;��A�HR��d��tq||�<��T0�>�gc��+.��u������"DX��l�Mx��w;�X%��W�r����m��9�b"�^�V��%�;��epc�a����Po���8w$z�ѳ~���R��h-��! �$Kʂ�����+vs�E
�6�`6?iR>���%�r��.����V�5H74i`y�Y�κۜ�CY�0�<~��fm|���(-	wa������5*�����M82D:�C��[�v����uG����f ��A�-J���C+9ke�P�����bt�;�q��q=�B������^�o�����s��ǲJb�"�����T�|;�)�K���s��=�|ƴ���*�=��*�"mxp�[hӕ��<V�e�%.ፍ���L�1��<2�T>�/s`���g�ۖ0��G�Ne��)��}@��=bz	��-��h����n�M��Uzi�re2!Q���%���d��k�c�G�[[��؜�G�1%�n�o.��O-E/ơVUVǗ�ق��>�f�K��(�G���W-�@���h�T�-/ -�_ڂg����hv��y��FW�ڐm��׊����,]��N1��D̽ku�y�\IeH]0�d6`�rN3�؇6�s4�����Y��z�o�T��>�ң��n���OO���۝ˉ��)%&~�Cu��,
J������E$�G3���QRt��R��X*Y��FO�lq>��i^-WT��!�4]��I�AV�X<��A,XiXN�����s|t�
8��|͢&��kC.	�W�@&w�M_�p�D�=�a㎿�����j`}���i8}��Q	�I��^�*;�!G�1D;�`�?���;���_�H��>�`*�ٖ�?����!6q�	L���Qm b�:�Y���ߝ�Ԧ�rc`�ě�=��-x=#a6���:?�_׎/B�_�ּ�p��3W�,�ZB���^�����ark�!�k7�$�}O�%SZ$i��N�-�Y���F4�����}puO��a��;�u¿s���P^/p�A�Ը6�R=(���1Ec93	b`�+-��<�K:�A,��G�^'X����qI,6ޕQ�Y�
u��h����|Cm��{Tի��n]�Eٲ"ԣ�[B�L��Q5a����gl�9u�/��))o��C:�]*b]xA5��0�:Kd��!X]<����M�=q��w}a
��nX��Ո�ٌ����h��sb6�d%IDJe*`;R�{I���O�TDS$Q�C#��uI+�L>~]�p(��A���2�J�l�����c`�γwklX���A\��گL_�ęǒwG���As��`�o6a�K����C��#���2��-Om|MX��WE���7@Tb�?m�����Ř�Uֵv�7���+�>�No��0Š�$�6n�4P2��/�]�M\�����ã�S�q��(x�@�ZO`P�$����32^�jV��H��1�7%RhC֡M�:��z�Z�7S�Q��=4���z �۠�@��|O�Y���Cb��<!���2h�Ϗ
{�x_�*�O��&�6�̴��Z��{
&a?�2� ���JNbbYޱ���F��
ޙZ��DH Q�:���Pk��t���HS%�<E_�<d��7��uJ���#4�|����n��#�Y��x{{\(�rt�8�^�M5��ӳ�(�T1�q�a�@�]>��r1 �?���a�CY~�$�g\�j�&�2QPR��\���{a�0�*g��j-?��F<���$�{���<L��b�}�EY��qA��QPzŲ��y/ċY�Y�(/����tQ�r���[���o/I�?	�?2*�����?����J�T,�kZ��!���/�3e�5y�k���$;.^�k,��A,�?~Kc_Y��F��6�kbb�@"�Bs���.�� ��
A��[���(T��UL�2v\�� ��T�����(l5�'��_�	�)x�4F�Ą
A`C�cy�v��D &������x�$���HYr5t�$8�"zD��ܙ�s���^��`
�q���D���|K�{�Cu��ȬZ�-bvy��<�����y�`�>��6�]�9����h5�m��N�����*'�˥�oh��)W!�\�өY^��Q�zl�T'�6din��
�Y�#u�r����3������7�7��p]��P�j�#@�����{`\��]��˯��ܠ��*���)b��W���HZ������E�����{���e|���$�d^��̝�Pk�����$ �S��~��e����鋮~`��ul�+��� ���B��K�ՕE+SDS}u9�_����>�eu��VgH��WK���&�Q���Oc��`mz{���Cp��E�ֶ@=�<k�C��N6侩��Z��az� 6:#	����_��R�v&�����3L�R��2»Y�S�o�+�H��}��r6�3vG��>��{!��G�ү7�AS�v�Z#��±�Q��8��M�XN��e�E�Ϩ�_&=lZi�1� ѧv���SvA��E���\���`h� �G��UV%ł̷��T�՞��.��^�qH:K�@��/�Bӓ��Ir��Z�a8QW��%YU��-I�x�'�*��p_���ו���EkCiXl$<
���X�r ���o������Y�~%t]�(�Y�X2 Ë�?�O0�_�ٴC�,SF���b1�a�a�ba��а$p}p2Ā�<Ό�Sj�U�o�	[�f"�̧�cDaFC�yrl�[���r̆�p,�D�˘T�m�8K����z�͔G���]*8N� ������ܾ�[���]�m]�X˖;������2~L�y�Є1�����x-���r�y��sn=�ީ�n��Դ#��{�_�a����Y"�ΆgK����v��%��E��zS��.�i�`�73M%8fN�̙%�s�}��QKJ�0��<�}<�8BH~���,,vm��\����4?�9�|M��DN=mb/�_��8��e�������yؑ���T��a��e��pg����J%��+<���ۋ�"���AMD�p�FN�u���	U;����/F`���&�)`	���I�x���ې�r�|���@�l�ׅ���	ͥdÄ$1i�u�"Ǫ�Y�qǶ�@ՠ��F-�+:_����wj�����"���kL��"�\�1���=��k@��F��Vf��<���v~:�1����*@S��d�/��x���f˟KlV;q|loۡNMsnG��T���gH\-Ξ�E���[`�9XgZ��$�(HZ��2��h>b)���_���l�~uC"0g8�+�p���[2��Ž#J��	f���D�.�m^�|^GW�a�����=��d�l�a3fѸ�BϊƢjg�����#h�� �b:#�ȥ�[W���.�E�_~)�7���d��r�ϔ�K�鶻5��Q�ᾫ.x����� m$���UM�J|����fu<h�l�G͓������|�~�K����HK��un��4�<��T�?������Q�g~��d��l��:��L�Rޞ�e"�[�����C��9�1�w�*�#�l���љ�SqI�+Y
��;d'y,�?Һy*�x%cj(���RwЌ���F~ ��qoϦ-��:�fDR?	A�gfP=�������m���wwR&����0�m@u��`
��}��Aqj3$}meq�o�s#��MQ窪O�����̦��sĪa[`&�\0��"� �h.�uٝ��p�(�F�+�Ft��ߣ�?K�4Q?lM��e�����ڷ�I&$�L�dpp�yz"�nL(���2ԇ1$���~c�%/d[W���E��b�VL?>3.���`m��ossM{��r0�2�g��_���H/��G�G�L���3�a����΄o����x�҄A�WMc��`1�<:W�<�!�'��RUߊ)��}AO��2/aĀ��(ZC�_Oa�`ևx/ϊ)*��?h����
v �͘�c�����G�e�@���
�[L�4��������γ�t��Ѱ����;)�P���I�0�M�����V����g�X"|ߤ�B�t�[�e�z ���g��p�#�y}P�ˋ�����T��K?��~�;A�_�8�ϗ�4O`���HFF����a�Q�cwW:d�Φ�N$1�C�w�:�=��[�i�l���c���'=j�Z��&K�r胧������h�/$��'V̨�%L����K���Gba���s���t�����@�
�C8?{r��_02�K4`�����:LCBf0!�
WWVe��=|	�9���������mk��6b�+WrF�n�cZ{��?��ɢ�1x2_)î"�t	�C<�E��&�J���y(�����M1����݀��݋����6F��pM��z>{�<��Dz�"�b�3�5�n�I�K����.����V�J�0��̢�qn��B0�V�O�.e�v�����4p7.�8b�����}ڠ<�DQ�]?=�&_y�6����nބr�cA�Pc���=N�����i�'��Ȩd|S�c�7M�"9�G�U��!��V�����nlS<�r��b$Z�Ci�Mk��Ɩ�5dLf�\�u
��8�B��>Z58��?���S��-g����\�g���E�Ɂ�(���w��|��	�"�h�%�e3KbR%�Z1�k��ő���Y�+��p��l���?�{r�f�$*������6�2�G`~�U����Wڤ�~��8������v���T<�C,�Cb=o��Dw�φ�q�:�q;t�+ӓ�yX4�5���e�ejsu�����}��r��ed���M�M��yݬ�a
�	���|7o�	zl���T�q�{�Fj�x��<��MY�T�?�,4r�o*��:��jY���������q������AO)�_&H@W���m|�͑W���icb�"�q �}H-Je�=�U��'�ں5�#pU(L�[pY���E��[B�ɳf��0��������杁�%״ݽ�w�VS;����>��D�t���0-�7��r�
Izย�/�7��G՝^�lk�+D����Of�qn B	�\\�����xf�L7�V�,��_9U���aS�VABp�G�6��yOx/�M��0O��wM`w]]O���2�o��4��ک��~��	��L������ッ�����m� k�K��딢��Y�����ѡ�qdp��˫��䧻�.e�J�z��?B�ۣ�J�)��id ��~.�*��j�^�8�����h����\�B.-�Flq֥ݟ3I�,J�>� 6�8q�3K���aLSN�5���!�9z�mT�A�q/V��x��B�������ϝjjV5��x�O��V$4��\��k����B"�9P�MZ7�q`au`���舷�=�]h��x�	��ZE��+j��%/�1.��\�j1���Wl�a�Nhe��� �ЎX��2,����o���u�� 8�9�����1���YK��Ә����Txh�tL����s�܌^�`��숅>�}���Ǝ�;�\m���@�3j�`�탽�" ���Y��}{��E�� �ʧV ��^`�=`�ߜ+���
���<"&��@��=H��N+�%�/��J�mYJ]^i ��v��͍�Ү�����G�]���e�dJ/�䈃&��,� �-�!U6���u%��kl'����G�x���b��Y�k2�Q�x�,%���z/�t�ĎY{��o�U�V(��"�kR� 
;7P����Z�l���_X_^�H����>}[@V�we�s�a�F�s�/�vո��]f�~�d'X�V}$c�\�Q0��;���m}��<�����C]�ə�8qb���+��[����	\�O�yI�Y�CgW�Q8�%9�G�Y�X��l�7�;',��PGk�_^Ͱ�I:���2�>�b!ࢂ���t�IƐn�K�dh�ʖ�o5��2�_a�?���ֳ�hx�V�8+��e�vv6���gN��^�;B�VW�C���we�L�	a��ݷHp��64����Bt�9�k#�p�O�n\~u6ᮈ��.v��}��S$Cnj���2^�����Q�9�c�n��-
�7��eT��c����x��&(CK�R Ϡ�`B�?�U5.�q [��;�0��x�O>��z�nHS�қ#+e��st���X?y�.X�� �EŊئ�|�F H^��u��pa��~�ߚn�Ӊ��%n��bZVd���"�pP5jf3<:�0h��-����-+ ��	�fGp�(,{��������������Z�Rd'��O��	���i3�
��l���QEHf��dZ�'���&��L��.��8뷕�+�(#��R~0�vj� ��x��<�ͼy ���FAY�2A��G(�3I�
�l8V#bj�n�� �Q�z�?�>��W�h ��23jF�F���"�2�8�M�{�ǂbTM���g� Gtaup=�dU�gη� ��"'#5#�������M6�Z� ��re����(��ꥉզP!A�@���Od'8H�JrzP���yݣ߿x���@����uP8���D�U{r��m	�����[A��5�Kb�H3n����1��eWC�Ky�,7��� vCB�-z� ���5B�����H��)�QAPs9Dȇ(�~�������{�J�����e�!�]E� �B�Ք'���ɭ�����p�6*�}��cܯsY4 s�G�~�n�q�TT���ԋNƷMxaxd>ۇ�#~��[��Q�R>LiM����������*~wa��9���Jϩ�	���Љ(&�����v&d����͇O~>o������y�N��4���9sq3|M��ƒ:9� �;��h�{\�xm��;��X� �?�.�6J|z��,�dP��[�!��)�Q)W��W&O��Jإu���U���6C���X���t�\�P�v4��@�ͪ`���g�^*�m�SN)XU�>9�8(�%�� :hE��<nء4t�
���" �)I�-5z�X�[,ԩ<�=�`[Y����n� 0,Y95�#�_a�o�|y�p+���MDx�S� 	NJ�E��@�̪��ȖF��D<���--I��km#K��~�E6.K��f���SU��D�폲�K��V�-A&£�n-d�/��
�j�̜�/���A!R���Gb���!�1�;3 >:�P��hRS��Q����zd$ob��}�].H}�����z�����+:��%fW�DKUm��r�;䠊�Ɛ�?-����x�Q��X���CM�C�����d�ɀ��~�ꧣg�Sr�\Ki`Z�t,s��|*Dn�wfq)>�D`l�!@+���1��.�� ��Y��1DF�$F�v=@���a��ǧNM��m���ܨ�Z��G�+0��BnH�|,O��M�Z��D�����J��wJ�r���g���M])�Cln��l�h�� %�.�1��k�p��x��u���Q�����7��)�"�UDn���h�t�q
�Uw/��A�Ps��u��;�9�-%a	�c�9���ݕ�snA�����1=�����^�R�x�~8o1�=�� 	UB|x���%R}�V��}����209�$��r��Nf7n�-p��@�RqŊu���N<	��;y$��r����O{7]�˜)P��eP�b��&��C��S]���h���:Y����\��{
�~�������y6.��:��]����X���|���6����i�#�9�б �����(8�4�U؀��6�t�8%h^�l������TF%c����e�����:=�Qڠ���{_�������/�6�¸�a��4�� ˂�}��]͓��=�[��UO
!}o1�Г�Lǌ���Z|�?jӄ�I5cS.RR��K�q	/5��uEE�����u����4�u�> M��@�#&	��w��-�{0����J����L�
3X�u%|GEZ��F��1&r0����d1�a^��t��nC�� wZ~�S��!�%5��G_o=W՟=�̿�k��\w5�ћ|	b��� �RQ�n��{��x'�a3�9�"��/�ќ'�e@pA$t��N���[��èK2Ք��i�D���f�?�=i�,ӄv�}�na��n[h�*�-x��BQct�F|�6�hw��
���|��F��T���6�N[�)��m�jN�p�)jS�zC��4.��GA�+���L��`�-M��8J�c�A_��6�P�G*܁sl�H߫^
G�^�#r�9��dRH����|����?@��qm֨'����.d��=�읁}�sҚ�u0;��.���aE����r�������!���x& @��go��Ț���8�;���ěި`�g+�Z��T�ә�<���HHQ�7��e��b5�V�Ĳ� uT���#|������;���k�� ^�HRY�g���n|�i�̖o�~�d��rOu�L},Þnw�d���nM�]o���'�v����gguZ�O��1�83�e]E��0�.��\�O��"ӂA�����˂�E�{t�!�+���G��	�U{'§ҹ��K\:�E7� ��p^-Q��:xa�o�8�m���1q�F�Aw�Kb�ޘڄe{�����}@ 3����&�i&�t`h������u�\+�� 0e�\��h�'�r�-X3l�U�I����d��6]p�&m �⴦��+��.���@�uv��!���Q�$%�	�K��Z,�G� ��x%ǡ����� z���X�8�Q�i�7�sr�[�t�Β���9]������n0?T)�rjj(�������� ��[~�����՚d=�����G�4��q�
���(�ȯ�h�� ����
�kJ��N완S�U\��K�$Dc�:n�_6�2�v���oU�S&4Fio3L-^9��:��c<�+����?�tKϘ��y\lO5=�"9�h���ԇ���5ȴZW@x�A���[��(z��Dln�����7l�������@ed|�q��?g�Yp���Pw�/�0�N�N�gJ�늞W�_�������I���k1�:�g�-I��C�꼇�(vW	�$+�Ę��N��̶Tpv�Y�B/zE9�G���܏�\���N��E��,/m�t�᪻o�׃�9k(��{%m��U�q|�U*7�Nz�#������t�r���j\D���a�(�`14 �>��Hw����M[A���N�|0ؚ��U�~��y�����3��/�О V��A�(?���֒ S0,�9����ӣ��x�!����.
���[2vLvK�߱!���CM%N~�0��:��[��>�"���\z6��߾E접g��4�k��P+Zz�Ç��}e͉�E�P�q��zK�k^�i��O��
H<;�� �?O���{`���Ot��Z��G�m2{�@�/���}=���d5&i�e|�s�i���6�i�V��5�Խ&U�S����~މ�>���� g@�\ɤ��ҋ�.�P]�^#�n�=:�aܦ4��;܅k�`!g��+ p��ac]�G� ��H�l��F'�Z�i:�&�M2�f�Z�bo��d����LF�vĭ��a��!��6]%���Y�橕���\f��t5zՎ�XGn��_V��<����F���p��7z�@<��|�6'�Z5s_�s�e�<�"������(�8w��y��9�?���.0X�x�v%��~�w����VD�f:���{1��j#<m��dPi��K�t��hn{�˻)��ߍ���5���Ը���,��a�b��5uSGʰn�Y$��I�^
���(����I�76*��RɈw�{}W����D�"��g�˃PY�~�8�Đ3���"Q�_�����7�ceYO��r���Иr�|�������S {чY9
��h/1R����3���Vv=����=�.\�A�>1�&�`T9!���H�!2D�ո���t6h|ƻ<�l���`�<V�4�h�"������M哋��V֊`g�4� l��E��!��� �X�͖��1�r�t\X���{�(��-E[a=Z^�rZ�(�;<�a��W�Օnţ$w��g�C�NNyF&����5HQ�c��˅�4�݋s`)��m��Ĥ6���6h�bK�,}AHp��91z�i�:�a>H��B��T�bA�n�_
���:L�m�1�'5�m��l��[̧s�u����Hg7,�0��i�j�jB���IN.S[sX�S�׽�C��Kfbx���0ʑ��� B�q����#Q�38%��@�Iܯ��[��iE��An�l�S��P�CW<@�z�b$e�\z3@�I �h�PګRt�ղqD�g����-Vl~Z�͔����ꭦ�h3J�f�*��y7;����������h��Ή�_]����A���H��!ᆬp'^��V��(�H ��Qó�+�Fe
➁@ �ް�KI�P�/�N��oθ��o �.��*�\	���{�,LpG�l��G��-2�d�T}��W)���/��¬� �KoX�eL�=�/ւ�Z����择�2� ����~UP';�ݪW�\�s�z�O���Lk!��s(�S�b�m<䭍˨!���'�b�#���J'\|^�=��mA�A���~�H	q���l��l]^�L{����+:�(i ���8����ۜ)�Q;{P=|!{ekC�k��-�;LW �E�[�D���3SH���Z�4�C�%�q��(��ƊI�a�SL�K\�,�\�7q���kQ1$�����0@_*R�i��ݰc����#p%�O[ـx�ǻ��$CN��+��h�7M�F0�J��P�p�����h����2\�cwђ���4��::�[�����:
�_�
ZD]��{��/���s�/i��0o]���ɬ!�xFs��*���?���	p]m!=��I�6�;��������r�&�vY*�X�Ԝ�0�}N�|u4R&���6�WfW�>���2�'�� ZY�8��RD+vD�|�0��3{~��(ˠ��aG�؄��ޱ�M+:��s��0vX�t9*�lс�ſ�|�.#��1YZ&�61:�O�	71&ֹ1+��3D���D`�z;�!J�/1���L�=�-���e���ƶ���>Jd�]u��C;�桎?9#�Yϕ���S�7_ ?�A��Aԣȵ��n�%t��\��Y/��wfdie���zivAr�㷥pbq�]Y�<oaʩ��7@E%Oz)Rɹj�|[��6��sZJ��/(�k��`��zas�_o-S���PMYr�e�J T^��V�7A���' �1^W Ǹ���X�s�r��c���Q��������� ��gM	e3����Ϳ;\�|0�G����	��P��ق�-X�iI�
劳<G�����p��S���(�C��ݼ�s�
�hT�Ee��p~���'�0�FW���A�|���mXdT���k���f$��3�+kBK��Ù����%G�}y��:\���x���^�����x*5���x�7���(�\g�.��Ⱦ�6��ۆ����1$'�<B/���:�����w� /}3�z����U�ߜPb�ަ��Tu���PD��n�@p��o����8o ��b��x�|�P���ý��\�r�F��'_��ͽ_����s2�bN�pN�),������o?�P��s2sJ���wn��l�J�Zw�������h�K��,��To?m6�U���d��_$�t"�Z�k2�ٴ4��~,	��X���p�rjulaq�?��6l�LП�߶��CD��\}����4$4��Ψ�H��W������&��`u �2ɲ1�:�1ނw8�JB
!�`�>�B��������$�7xZ$SI������(�ˇ{��/��k��OU9D� ��;�	��'���hi�ޞ&�^m��;�}3���F���Vg�'A��AC��f
��Oir<.�8+f+����y'S��6�~���u�I+��=l����o��(���-����J>�G�B�h^�r.�64y��Б2зڧZ��&�<��<%ߩu"�.ۉ�!� �h(��h��?����Al�`M-�N���"��H3������鱇e�*�����@6�~�X�"��B��É�̓DcNR@���p��C��H!�b��xݡ7ƛ�w@X9�w�q�	dY�c���5-��.�V݉K��T��������F{ѹ�("{Y��El��KH�И!��\kdL�c���o�.]+f>�e�?'��,f{�6[3VC���O)�nZwD*�>-��TwZ?F��'�3��R��H@�����ˑ�E����'+дuC�?خ0���J�Q�Q}j�?tϲ�}Zo�>�プPr߲aj��<҉ٰ'N���D�Fl@J�^2�X)*q��JP�b�e�;�;�%ƒz8��[T����h�`�� ˥p�=��wOY��$��t9GY[�{}�F_����Yg�;�KS5SW�|�:~Q�oG��+o#�Ua.��E<p`P_�a�?���A��5kIb?��R)��Aϊa�h:�bSgQb�B+�>��?�b����Z`�>������R���*��t��a54;Xl�\Y���>)�QU�oa��!�A�=��YФ���O����ɮm���b����사��,�Mc$㛪��	�E"2��/�J�=��(�O�>�6B���wj&``��>�N���Ryb�V���+��md��`\�!�%��tJ�����{��~��p���N�䬤��?e��?�q;U�P_q�����C�/�� ��98�ڔF(��v�I���Up�!�� �,Wf�4�g���,u�.匥(�[�vN8&���ՐklUr-ל�_f�:��jhW���d�n��Ц�/�f��4��#�!X�����k3�[�T�vX�J�Xb����Q�1Mng��<��o'�P���e��xV�UCސ��8�mKѤձ�ұs��I�olT� ��L8�u��_���DO:btZ�d�-����4�o�vs�u=��4�s�ʠ1:��A*�"�َ���f���T��*�CQR�D�&�'"�S3T���`;��z�2��R �`(l�O+U�bH��.9p-��n��%������}^P?+��)�s/0�J�KU&��yf5XRb�Mη����Zj ��uWl5CmR%�^�Ҍ�u-�x�L��^�(�yfn����F�DF�s�w�QuJ6���ʎ�Y�ծ��/+��o��?7S�m���R�:�8�S6��b�#��됣4�ү��Vs�T��׆7�� �&G@��i)���
�1����H���̋�g�IP��
u�K����_�R�S��C����k҆�Ý�zᔸu|���@D�y����7ÇE)f\�A��wOIr�a><d��:�1�G��Ph3BJ�3����O5��oWA�n��et1%��`G nD=�)�j���M1�Y�x���{ �I�*�̯l\��X�k;��t�]��v#��l��ߝ��w��kQ�gD��k���2�oF���������è�S�,D�)�0�l!�]�!;!0��3�&���9uO���� l�ٓB ����ş؉�w��_EΚ#��Q�6�y�(De��QٍNXu8�%��H�C�&�C���~Ⱦ�kX����Z�����Q�o
o}��4l��~sj����J���V�}�e�1l�f��ईJ���K/�<M,EI���Sw�l��fѭ&\Z�+Ύ�TR��9VXk��}���l�{�C�h��~z���|�U'�¤yr��j��Du)�~Lؙ�n�)0彯+���sY�U��d�ԁ�&���H�4��2�r	�]�f�gkL ��
�y��/b�8�nU��n=8A�橃�*��=�͞��j����ze`o�UZ2���Ԡ�~→�B������Z�֕�QW���+���ke�BK*��rCn���2�𿍕ߙReOՂua�zZ*�g+A�\���=#W�L�d�R����hI!qq���Ae�r�=|��$P���=�盉�꟬ϔ�nnB���s̡�0���S����Dcm���9n#����|�QM �-#�x�>\Z�Tѯ{g��r}�uE�4}�Ƞ�Q�*��ŷ>*�Ts�c�ԡ����Gi��@�!�%-�i��-�@b�s\x"��/-�>W	=�:'��l���M�`t�D�馛��X��[z�mj���n�����<
���C�-z���)>�1��#}�]�HzEx��0՘�^�%L.�4e {�׏����zG�.V�%�qFR�6����k���]Os~y�h����9-y�y�7|XqV^�ƿ"s6�g�
�/G�O�hp'�/�6@Wr�l]�r��ExJ;w]s��#�W�n�-y���Q��\���n�]2J�A�&�e��*VW�/�l;a�V��5��IF�>�eƭ����������c�@}
��߽w�A��)�����4b܌��M�n�Zd�e�~��/��@l6*183�&�N�ɠƞ��2����ALZ�B*Aޡׯ���f��(@t)�O:�@i�W��7�o{���b��Հė�~s �v_W`���6P���k)xY���0& �4H���BC��i/�ʆ����<��'舕`�3��m{E����Z^@;_�S>�D���H���u|���	³u�W�ЂF�l� ���hiY6���K�l��qz���A�|Y����tN�☤S�I�7��������G��A�&е�ޣ|��x�k/��'�ϭyN�������)���������N�GV�K���F�WGm_iT�ɜr��\!��w{y��η#��oE�=���p�ԏ$��05�T�n�<v����sBV��й��ݴ��]7��[���'�[�	�ٔ��=��	;'�K=Σ��K3��&���&�>�X����d�d~�1��b�U�V�8�o�H��
Z��nn�<��%�٦��@R�[=Y�2*s�G���n��t
����ʯ�`��7*�t�@�i!��騚��Ɛ���Y0qn`:����2��c�f��:�UJWZj�R�W��*?�K8��wQV�KJܗn�ҩ"A��Y�$���u��m.&����!�-�b�8P�b���e�M�}r3�9\A�p��B�����hTd-�а	���\ѥt����DOSdI��x�%*���0ϒ^�V�f����:���M�5K��oJ�.;�\L})&�zu�$!w�����cs�* y����hΫ�����21Xg\�w�;5F"@7%S��j�yW��~���C� �8p�R͗���h�� ��������f�m�;����r�m�(����^0���an�X��-�����(�R�`�C�~:�����R�;a[�E��ъ��(i�Ā+�KM������$��nK5�Y�Y@��DA��b�f��(5m+[���B������Ƙ�5^�_�WU׷�xq	�m��Z��:X
����%��O�H�
N��R�@�Q]%��S{��hdE��Oha��A�6���� clj�{7�YH���cc�O��Fga1_>*��$�F���_(bР��C�gյm.��YMx����C#]wT��_��v8��59�<��a*g��eƢ"^��y�d�ى�qޓ�&kL[�
�X:��q�o��wWX�c��B��,Pr^��e��hr.���t��D���^om�J%Ҁ�o���o��m��"GTD�q���P���]٫Sۘ�5�� z�v�=��s[�tɳ�v��n�n׸L@)	c�z�����)�3�j�8
i���Z�if����-e��p��$6yu}���	�P�rpמ���'�2�m��R�b~���[t��n��)B>7�dRSj{��Gϲ��(��x5M�3k8��G�ҒSv`9��v��]�F�Kc����
a)Hm"8vt����&�w_	�Ԗ�x�!�'%� �U��4��Z�A�D^���Q�a��@,l������+�8֩�ߔ6	$�G��"L��*|����+�� �q�d"���	淚S�s���D涚��n���6����ǐ�J�d��ۻ*�$�ʎc�]-X�-�.I�'q3U������|N|2p�`\H���ϵ���!��l�Xl�_]��{'�e�p�g��Pfa��,�p��*1#�/�Y?���I��S?e4��eO�hW��m��g&V�#�:��N��ZV/3��������*\�vP�<�wظ���	�!���y�Rޭ���=�Dݙ,#�P�0�����/��=>5q0B��MЎp
�H%Zc=vq���i����8�T^��m������'�V�Z2���R�u4+	��2f
�J���4Xc;�1,k$ǫX�]�n��\��sh��pC5k����Z@g0:��~pp�vI��}�wn���A�o�Z1I���Y�jԵ�ѡp�V���=������=��@�j�p�We�J|��]loF�aU�����W	C���5�G���
;��y��%U�7�*D�m����'+c_�69*���I�&H̙��9!u�T!w�."�?��|�_�@�~��(�|$ݝ�.���K?_ �Rbe���_�:�����NM1@��� ���Fw�i�UQA�E��������jAv-�\c���7� ���b�~��H42ҋ�5�	D�
�5�1�r�Ϡ��uqou�k	'\c(�B�|����&��ԥvv�۸?��	_g�t�W���h;�1C�o����� ��[��+m�\m ��GX�6��'�E�Cu��x�)6�yh�fz�6w"(I7-T�Gސ=���^Dx�U���V��'Ʃ�I��[�F��a��z�l�G}�;�ߟ�q�<�o�v�L��F	q��T���9n*͋/�i�����p������Q6��d�3�]���ɖ�esx�EG�`@І%aU��L��YKcv[�.�,���1���E��{rƲ�96��|�!��,�����?e1�AQ?h�Q��I�����%� �W+ ,�?�3����6	�P��0rs������m4j}�k�l�.5��3!$��I������0q�F���_�>-g�/ٺ{ݍ���*���׋uL9�W7��u�i�j*m�$���<K% =`��v ��\�]���q�i�����
���FO�3oDn]����=���I7Bbq�	9�Ѫ�#��OH4w���ӻ�&��>��`�\�<F)Qv0 �Ke�{���'�C�)ݷ��W�M�Z�����^Q/� �4��ң�������{�¦��CrYζż�lwKA���A��k�31�!�Ng��D�Bu@��9e�e�	S"�k�]�z������&2�G�}�%�o����M�r����s���lIs\��Xgm�WY�sw�
����N��B:L�"I�SEw7��U�\w�Xt�eRA~!���/�Ѡ�7m�?0=�]����ʛ��C*U���Wb>0@a�va���%6�.᫰�J�-1%�����F����E'�k���B�^C��V�d�2`�|h�>��Wݮ��}����`8�M�]#��%��BH������'�d��u��?�BY���V)�Ρ��g��b��ׯ>��TEG�s/�k�VZe<�*J��fIN���|HfZn�ke�rL3�M.;�R�u&�3���V�������ߜ���ԁH�:�,��<�����J�E����m���kβ�3c�?�Ōۋ�6�j�_���?��k"K��4�_���r�����M��f������ȡȳ���щd�4ar�E�M��	kY��LKѯ�J*��Mc+���?XeW�O\�l`1���ߜ_;
Js��N�qJ?-�%C#p��m2�W��Kn�cEq
�<H+�&_���b�7x�.�����Ğ�pU%2�c�ܾ6��^C,�?��R��]��g�tJ���8�\�{==S��& 2�Jho�P]MQD�m���t?�?�G�Hn�R��))ʾ�U�]f�t�<�i�i+=f9�<���ky�w��w��3?`�_����oU��v	�RJ4�`�8ݻ���kJj^δѣs{$�t��Ee~E��
M�W���r��p#9�-��A�,ŝX.I��;��&��g�N'8@�3��f+y��`�������)|*p���܉ 1͈�����;m���w�[
��홵� �&�~E�_��%��c��S�0���e�.n01�V?AD�D����C'\TO��9d?d���o�锓�3�!�5���R����у��H�q/1k������?��������v��_Ŝe^�q��}~}Gr٣�W�( /��1�0�]�E~��V�r�|Z�s#h���e=N9��$�|�5� jJ#��Z��&h���o섻�g��./�)�l��h���ml%�?�}�������O$�w*x��h�0&5W����Y|��Qf����EcY�a�8��@��G��)��C�m�0�w+�KaB>��|ä�y� �B�����,��$e�9�Yٲ�bA��x��e��.�Fօ�s}�����|�;�^�e�� #����`��������%w��/28nDT���N޲;�.|����YO��<�³�2v}�	�HC�K�+��cc�hg�%���S�f�B�{av�s5.؉4	��v����cӗcW�;��Ŋ ܪ`��#��d-���d(C�/5$y,����Ӥ(Tfq]S׮��^C-�}��  �[6]�k��ư_O3��R��Z���fB�.�5���\����T0<5�S�m�c��w�mI;c�,�@���� Y�ޏ�;��f}5�c�h#���>�C�j����d ���L�&�{Wl��fK�u���	;�Ջǹ��4[�PF����V,�V�bXI��P`�KP��-��H%�B�*oy�����3���V�kR��U{���5�@�����4S�`.1H4��>�Z�p6,��㖋H����so���`j�QO�"n=���h� ��Vj8��������$Ҟ�3���M��Hk���{k'��A�h����u�8F�!�"BN~B�ҡ�v2��ͧ��܏�Gj���r�#04F�n�xK�|��י��n�Z'
ok��e������̚�8V��u�Ģ/s�N�0Fh���1'��ty��:wie#�WIj@7o�
˨���Mj�����[�@f��x��L� ��cN������}&��,���[�(-�t�(%�����ೕ(+�����Q�/RJ.VA�I	�IWj�CP~A�Yt:�oK��4M��p20}6 b�} �ۏ��u]��l��pHLk�.�RԢ�Ft����(�^%'��{D+6�WHA�3�K&���:���y�Cs������[�Ń�΄�D�ݡwg���5�i�#l0���K1K��}E�yOc�dyY�{5�	([΄��˭��� �,�7��������~N����g?h�C?w��d���LH��w���؁�k��(ФVݓC���G���Wº�زVԺ~-�C���Ǆ���w�1�hnt�g�|K=��lڸ{��U^@�=}=yֻ��������6���;��]�-ı5���x���a��@{��';�J��L���Ddx�\���Q�ӿ&Jm����B?a�2�C'��7�zQ��+(	�U��?��b�a���N�|M+��!��"2�/�ԧ�3�q娫͓�ԕ���V��[�������JF��=%h����� $�&GHd�M�6�~2F�L��I�~
�4v�8���%����
�o���1T���8N�龩t�v^>�����'�,�Q��H_R����fk�U1ܚ�L�!�o=Q�՛�u��g�����L"���w$�)��Ztdr(�ia$?o���׽U2�_G_O�0?���~�/�i�;$d;\�	v����[YO$�ő�Nk �-��-���
���F񤘅�v���g�`�v��������%�[���/��i��0;�����aj���(�K�IL�����I��/�g�N�B0fܶ�mW�aY��F,Eh�ژ�O��%��o�2�u,!ϼJ|��f��G/@wo���=��=H�b�
'��>� �/s}�@�E�`���gj 1NtB��+,k����$٢�R�a�rwx�m��3)a=~�??�2#�(�7���V��	�a{�
��I�]��v%�������(��ʏ��*��W�X_0>ٯ	�{\=�Ne�����2�ˇ%B���o�� ��&>i�Usy�O����N��d�� �xb�.�ڎ p�ӆ�?�h��`��&���-;M�瞹�CH3��F���y���fkҴ虢-!=�OA~U!>!�Zs�i.�ǟS�L�·C}���R��(�_��AR/�3C�4�L_i�`jt��'*��N�'�_�LeC�M�ȓ�a%����.��gЇ���n��օ�B"�U[��\{����h��qV	r!F��~"��s/�����+t�w���̽�.���ȓry�>N���:P9m1ǽ��7���+Pe��	2ˊ���A��+؈�?PY�L�n,mj�2Ѯ�L���J����IE�����H\Zơ2����l	@p�8\nb�S*A	43d�	������[?6��&d	5��a�Z��sG�=1�=4G��S��'��d�4��C�K��YH����HvN��&/�5|����"�q�:.fܭi����x�	ۍ���K������Ѡ�!�Z�@�ŀ��}Q����Q�_#��?�L_�;>��]{M99Q����xq�!όhw���7��%Ac��k��j�5�0'�~l�(m�H�ǆ���̇Ḵ#�yz!�M����b�o~���ž6>�n/&S.^7�)�v��:���|��b!���+����F|�
�C+�Z���ϗ��N6	�T�JO�Y�R��/(w��`���?l�pwl��	��eA�Mkd%�a���2��1M}��4W��`ۇc�_��t������k O{# k����N�m>x��u&|��M��ޫT6����{+,d��%�2ðm!��q��=��LȽD��R��>���rj�JQ-�.�p���� �re�9��biH_
j�!8���x:T77���Y�
4k�~}��w�7��?��Oj�ܰ?�@����u%E���s��md����õ��v�2�X�+�tz��L�
��P?�=U4���Sl���m>�m0�������W�F�(�\k��&#xa������*���q�#''�W�����F��Q!��_�<x�*�7
� �m�@GY��/rzK���D�4���%{]ƍ���2�<�]�]����X[�D�Z��'�M�^��CFx����z����`��;;�ӒLɐ�.=\ka+*���-��qA|UW��P"���88>��x�'?'�[�-E: �8g��,t�[��GF����$+�A�`&����ox_sQ��sPgz��=ɭ���_]A����V���� ���Y[ѫ0d�5ײ�]UW̍l���aF�1!u̟�K������ \���C	��a+�Dyuu�i��U}����e;�����Ը��~��j�I�(=GMEZ�#g�ݍ���l���y�H����_�ˆ��j	b����K	�/`E�.�]��`�-����g� ����ݛ�1�{�Z����-�
~̟.�=rt#��r��3�]sHl�ʼ
�y�{K��x�܃j�u�i�P��
�*H���\�nB��J���%i4���Zt��^Ȭ�$��Wz<�K�R��,}G�ٙ���!�M�A�m�-V�_T?��Z ��y}E��撀v���X��Q�Pb�"��{���.�A0�߈X-� �o%����	*8�]��Vy�¦r���Q�5�4����|Ǉ�L�,c[	d�.��P}�$<>��<!�!���	��]�8�&+{-z�u',91&%� 1�b�Ȅ=�	C%�X�9�X�8m�t��ba*�$<�Q��{�Ҏ��Q"��`�R	L�N���	f�����xw�arT�uv~��<I,��V&��g���ctuIrGhԺ�����xx"���ѢX���=Kuq�ʈ�Ѥ��0#E��]j,�?�<jx���m��M��+"����_�����ۙ��6�+�"����db��#܃e�;����^��H�rl��0*O���'Ix�P+n�<��y^۶%���1���גE�j�M�^����#��l��Kv��*��FIF�{Y�k��\c+o��sǒ6.��UꝘ�$�\�mK��<�o*����p������\���c�/���Y�t��z����n�:3 If��fZ���� �+�;fɃ�d����bo��u�P*���Q���[��Kk��=�~	��5#W\���+x��J���V�^ߧF?�#.d�(��9�%�z�����O��6x5��AP�kgbmN�u+y,n�kBa�B-�0�WK�����C�	��ze��G�Ǒ60o?Y^ GVh��;��Mtf�^�,(��D?��z��.�>x��uи�z��7.n��v��=}v�?=�t�0���Wܦ�������J��ϛ<�)#�w]��ֶ8��_H�$�C�\tD�i��(���^΂g�g��n����	#�:l�!����D.������nU�P�5Hmk\���W�b��z�&(�h�g�&ף���⒞�l�BLOّ���͔����;��?�,��I���L$%?�dW�3	�p{ZHl?��+�����v�N��W�8��O�I���9uM�z��
�%�&��T���'<� �(�'@8ňw���,�[��i�2Bٳ��74Y�h�
L������wv����8,}��
��`9��-F#�1t?�v�/Z�/��{G�Q�+,�o�" :���-LgP��ؔ�cK���&�m�q͂hj�3Hy0M�Y4��Ȧ�p��匵���0W��}+�� v��{|�7�j�e���>Fj��r
���|���M!�FՁ��"Q���o^k3���Ƭ��n�_��K��h/���]z�\�|E�-N��BĄ����N�%7�'��0��?]��hvl�z��hL��_S&灐�#�D��SHHŷ5�w��c��!���A}�^���,���J�7���c�z�0[y[�We�"8��B�$y�zL�^��7�&̕�������>Ê���Dx����H�[��3������V*ۋN�j���~8J�}�}��P�u}S��$�~Ҋ���:'�������F�1�@���<���4�,ã���Hގb�Eը|���E�v
[��TcO	l���H\81�:�譾��P�/��h��9K�zb�2\���/MxA���_�
�i �6b��(į)�AeCb�-�����WŔ����	��o�tյ̾�4qm!�e�P�և�r��d8�,uE�  �8�vK��ܵ��1o��&���jY�w�A�1`�Q��Y���a&<�� .;-�FSB5�o�����3��[���	�Vw.v?	�r�'_��;�X3 7��{�igT�vՈ��U��ɆU�G�r�Ȁ.Y�d g/��jI�o� D�4,W�k����	_~OxC3sQ!Ld��I���PT����d�l��q�DJ����9�&7�Kfŉ5�����˰-�`�u�l-��������)� ��k�O����L�>�`�ף�O�A��߹!�P���٧=8Z!59���	YXu!#�q�CxW����Xu.��uG�w��">Rn��F����\T)��|����[�*�p�NY3Iاr��h�T�ޚ̾�E�R�������&�
��� Ǔ|�"���:�n_��yk^Z����)Xp�P^ΡK�?6MZ[<�w�V�����\ݒ�0�P�L<�bχM���-��1�.'\�ًK�W��{��y�L�lN�,1�����q�S~ڞ"�G1
�a���ۦ��>ʯ7�#�j	pd9q<''J���M@���T��:�\`�+��-�h)3Y% l����WS	�}w��0NÖ����ԜL�k��]a�O3�_�Hd}<��U����FuY1U�Kb5/W����k�7��bL���'�Ɋᾥ��r����@l;b�JY[.�?:!A5��YfH����-�Y�0fx&�?�d��~2��\��!Ą����?+|w�@�!J ��Y��@�g�L3�h�WqkQ.	���T�S�#����\?1�n��
�c^��u�8p��8D������5�����\T2�m�3$�yrBp��KE�G>m�	��X(_��B�1�����	u�9Μ
>=������0�ѭ?{XS:bn�f�g���ن���O~%ZU��FR�np��H��#",�������7:�"H��`GO�o^vF:�E�/���׫��'Mf���~,���:�.A�
����P̥�Ta�kP-���n
�����	��c
r����5���-q'��e��[�un\��h�/��� ���K���T��	�[y�Q���{o�*�Z߽`���F�+�P/�-R
2�e���{&�|��9(.]��c�����Ts0�/�y�q�Dм)d7��
Yk���s�^i�p�#���B�M��,g���k��Y�Ynԍ)�;�d�zy����.XK�13���h2tv� �q�t��k�8�M��kY&V�S��<)g�B5豜jЏգ�Q�B|R`H}���:����g�y۱��g=Q�@���0���7��OpF�n�[�����5�d|�]����r��z�#m�]���&�<W�j���:Tw9��q�|���<uŠ�,Ň���O{��o��9KG�V�5��*-�虅碲��{���ӯq�t�-6����*2'��▙�uY��$�$x��<k�/�7S��f����٧���.r��]g�P�L������������W`��?hkr�=G������V~����al\�y��P�uY��(�@�kƷ�8�Hh���M[�8w���uv��	$p��oW���y�6�}�M�����fNįi�֢�Ȁ��\r�f�A�(�Yu�1Yz�e�}
�:�֠ҍϚ�$�ړOD�pAH{/gÞ�G�5H�z#�q�3�;-����^�hƌ.�	�D��H����gy� T���0$1n���t@��զ֩��.���fo`��:"6a��r�l���[3Xb�ٞ��հC䴱�y�`�L�VX&A6�:l=�F�a�UR�}9UYS��?��6N���7�2�V5	��)�i�|� JV'��n 0���0z6*���ŋ?�ʞd|��+�2�v��+�l�a�o#pƇB�d��xF�ui���kڑ��c4Yj:.�=��'�][2�})��}��{�|����L嫮t�}38j_ ��v�� �8���`7)���;���劻���2�ȇb�!M+=)��V�jp��8)��]��Q�\κVz�~8�ѝ��6��=�~�1X���� ��τ�2�O�t{d�4�~IA��3SS6�.WhF�`���=�8ڢ~r����(H���/[����M�A�v�ف��������K��!��b6A�yN����>���Bnfu6�����;�w��"����Mir�n qP�DɮFrc��(�'�]ǯ��ĵ�jʽ�G�m3]�R}Hk]��v�9�S��z?�
��R����-�0��v�CT�tuq��d�E�X����x�����x������.���N�OTx���U(uN'��_�¥ĺ�ĭ�y�ү*q��>���o������Db��GJs|�3�C6����(�n�56U�����6;P�h�"<�l�&�2[׉�1M�1��}�P��[�����5�t?�.�z\�,��Q���Ӫ�J�%�y�D(W�O$er(�(�^n�^���r����A92D`�~�.���(�:�Z���������\t�1Z��r���{~:�
d$R@�� ���Y��pc_���_��C�o�����,���6E��U";����z��D�d�-0�����R%�yۇ������5�}� y��F&=v���E��AC�1��-���c,�� ��q5'�q�/�^}/>�h����
��$�u��i���"���0z4�������fS<�H�)� 9'�ϕ�1c��Zz��#G�m�#-pT�2���1�니=��ڢBU�f8Z�6���s�l��*�׋Hh�b�(UW��6�qJv��K`���ݟ��iu�V�땿���?�@�a�:L~H4-;�#@����tx��l8L�7<�� D��\Z ��E��^��־̜��$�_*�u�sy��Ē��j�$o4���ۗ��y
��GKe*O<J`�o]���l ]R��Q�v ��ѐ��6��X��E�t�6�]�<���*-m�D\l��]Qݎ�C�7k2��׼�D�K�P��U}��Ѽ�Ok!
{o M��uog�l��m*�«b	���O��w�=̀������/�����H�8�����M��pc�����|vqǁX�2��ǥ��(ـ�ح���́������'�y�c�\�&G�#b�@g��ثZ7��UT�t �f�|��0��D�T%5���ʝ%�"[-�}����	>0�����1�%i�L@+�L�36f�{�e�B�/t"��#"Pm]���Ov�>����~���Я7�'YI�nO@��{����0B�M�W�d���*����!��D#{���cJ��z������ԥ��9nԇi�ǃl�e���R��2�a����*z.��k�<Q����ϣ4ӽ���]�&��"e]kH��t�m(|c�CV�J7��||�a�5�zo���hoLy�'��-S�#���g�*y�@�t�7M���=S|�nq��=J#��~Up͛�/�6�����b�SpcI3hA�ȼN�l�H��<�����Y���cI<�ù/�h� ���T]�1D;PT�RC�_����iՐ�1�X+ �wwVw.����l���<�����sAr�3����8�B���JpĴ���K<�p�hb»k��t���<y�����Hw2ϩ��(�	�}ߋء�1����LZ�v}�{
�n%Tgu�Ч?��@�q�,̜d;�(����X�Q�Iӈ(B�.�Ysط((� 
!�`�F`��h��"�pe]}��k����N� @-.$��Nb�NL�"{�ø���e")���͘j$����������n��6�Q��t�HQ���	�@���îS�-�@I��9ݩ��xl�Z�o䄡��:��4I.Ӛ�@��!�Au��γD��/�̂1 >o�H�r���A�Ȁ����Eto�( �o�*ы�\����k[�~��Ϝ)�7���R�����?���(�B��#�E3 ^��W��B%��>�����ۺo�PᤣX+�#���t�[-���?�Z�F>J"����:�Gm��o�������F��� �k4�%�>��rj���F��fGod��dYx^ֺ���`�:ưv*n ��6��a%t7.z�;r��8���E2���{?m������[��s�.Xb�+VV�ĔZ�k������~�*�ϽSQQ����`��cL���8�W������+]J?ն�#�>�1a�Vʆ���A��M��b�(�;�o��+�DA1�7�*G'���Z�kd��Sh��V�
�m���:�=�=&`�*�cR9�.���{���g�6\�%��+?|�����wR̀�HSA昫��E0y$)��J4,5V���3c�\	�-�����>ɱ�\gV'{d�tξK^���W����r֗�	�ϊ_g��*�ɝ
ڕ�h�_���6<>���ݫ�\C��"A���"yG\pgY�N���)|Vj��ɢ2�1����wL=%��ԝە_��1pu@�؊I���N�~1�}?
�(�����2χ������n[�ʏ8Ɯt����cE�(�U6p�k��lR�wF�U�e�&@�N�E�F���y{��t��Pw[;���S\ЈadX�s3��h��Z/L�ኤ���-���8]����=��N��< 3|������F�9\+z�s�)�s˗�o�x�D�R���_��i� $�ؗy�u����$����ɝ�
�RgdҺ:3��nQ���<�m�Uq��,�(��1 ��m%�މ���8\�\��H�Qs2�1�v����S��������cQqŎ�����FD���9��D�HL���Plٷ�kW�yX�nc���;kg?]z���H��1ʧi�-�ja��Q�d3 X�?���|ȯi�7Ew� ��Q2�U��v�[3�{~�H����⻉'����.}�AZo�|��t�,1D�ےU�x/^���SH�!�v���������6v�N%r�:3+pb�^0���dbT%-�7/�q�K�<ٰ֥�f��c6�4��R��5����"����j,5%��.ѵ�3;
1��tPUx��,�f�2,2[Ƽܙý�s[x�JI��Nю�N�� �]��C�Y�,�[y C��\�����|�:d�rD��x_UT�'��߯5ܡ����@�x.�\.�'�������)�:�:
�^Jc��g4�r��]��V�Z���w�&�A���^!�l5�[
�k����%��ѭ�1^��� ��TM���pw�QFK���|`�z:�2�O(F��N�J��j��o=�q��	�%DZx,�0���r{ZD`�3�O&�(1�/G��4������م&jf֚�6	��z��<ļ�L�W��@�����ͩM��=�vNx܅�1�o7�\���j��e�ݳ����K��-�Kٰ��@����G�VPnT�k?�i�ʚ�^2�d8�����XD�C�7T}-#��(h�U�x�]d7���9�<�:�q�"����)i�ʡ�����#���F����i���]�g����EU�*���{ǽ���g�{�[	�{7n� �Gb�jI���X�g����Yl4(�;g�����<[4�̮�1�hTH�]��_����7gw�0M���UݕB�EIa��j-X�����yH�\�2\�]^�h���K)fK=��<5��cF=!F���td�i�[P��$��5Ó���2�l���p�j�w�� ?�� /;�s�p�bA���Fu<|O��Lu�E��X��c�QN~����ft��"��!�M[��҃�vkۢ�#ƬI��2qi��*�9J�z]��lu�rрG�US?��ˌ�B�u���Q��]�zfs�Rj�2�;�9)�1:Ǹ)�͸�l�u>�<�����K?I!�r!3EͰ��x\<o��X���cB����Ԕ'Sݏ ���o%�W=��Rp]��!-�n�{#�6���Z�t&�'%�1e���*,�fu�'���L�����x=S��Z�Ծ~�<I��������S��=� �E�fc����^�J�ž�]c�'����5�����BZV��z�����^r��iT�<,"�+´�^8���ʽ0�5���_�v9o��I�-��Q�/��9�qj�8	cog��i�׳Y&6�Aw"��Z���{��>Pt�_:�s��{�M ��<BՅ닞A�V/׿ߵ�1������e�BE�;Ѝ)Q;R��G��br�����a9�\ź7��TVb��vTV����*W(�x\52�/չ�j�,1}hι:�k�/�/�
�ԓ��B�/|[��Fx���2�؛d�bR�Ш^\����϶��!{9���|�����C��]����U��NVG{�s���Z�����o8�8�U:���@𞶊(Y&�&���·NJS���Į��C��,|�r%�c�)���?͚��H������ۦ�>�����\��c�3x�;�ɆCO��4�sŐ!����*:�T����y��+�^�.XR�ֆF��]��\$ah��f���cF��ěa��#������S�,���E���."q�L�P���f�Mj]� 7$���ן훃:��+�J=.�g��)d>�{5x6�C^����	;�4;>1���k���m�m���w���]��)��SI"An�T��j�;�����J&�^��[�6e�)��T������'���,�,���N����օ8�˶G`��D6C��uջJnAc�W�	�)fՔ�vA\�~�X��`��m{Ս�L�1��՛B?��	�Fbd*��Q�Cc*�?�ք����#�p����"�s�]�O=D�.0m�w��=.�����DM����Bb+������-��9÷"M��y�Ds�Tn�N�a�W��A���J�n�x��)o,��� ����HO����ͷ<��&vr�.h-;�������a:<�($��]����ˊyh��hjՍ,��Z_i�{�R2B�bcM=���Lyq[YJ�O"�-~L�I�d��p	��6T�9�����#N�:�r\���R�~[ޟ���?Z��.kH�Z��#��,�ذگ����HBu��L���
m�\7�����]:�7$�*�h���H�2�!s9�[G����"�v�\����d�XR���r�Ak���o���Ӡ&�# G9��-���?�lYW��4c$�[��2vqHv-�C�x���w�qz`�)���':��0�!t�#jizC^F���=P�t8-DG����0�" �L �R . �
h�vx��GY´$�ۚ�߸k���5e�^.�������J�k���»�C�v�2��>ut��n�U6�����CĢ�#��H&VȮ��V�����7�0ڌx��F:7>��%���ƾ_��8$��)?�FI5���f�K���X�L`0k���sa�]�lbC���z�kZcl��b�	5�f��ݺ�@��|&O?��֤Ƚ���m�Nx|��d��"��o����R�u�ak_`a��ώZu���ԷN����5�e�W��m@p�S޳ڨ���R-U��Z3��o�R,��p�Zr�#�q�����2�n8+�_O����ͣ�j���H�� �G2t�1�DZ�)�e�#��f+G�V	_��#��c>�HH��s���V	��}v�V~�\���v�4�a��+��v}������`_T*��R�D�@9��دL�zv�/�4����Vk�C""Y&7 %�#Dj0e�X��s�q�+�����%��4�wb5��CMp�NR��S�TK�5dV�6
�ehQd�s�G�5����y!.ûu�5���52gy���f��L��� ��/�qfWL�\hau����r�Q���\7�L� t.l)�sn�/�J���%t�y�%�z(M�����qLn�JD���!��dB�S	��
�(�0jEN�ɑm Ыݞn��GJic�	��OV����Ӛ�@G�a�Ϫ�ψ%�t�=f1���˂O��)��DnC~����&���V����i�GJ��UXt�"�#vYR����{;IXܺHDk�Ӕ(����Q.mP7�Ѯ\�o���j��z\4T�p�� Z�3_HD� �Yp�
�c��WD�2��d�]Yut!�%b���-XjO��F`h��y��7eF����Un! "�Ujj�#�:,��V��"�L~3UǗ�cа�=�ϙ��8�`��N_a�� �Kf�>(��.�l�_�h:�[nA��)�s{{K`����@��� �O�b�`�=��SI� ��{�����	��d���aĭ����S���<E��M٤B�O��� ���b�����m�sV���m������m@���fk���:7�@}Y��p�w���2�WM2���Z�c�F����;F�M�bß�������!"Cd� '+ߪ�.��3�a9��7���?�v��=)��W�>)5n�G��4q��������W���9�'�	��)����t4*Zi�]��VӬ|���LOY���޸eଢv%�����䇙�t�$c���,��*}�����䍭���Pφ��~�+yT��cF�ټ���5	���&�2=�i�^���V�%�C�s�O�a���(�qQy�	��QR'Ӌ��MBH�6� �d�e�0�0n�ʝg�U��:��aԚ��('�mt��!��������sa�\�x�-����;u�����r,��^R���#^�U-ٌF��͚8��@ڧ��zy���\G�Nk���aD~�y���a+�B9��~1���8���H3�Sf.�Ţ��NT�2��e>��#�������5H�a��T�4�<�?�J�v��4C!�&�T��\[W|�a{B�$T�k]����
��35
�ҡ٧�S6����"�-u�� 8�3������|ӄn~��LI��`�p�X�w�7E�=���EX�/� �� ��7�J��8C�k�ou�9D_^6r��@K��� �|U������-�-:�v�\�et�c��V{e�"�.5��!?�w|\�I��;b�����ԟ�{�ₑ��L�	�`�&h���y��� �������M�³�Wf�9��GW\)VA�����K�:Nn:a�� �[�E����ȋ�؋��:Ʒ���1{Q����:{=�/����[�1��Xb�0�xDi���6�i5^���v ���W1w' `���qK4t����_ɜ�E1��C��ϭ%Q\h�;aƸp��sFh���_d�����ۅ �d��K!��h���(��ӥ��8>3e�o��Ċ��ȬH)8���ɖ�3�~H��������dVf���+>��Ԝ[���$Q��cǩ��ϛ�aY���@�ΐ-kK��XE��\MH���m��c�C�+���'{!�jys�8G-�@�0a���t;M��/N�tm�?�|S�k����@ޅY������?�Ӣt	s���{jà��6��N�S��F3�թ��)S^�I������H6�������]Q��n�O�`Ϊ�bwJ�S��{�?�mc7�c{�6��Y�&^t��w���q~?!�$?�����8�7��I0�_=�)���۴YǄ�w�����? ��1%��UA�Dgý�������\���1tв�#DY]Tŀ��(q�R�2)5� ��ە���v�~�1V]6�0I�>c	N�NK���Ƴj�� >:�ڇ��^�)�O���!$  ����U"3�i�7a�A	��A����,o:�㉯�B�;�ͅf�vcg�ۇ�p�y��k��R��s�X�{M��%4��li>^iF�m-1N=\��Yi����#O])�2�P"�t����b�Y��/���3:U�g�=�V{�f�}����ͪ�}F�����f�ɰ�\{E���ܨ9���Q�X��o�J6���$��?e%>��W��3�����1��r����/u�JTo��-�zkO�0�O%&c��,�eoj;=e՛��Ѣ�Q�wwL��Z��$�N�Aٝ������r$٢޺�T%�玹�4 �U���X���B;g�ʂ"�9_8�<�A�0�0�^en��j>��Ϭ_�|�ߟ㢔�}�������|w"W��dK���i��4^dߨZ� �,��*+m�r���av��K\n>b������ڱN����kQ�6�T[z���`�9
x��k��ZX���ݶ^��|�;�:���V�L>$��,�Rr�wg�5Y���'j��NZOA��8t陙N�/�yJ���I���Y��B�Y�Q`���*�Ή�z[�fQ�O)��֮�Q�> �h+
�M��c*�Y���#�i���({��[����[�vW.W"�Xe��p�6��q?�4CЫ�4��	�
�=?l.�N��S��5���@lk�ȥ��XR��@2o=#��WH{���O�Z�t��6�,�kڼݵ�P�R�����|E��)�}�����8��� l�1��ķ�]u�S)�f}?��ț0k���ۖ@����?N����0냞���p�nåB��Ȱ������3���$&�Bi����T�>g���ԩab�f�^�j�} CGeU*���c���	<l(����C�e	_��9S#�w����6r��U��!�o4{Q5	Ζ�B%�Ckpm#`�dx�����.:˩�7��(5<��P�.pt":(�(/EWҬU;��<�o�1��-G#�:2̵!j3}�a�ʻ?�!�hq�bS���5��fywP���ck�&>�f(d��Ѳ�䗂�o�4s�D��S-	���k�cE�`q�[�w�#&{���ϖ�-�\g��_��$��������|����B���O�ŞL$! � pn�M�p�����%Ѣ�Ie�Ű�����G�?x	`�W)O/���u�IiHK��n�N)�>�L%�[�|$�G�H4�v�zܗ̮�� Hŋ�����3[���X	��0&ń7ߘ?�����Z��2�S�ߦ-(i�t�6uWq{+Q�Ś����LaԾy�c���^sYt�*~����E]�~=��B1�3G������;��G���� �� �2���޴t��C�����a��p��9�$=7�\�}���gĈ����6pB�[+��s�Q�w�������z��L�~_a�C��1�|C���f�(#^���`Q����û���=]d�Bβ#c���s�5��X�"�j�����c���O��,Х����YX�A_���mhf��b��	�z�y*^�&�!�:�E�(٧@v���W�ɛ`fVC�e�ky	���WpC
��c-ص]�/�OQ�ƽ�^� �F�OO+�k��%�9�j�T��k�,����&��ZF"#��M���?�@udo����D5m�S���k;�'���s���)�.֌r4���@pi�0�	�^�����N�$��귋_�1}�u�� ~�-۽N6r�xQ[�<J���g�S��{[b4�$�mv���B�9J/����Щ�íĲ����<˒A��>c"y�]�u'Ae�*<��R9�=L]ԁ�nEƃ�[|.����lU}���,��1k*�$`lL�@�&����
%�C��#g;��B���n%=�:Vͬ˳�V6��MT(�8�v�����.��p�Wj�`2��`�F'�&�|�D���ē��+F͒X6���N�Қ���Wq�l(��T��F>����-�����Y}n�7���N����g��,�b]�Bc�=9�<7
s>Y�~Qe'�$-ڍJ�s�B�k�},XN)k��9���l}�3Mi̾���p��H����;ihI��@�	����΁J��P:�1�b���k]�%߳�w ����V_��Z�^:á���▔暞���p<�	�q�*�F�� t��2`��&M��h.<'`Z '�:���b9v��%o��`�F�����Q�1X��j�T�j�lYn�Ā��s`�������L�@��
<�ѫ�^�邦˜��u��C4���0����=L��l�[�L�����yî`�H_�Z��=�K��wTSn�U�{��XOE�[���2���2K�*��6$ =�z�`(Cܬ�7��:)���n�g��@���4����4	�=;�u-
k�Da�.w���NZG2�e����<�!9������
�@�cV�_�#b8
�鴶����A�ކh�q?�����)��@��{ �4^�x�Jċ܁,c�`��ov�^��Ӂ�B0����a���n1M�� y��	jhYb#�V�.
���T���9� G��$��kwL-0> ˳:�݆�1.�Y_��'�&���f���W���X�-�_=RvdWU�0?�y�@+<�V�c�	�4%���Cm$�*p��5j����+��L.�-�.A�V3�����#����G��F�z-�HL�!8�L��K�q�0��SbX�]�EhԴ�oo��<�����:���ڃ��n�=R�*�ho��ajA�����@��D. �a�W�4<'�M���k�<���q�$��ԛ���n��7�o�
O���+~u����(�\$[���8������%�{�wک7��G�S�U�!�u�UWS���sS.gN�E*�1;%��󕤦�2KX
� �YR��z�[���-���F�:Q�L�?��(�D{��o��c�,3�D��6�Q�PYm�A��T���Ҕ�M��g:Pe~�6ڣ;�����xрߒ��u���V����$? ua+�P���O�Tl�)�'���[�gt�>k������Uƛ����3c�)�ܿ;��TeҰ�Du	Ļ��n��i��C;�W���[%2 ��'��=؁4M��M�c�����;���>�8/������)S���tH?�4�խ���YE��2~��T]��=5n�_����<�F\�#k�M�rY�U��?am��	$n�Џs��k�Y|���S[��o�w�|�)"nw�񣸱ht��o�e�_1��i�V認F�1��9�&m�pS��'�go/hDe�tAÑ�S��BL��0��e��s���q��%��ca瓑�S�X|T;����U׌��]�_s�q� x=��Cґpk���>��H&��lY1�P:٪�����W�I�'I��c�yl�p���p�:2T`�;;
�ћɞ�t�f����C�ε:v��b��P����ckEA���h�-�_�v�#}�r���qv��b�%৓����1
ed�pi:���0Ґs��D����][�6DSZ��zR%��;`kFј,C�<Xe���c �!BPw�\/^ğ"}Vn����%���lI�A�w��Z�"ڊ�#�n�68�Iz��%�S���iKǭ��2����>&���b/�$�]��.�s����n��o��1z�&����x���֪��t�J�s���s�$�ʸ�M�m2^�J�2��� ����ӕ�P��#9%0��	�O^^/��+&'�<E����>Vd	��������ѹ���u)�B���u�\��T��K�C��ɴ�����<� {_l�J�~>�0�d2���Y�����4�L�	�D�֠]�H��͋-�q�3���=��"5@�Ր�,�	�*Y�fn[=%X)�d�1+рL�v`S�֞��q�E��+O�5��p�i�N�Y+-7 �n�yԈlg`���[Đ�xKf �{D��	H�}�A�`�p�-�f�r���2rE_���nz�%�l�Zdt�3��;���
:4"G{�W���q��i���MW���K�w;5�x�Ҧ!�<���
D| ]GJ���/�T-.�p$��m�{�I3��"���l�oԱ|f�@�Fa7�+=ｖ~n�t+.X�|z��(=xBcF����.a�X̕Ɉ��z��dк�%FU\�tf�VK�Tk�R��;}f�/g�R��%���v�l`���*)��"Rp�E-���� l� yZރ:cW�ȧ�	�vǿg�<����[=�>��_�6��AU޼w���������ߓ2>��*�|��������0���N9 B���k��;��6 �!!�#��je�?(�}[��lX�"��OQY�B��p!��� �с�\��"�����s�	�鴐� T�kΘ'��2�6��Z���6nvdg-oH���A��T�{�~���@p!&����T��F�(���;8�`��o�1D�-�&P�oD���Sl8�m�����>~ص����&M�EHZ^�; �57�D�-�~;ڻ��3o=j�oA�`��!�$����U�bň��~�|/�G��9�/7�֒��)Xsug� 7+}��-J�nG����
h-����K��|F��?Ch�s}�M���X1�A���>U(L�Q9�:�fu2@�R�W�ڵ�Y=�x�[xq�Yw	($8�Sm��$����Q�F������bp��؈�}���V< ܧ&&��۔� ���v�Yܪ(�Q$��@���˷$��j9k.�/��y�?C1g�H�cs��G������#Ʌ�@�-.��	"v����,|��&�Ѻ����un7��m���u��=���zx����t/w�G$�����8�+a���L[ו�s�<�{x����[ճ�T���&�YV`�PP���f��s
��/���ЎB�;���%�Ȅb��;��Hi�RNXq����_�1a�l�~'전�Z�K�+�s��݆�-W��n�����Pn��N#�cSI�飾ǟ�]��&��L����h���F�Gð�^i/k�_�4���Ӭ���T��ރΪ�?N�/.�jϛ�h�".z�
O�D�+7��Dr0m���dQ�	����f�A��^�Ӷ����,��7����RB���ځb$6������PV�sL���d�h{C��3R����0}��	�=�����U3���S�b:#�0]O[����A������AG�SR�`O�ώ����0*f��/N`l?xJ1��S��&�с��Ф��F�ʚ������.�+bE� �ֽ�jJi@ʞ�ԉ2u����$�g����[J������#��HV]|��z��SYZ'.���1�:�P3��}e�0� ��ي�.M�Kl�iB�j���IM��-����~����k
:���"��ʼ��96��&;����W��9o�WJb����d�Vͧ��j���-K�Ѫ�q�8��D�a�)Q�]g��K���A���r98��ní���d����[<CFb%�e�>�9�"[��{8 ��q�璓I���5�mk#�iѤޅ���a��5~RNr���}���Ok�/�����Da�� Q�����h�Wsn�-��a�B4�ʵW��U�r�}����5*��g��5�k�k�<�,pt&[(h\.����Q�$lW(<u�g�DA�D[���Usf�}��&�ne�K�%��QzWmF�˞v�$��=v��N�aE}��F�x)ތ������SS��!�T-��-��鶮|��:�$`��s����k�A��?��r/x��u[\�"��(�2o�Z�� dn�W?�}j��n�.U�;ó�N��о���i�W��(��k��|�X�|�һI!��6S�0DP�Տ�"�oH���g���ĵe~<i��%l�e��>�
��HԥA���ҍ�P(��N���a�f�����,|����4�R=��&��n�Oܕ�u��n/G��G������B��Z%WܞgߎK���|�lx��>��0%���5��NA(��%�A���81�?�g����J� /��[���L�2��S�A����0�ؠI;q/ܰr��\�z1�a�9���y�Eo �4�/��<�N�p��鯕b�0��~��W1�m�n\�����1M�3��Gފ;��ꨀM��<T*\���y�c*�}�^w��v�7�EAo�_ݫb�9�6������ג:s6�I���z�(�ŧ۴~?��9�v�,ݮk*�|��MkŹ�{�dǅ�B{�qG�Eh8�i�p[�l�ұ�\�v�:�넡`�(�A&ݬ�VO�ܳq��(
mw����D��ѓ)���1魺6�&�lk�$���M`���C���z�4
�L�r�~5��peUd�a8#�R�BG�M��d��H�.�������1�`c��L������W�I^F�$^Z��YST��#f��_]*���]"i��$U`�����~([�XՎk5WIP-�M�vyP����<Ywd��
�t��w�0<#�����(����1(%Վ�N!����c�g\�E���q|��-RdŤ� �P�+���!.6T;e�c�Vτ@���ʉ9��GĒ˭��o%c7��%7��WP��ԪW9s�P^���մ����i3�K-� �(�cvr�Cb��W�"���`U2�c�K�.H�{��)o~����2m����k�P�]��7�dUd��h����K:���l�P�o���<���z�H���3k���C���o猋������:��A|��݉=�J��k���Y(3eA�(\S�ZKpM�F�Y�k�*���m'\�ج���zz,̫��DtUA�}�ؘ�	��y�/�v�۸:�R�|q'��u�iך �Z;W����}�8��eR� �����C�:ث��5�E��s�֡�6�
�J�Z�R��?HʵMc��h�u�w���i6�İ���������
f�B��OY��*��4=��C"hߘ#T �����zH�J�� M�hV>IZJ o��\Aћ��9e�}p��WK+�q�*(�.� ���u=K)hI�3�]��1�9D���a�X��L�c�lx������j�}�����*�m��RPB��~ \����%ç/�ku��>�ͱ]a�gW:&H��Z�g�4�A�.�q��=���v���@�	 >���P�"����M�h��[rH�����aFA����{�h̋s�1��la��E���T	V�@���ٯd[:ξ��kˎL��ӽ��E������k���b�v�=_��l�y��Jhx���`�����ν/��΢����o�o0�DX},���3���`"�1Q3���H�d�#l�&`�8/��#�ES�x�0�"�n��ɬ�~�u���l��4fX$s8���4aq�A�R��Q�Z����ƹ�;F$"�+ж�l�d)�R�F}1R�k��vL9]���)2��ׯ�MC:�7�[�CE1d�O=&�}C�i�š��/��UE��Dc)�"CG����$d�/J�H����f�dS��.�]�R���@MS��|S��R43ߛ6���4M��q�K%%�9`H�������-��l�V7�,����ς� ��g��&А~�;õ�1LK�#�r��Ͻ�.	�=(t�~aB�޼�3�{l)�]�0�H�nm|����C/�*Jo˩���7�����M����|����c'�I[~�b�?�?|$o=�������'k�).�.4�|�~s֦�!á���Z�cd讻5x_��b�NZ+���3x�t
4���OY��G�h��cTk@�j
"m��t��4�I��a��ju�r~*��#;-,�BH*�;���.o;�-�/-Ʈ�;���	C���]�C��8��� �����a����
��ɳ�/v�\��ߡ��I�:�FgD�� �2�J�� �v3�''�A�Bs�^cg,��H�@å��-Lj��8e_z�,;�(>���}5� ��rpY��p�(�OPYC�I������F���a��;�r
�}�c�\���m�gͷ�̋��v2�\�e�dA�K��+���R�͵���4tO����]d������x�u~������3�xN�.F�Z����g)k0����e+Y����У�.�� 2i�-���!	�r�p����4xosq���@��j���g����iDVѱ������v��C��L�XR��TȀ̜�R>��E>����K����hA�9�I�P:7���e5v��iQ��hJK=��,Q�d�ˁE�,�_�
�s֤���!S��������߼B-J<�K܁M�y��h�2$b^1iD��4���\��K�zN��ec�S�,���������tJ��I:��8�s�f-�sw�^ef�F��V����aꝺT�]h��� �*��B�p�e�����E���/&���~�7��]ޯv�`���<���0\\�j%װ~������yiHm�fo5Ӧ��*pgMV?�'<�zڀT��xs���8y5�Zl���;�懧`��;r�	��<�r2�-��]��:��N��C7��(��f�x�n�]�2y�(���d�
-�YK)y/XZ�0�X��?�(�>e�a�JV�po�۲G���o��j�����`�`��S˷�Wk���ͩ}������(f���xO�ź�c�H�0SoyԶ楪�s\o?B�@��]Q�Y�~Z���|X6k�M;����m&��,(�Na��W8��Mx���5+����CǳJ����ہE�@r)2�m��Q�1q�N��M.>�/��z�~��{t�69^�s�E!�{&��'	u�#��I6%��!^�C�'�����2��Ο|�����
����F�f����-S4��`�U|��u����C�S!�G�=�v �K���Rd���)C+�=�����)d�h���܂HW�vY1����߭�٤�Y������[ߤ�ښdG;�y(S��&0ڽ���y��3ڲ$̍N��T���cĄ�`��ձO0N7ݥ#��F��3�E<�Ӿ�T'���N-5�4$�jǂ��y�Rm���?y�U���Z&��c�/,o�\�������Z����'["�Zs�!��&����Px������e���Xw�l\��սB*c�/�n3k95��5�vg?��ِ������=#H�뭍�wf���\Am�]� W.�I�Fm�퉼d�so�0��~Y=bv��M�P���A�������u��#����j��r�
��R��>�]@n�X �@�*���������xx����~�Y��=��|?�B�~�������)�ۓ�T��U+X'���󳽭V�S�5�zH
w���
���/Y�'�k�i�.�H!{=�k��Q��y����ߖ���;�8���� �Cj:�D�q!|%�k%
�ٖ!M�!��ӿYs�%�|����y�!"��М���ჭn���j%t��lV&�~�<f����ʏo���P�&J�rlX+�m�)ۄsc�s�?ݽ�\�ߥ/�� ���Ź�@D��o���c�I�B�O��л|��V�+�d��ƒkq��#l��觰�g�4kw��x=�KE���JN���֡�J��`��Vp��4G6�ؙ�E��Ѱv���g=����XL�����[{#���W�����T��V��fՌ��C��iu�<�1��Y�n�}d6\���T�� ���֟�g7�����@�� ;B�DV�v:�T��Zu!��	���lG�?�_І��O�.;lT�o�: S��K�}���F)�M�
�ᄏ;l��!�:P ��ԎH����<�e�f������I�o���k�)�۠��(�t<����k��Fbt'��e��G�@���f��!j���J����Zf�,����n�10A�-U=�9jh��W�����1R%Z��$���A˻pT6�z�{��u�=|'#!L<l�7�����/�p$ID8�����Ʃ�k ~���I��m6�엘 _[l;z��lSس����]2��܁��J��M�yӜ�_F)�ys^��$�'Bԧ@]�*^¾  �밟r��a�(��BAdB �aV��x�h����Cp\@W� л7?��&u��+WXΑ�&��}�s���v��σ|Jm��bP;F��nUO�#@J�p�Ԧ�x*!y�0� ��R���B�'����ֶ|۶$�� �UΎ���F�{FF�Q�T�kM��PY�3�[�u��c_����,��2W>ɨ��d��M�g �N]��wa:A�F-JǚyX8���z7�BR
fN�*��-���<
����J&��Z$Đn���������0v��Γ�i'�S	�}��w����yz�{�r
Ў�B��>�+G'iq�< ͗4o�.X�P��A�Du��7��E��*AM��Ɍ�S��SK̯z6��H����� KSJ��7�T�j�F,�M� ���j�<�Hlب�rx�әh�=�J�����v@�o��Ó	�7��)�7��6���7�ދ�"{�؈Ǣ��!}F����������I(`���o2�D�_z�?1>_�yw$���ŕ���%m�o[�9���bʰ^8���1�B=��w���0$GnӃx75�&��v�N�_����i4�%L���4�a�j���/���2<��w�fWP�cq=e(min���H��"�hQBy�w�7]O7���zؚA�7�n�>,�2�[8��O������Th/!�!��K��괝8�.}e˼�a�.�5�ؗ�ˠ��V䌗���u��5�N�|��>ɶ��F��+��*��''��d=U8�o�*a�`�C"����]} X\t_����J�A�R��ү��`�P���������9M��p��ML�����������XhV��<S�OheC&���Φ�/�W�u��.��xR�ɇ���딛�tu�WE4ep���6��f�|l}q@]YD���Yem��?~Q�
}�J_��˜$�f��׭��.Ж��&���@�p��B��4��bW��n��&�r	>W�,+bVUN�4�x����+�dW]g��E'%�DA]��c��ͧ�U6s���hu����RVO��:S����U�rZx�x�jq!��N9X�UPD�;A&��
QoU\�l������02 ��������=���srt�����2��p��b���{P�zL^��J�����n^!��ҳd����DT�ѓ=�M�B�;�D��R�]Sk���EIF��x�v�8��M��:��^|H�?{���"�E>9i��r�|kr=X��:s�0TƓE%`p"p�/�x�pi,��j�ŒG��D��σ�P����V�|�*`I;cI����a�w �πQm��N�������tyAa�����H9�ǲT����k�M�g*��C��p�LJ��J�b{L������W���yZ��fKD�6��(��K�� `m'���-�u4���6��J޵���:*���1��ᣗ*��j}9u4u�!0h�
�\F�����݈NN���Q�w�H~}���'�����^9�*4�MM�>�{��6���1�-{��dh�0+����K�p�ç��[��n�)F�2��xI�mB���%����e�W���HIo���Jg���f��6iQ7��dw�)��b�a� d���}4�@l�2��ov��-h� `�{�`����-��\�S��Ծ<�����.�\�1�e=���=�FN����W�c��W�> ��9��Zu�)��ia����rc�*V���ai��pe��w����U�L���?�0a��S8r>�5n?�~�Q�����!�e�|���5�dz�l���0�z�f�i��g+}����iN��b��/��𮏜�3�	i�W���'�=����F9��l���������QC��d��6�����T�+�t)����!G��ݗ0@��A_ZB��g��A�ȸ�Ա�F�P��*�`t�FY����A���4)i�z�r�]����܅���@�-d�/7���$�q"�����Q5ps�ci%f4L҂S�(�S"��X>ۃ9�7Bb��Px�b]*K�u�<�l�t�w�0mmiO8Ъ#3i%��#�L�X��._A��Σ�'�"!�צ�� !����\�@��7j��X��P+���Sn2Ox�}z�eҡ��cԽjx]x,gV�@)e'�V�~-�%�;`�}�{��9S.���+���+�|�K ��'_�Ȍ	*����h�Jb$=E
�F�H��5n�+#�(M:Jie�*7�#a=A��n4j{V���̀��6���c}�������6{��C!
�p��ݱ�?���~������c����"1a;�����;���Zy�%��<���zv��M�9�]d�J�>Z�ZJ�&wV�9����N��&a� �V𰹶�JF��&��6�,d|��P4�":�[Yي���%�k���J`?ę������.���K�����J�?~�=7�����B����;����A����s�e��Ǫ *Ғ\�m��!=}f�q���-����!=��L��ăM�g�"?R����DS����i��6β�*19�:�]�j�yX�1�%f'����A��g������|�rbk).4�=O+_<��6��71�����2�N���ot����qZ��t�>na�Ý��tn,����b�v�4�EV_�c % ź��&%��ŝ G��%˯K  <�2��S��n�V̮T/GL�3H�	0�
i6�F���F�G��4����/�~,���w��X���Ś��d#,QEsش��]�ƚ�AZ���P���+���k��|0��b��~��7�b��oT��Q� @�>���s�?5��Ѹ+Hkߊyx�d�6��mk����jܪ��\��%������2$֘��
'	q�D1�W	 �%0�я�Uq�ǅ��&�Y��Z��z��;�z
~�\�3��T"�tr/�omF�h�ì���\˖�ӴY�c	�V����bTw�Nz��{7
����o��مL�_G��3��{�c��|2�)��>�NCW��|���V�"��홓	�_�M�Gt���wC*~{���[/#V����[�{�\?br�������C*�D��ኼ���]ǖ@�.b�j�r�c�+�{	B�E�uhno���(@���k��.u��Ⱦ�3��^��[aa�Eu����������z\$�c���x��CP�B(x���i��8�G�X8"r�'7ք���cZ?ڥ!'Z�"d$ΦA��[�*�-�h����=?L���;/����O�,������3�`��S���VB���D`o���1����xd.�kόE�ޡ����� �aI��X�˔�LX�!Ud=W�m��ɂ�T}�$������2��ޓO"a�K��{/({��vq n�P �l� �#���pp�Ö��*��m�� M#�� E�!������`�H(�92�9�?@E$e%w�l{b�������CM��_k�Yq��[�)5}Vݣ@�l�^[^�� ߋ��Eh��:�j�>^�5��u���<�n��H�	��,�YI��Cq�]$r�ao�3$�+z
���Eu�j<

�� o��3Ugh����>G���3�:��ã�Rߠ����50u�W��]��_�@�c�j3�m#�(g�-gf̀flh&��`���y��������@ke�UEքz�=j�t�Q�x޺�9����y��؋[�I��O�=::0�<[��BAJ^.��dC��,`3�Y��'o[��PmA��\;x�-v��`�|{�j��S�t�1��=S�����2@6ʆ\�/��D�� rO�H��E nkػ��pG�s�f��'�t��J@���/of��:��?�L�I�s�W�<���L�{�˖��۟�.ÞK/.��~[y�j��-5� r�lYu�����3iX��>Y+bXek�u��O�	b^rB"��Ïr5r��t~�bY�Dz�A��<ءu�1;t��6W�co|��kFA'�Z�&��"���ґ�����1J?A���f4��c��P�<���V����|��	}�Ü�ؾ�YT����/��E-��\���%�yd6;���f4Rwr�q�G9�'�y�bC�I ��w�״XM���κi�ǃ�.����At����V3�/3q�ɟ2�G}����A�_^��[�1�)PN���+�9-(Z��[ф%G�怞 ���"0��Y�x��C�̊q;��w`:L�M�#(���)ueePc�.��}�%y�t�Z>�� �H�����473�QyIe
b��e�~�QJ�L���S���8N,�պ�lxך#��^V��y�XJ�����Ϥ��������~�A��<��xЧ�S&v�:7�3F#��Y�	FTA��r�<TZ�Y�ٞY����;��Тh=�c��X�e�¬������<��i@3������D 
�Z{Qk|��|�����2^q|B��nz1�.���(v����|x���ʪ�~Dk>s�+^�C���9\`&hW�q�T�	��Z�Jc�"�s��������w����s/N��}R-�wO2��D�v���k{�ǫ�(~~�Y,a%��]�{��(?���6�0[P�[T��F�*q3�OU��(�'ve���l<iR���2���ՋIJ�'��X���+�7h��U�\鍸��:�T�:�����;*Ɍ{�:<@��� fL�h��c�%(�4��Ĺ�w�s@~m䲉A��9��a��h��`�S�qT���(|���v3�
�oi�[/��޹j9�:~�����f�힄���iF1������),���|E���A�2�����Y�1�flp��`긖��O���kn��F��i"�u��rJ?-����o
�_��|S�MS0k�!�'{��B�\�_����Ҕ���\&:�@3h�E�#_�����+���e��-���͎���OA�a�O�(�G�^�#v�X�z�
��+e�Ys��\��{?V���U��+	0q&��ׄDl!UO`�N�x_��4�����.^i/_b2��%����#pH�c�c�Ǩ�e�����c�s�g��1����B��%�A;wG��H�1B�o2e�B[n���|�i������*�k����83R��#����f�W϶D�A����[ΰ5�d_Cw k���n��#�>34�Kئ�zi�)�g���j�8}I>�e��dv����s��x��֛J���h0`�z����Z\3r:�=�ۘKX@�n���l�8�;�@9>�������5+�5	��ph��=hzM�KC�g'�dh ���+1�|?q(��'�	��}�l�z��o[&��s1g�䧹�KLh�`�S�u���kOs���o�pMu���k��4��ZP�q�.��a��քWpTG%�:�2AM�hy������;Z��� h�<�xS�� 'f�77%AVE�o�f��%�Y�b�^���[��)�gA��#�C{�b֡��nS�o��Q����,�Ⰱrq���S9�sp���W�+��'�����02u�&4�"�.��H ���O��H��t`��d��ND�KЩ.h�?�`@�ٛ?J4��������iN���9b��@F�;�����yR�h��U����X]�k��J�>D����K��f��^E����4\(�]ձh܀�Y�Du��)JneH��$�0��^m}����8�� ?��XV3+�}!��̲A5���M5q)@�ܺI����L!�ì��0�4�uOU�	df�r:US�����]bGn[�<���J�q���[����L_��9�u�g����l�^����~y�s珡�@Im���mx�qf����x�Q��(�ѵ$�`����s.A��<A��^�n D���1�),��[9�p4�������a=Sh�CҎ#ÈJv�?����!U��,�h����3mP�lFd�	�˃;rn{OZ��N`[��ہ����1Jn�t���v6H��	�^��|w�p5I���T)�2���!y�C㿃�}j<�L�l�m�(��8�#�i�0���^���W~�N7�۶� "��I ί�{�|�Ry0g^�r+(�h$<�8�&a4�v�9�˵��Wrg�DFU�o)�,���@u᪤z�q��Y��Iؐ��Ϛ�^�Wq�sSi������&/���T�M2D�4�V���HU+������Z:RQ��짯%*���c}�!a3���u�m�]�Q���>�rз@	�����c��xHS�{�FqR]���I�3�,zr=у�2����KQJ}B����|�d�zX�6�"p�b)���F*]��L��0��+�]�h[��N�JW<tōN�i���
S��>AG�
�nH5��翼�����`���&���L��`���io�n�q힭��S�VL� VUf%�j�kȉ�֯b��sW�W�_ E�E�G��IS����:j�]�0m�u��Z����#�ih������v�PI��	NՍ75f{��.�a$u�[&|<2`tґ�H��a��5R7�����'�Z7ԛ྽��̅p��!�>�w��.	���|��S�<v�9;�G5��r�d��|Up�v���>��Eh�@^��7�谭�@Q�O��	wh�A
z���
�w�r�\q��4(���E��u�)��)�n1��^T�K���@��P�^Gb1_�U���s��W��Ӻf��l�9o�ϊ,�;�Q��TnWO�bG��%C#(���Qh�";��
����`(\�ս�
�����8#���ڨD������ ��u�y�>���E��
��5��Jm���jj�o���,!s��m��x�@�4a�ܤP��IY2�l- �Ճ\E��3�Zo%iV]�2 �=�����Pb�sϢF5��6;�t���<O�V���<��	Mֹ~{��>��FI�4�)ҿn�7-s>����f�h<2h3p�5Rj�)�+~�g�Ⱥ���rB��G�LA^��-�������O��)7[�T7�P_C�(��UYp�2�d j�`yS��S�Q��{�+�<�YIg��2L��6	}�)�3���Lol�RI�AĎW��,���J��ݵ0��S<8�9C~ژ��w_�
x�������9�ӍA}6��D'g���������ޢ�g��A&���� ��p�	L	�� �w���󅕂��ū���o�ja�xp���������#S��i��f�S���l������u۲��FQ��ܷ�A>�>�Joh�q�� �1;�F���l�;fg"v�!�#�-���@�`9	1����K'��lqѢ~�W�կ���]w��裡B:�J�Ь��4����UI�&}�<�qe������+q��	�2�i~0��<��n2S��:b�Z�JqT`t)O,(H�t�e���]�:C'�ݧ%�@� u[��l���a��2�t�� �������a�3R�|��g�4�b�Z(E��gĮ���[YIb��gK�&�^,]Y�.}���Dkůk>Y�d���1	Cv�Յ���U�R-f��\�@ai��ZL1�9P_�S�e�N��3e��&I����;�S�⢸�<�ad�f�߹�+��݂1ǧ���9�[��S��X�Ub���;���@�\d��v�dX�ևov3kn
��ٓ|��G='?�.e|4�wvz�I�\w_IBG��h߱,0�o!4�"1�Y��A��}ƪ�F;���ؙ�gcD�U��~��~[d͵Q'��f��gY�ђ��B�Q����a�ur$:Y޸�>_�"&��:�	B�tVWv�b����"�	����Z�L��;�b����&ro�p�/#<H 8��N���{�Q�\���u��D�(q��`��f�B��Z��=M���<�vK�m�p��e�;���S689Bp+�C�!�hT��R=��
r�O�]�P��u?��ړ�_�cp"#�B�Y��� ��a��^�I��,ꞣ��W%'Yo�vw�qj��G�Li��fB�w2W��a�s��I���jf>��׋�"1��`-M
�BɄ�?��ߜJ�SO�C�YD��w���j�&���(�a��T4p��i-@i��-;D;�(XE
�Q&�x�[�3H�k��|Lj��p�oDa�y� ۡV��4��I>1Uxv�Oq~�Y�Y��bD�ܮ�t:@�D���32��[,��o��Pҗ�(����$��6	0S�QA����(����a@���ӌI6�,Ζ=�y��5�ǌ�^K�?;t�|Xl�C� 2��%�F��������mP�o�X�Ŏ�B5-��%�Q�qt��喕�ݯ�{�k�X�t�k���+�<ӵ�¼s�.�=���#mo��&��X��� �nI��n[d��͘Z���M|;�(��@=ػ�/��>h����k��̉�H`�"Z���5��b3=� e������F���OG\-��ǖG��Eq�x5�E�ol����Y��o5�ee�#�c�W qW��"R��@��~̹����U�t��l�<�<'S������2�0�/#��[{�:���TM�F�~���O��v�Pnat�����-c<��a)���\G<�)��gh��v�&N1�6�Ӭbõ���<i`j&cA�z �gA�[��w��=��vQ�8����V1��U�eu�uliQa�Ho��L3�����H}���V�CʌuI��P1��,@1���44�w�d�|���������[���	K>!	�^"k���f��c���T�	G(:D;��j���zX�Bj���I)�?}^��
D���,Ͻ��B7��mV�m���m
��c`Y���,|l�D%��~;��m��T${��"�}��(n�0��X��E4��<�P@�W��J�u-����;�|~ǞS��\�����o2'g�\1�x���o�Pl��v=�Ec��][r%vty+��}��9�� p� K}5�B?e�%M|�s6uѶ'	4#k���PŬ��&���03��p$���}+h}�W�*�]����pF���:	j�X{S���>��8;՟����ʚ��=�m*�X�'	W�q�����;������"<�*b����lM�*8U�Ȗk��;�]�r�߳w6����U�!��l�t�L!Iz��6kU ����1�C#��J��T��8��2/��F�@�B ����FukFx۝�'#�{�;9���%��_H(M�_Lm'#k6>�g&H����D���Q�XW#�4��Ŗ� �p6^v�<J��kO�h�u9+p"�2g�Q[�+R��~i�b-X��f�=C�>�v���ǿ`�ujU� ��i.�ҩv��A/xN}s�7X����~ pʦe�,����U��j��5RɩNr��ρ��i�������e���,�"�X|�����;��`�0��=h�"a���m�a�hq	�x�-�/���i2���2m�B����_�^����$����BZd2ڝ�((Ș������ہ�/]�k�׵U��ٿ�����[�s��ꕛ�Z?�ƒ]����	Y��P�
���qID��qb~���z³�^���9����ڨ<�����5���h���[��#�ѫY�2�1�]�m�c�f�����_����� ��Odo7��-�*���#�.���G��.�0�J��E6.��� +xM����0��Xw��W�4H�K��(���]k�8���N�ɣ�e�����U@���Y�4�2	=1{\�ȀVM`�ǳ/���&�����$��2��	'
�T���l9�����>?���hY�X���&��	�c~7;E�	���Z���\2�
D������4	�	Ԃ�{��E�R���jBe������up i@���2'���t�gv�Z�f�W��T�����LW~���E��;����O��t�FQҾ��k@�o]�J|?�,8�c|�y�:0+��<�R���ۛ�nc2�K�����,Kg��JJ^\� �@H&�jF�������P}���Ձ@4�	)K�ϱ��'�KV�<�dqOCSP���<@�D�}���0��B�n`@��0M_��o������e���>I�h kz[BHhf���c�V_���J4ɞ*D���Yj]�_(i�����I3e��oP7�m���b㞈�J7y�^� ^�x��X�Δ��>��0���h`�
�űj��fs��(�GUt(�M�f��5������)q���Zi�DS�v}�`�)��%����/�{�vf?�ɕ�H*�$�%>d%����*��.�?T�^EP��:�,�]�@�P4�u�jB�C.s �������4��&%	���ƃ/~)����^ ��."a~{���v��>���q���Xw]~:�h��4g�t.�Ma1�3�Q�+r��&콛Z�V���NlI�Rz��7k�)Hx:/h���Y;/�ir�<0C���8���Ȑ��2NQ�n�۩�҃�>���u'�qso��( 2�oȔ��H��M�����I�~H(L���/?�x:�Zо�8�;}�ƅ��n�A{���虡�u��T��#Z�{?���V��ԓ�2Q�D�7gE��GM!���R {�O��@<���x�I����v��<CNr\ڐU	m
*"+�^�s�d-���83ҷ$� u��<w��
4�(خX��7��͵����9X�Qѕt�`�݈�<�,�s���N�1���Ȣ�H�P�������n /�j�8`0Sҷ~#�O������9���˓ևa$�!���HDDǶK:����7������+�l��7hסnVQ�T�KE	�͆m�up�jYi���]�S�>|;�C�K���(,K��{��b����Y�c65�=�p��ԝ�*�
tQ:�ޜ�����sF��q*�ӌڌ����x��2";�� ���2��-���w19gg1#1�8�%⚐�M�6'5�!�*T&��Z�;~��3Ʀ�!�u�������8������d�v���U;�Y�ɜ�V��;p;q����ʴ_�Wdj���q��D7�(f�Op5/�,��:M�QH;�T��wo9�Ҽ����&(k�:�����Bݡ��#.����_�w_�Z��R�GT���K���K��<���[K�u ��8�p�"�'ί�u�q ����o�}����8Ij^�~�p��L�+?B]#� ��l��P��y��"����)�R�0�8޺���y
ߖH������%�G9�:U��F�v��](� �5{�Z�4�uǧ�̙�[�8��K����˪#C�>�2�U�b���6uGҟ�n_=G2-ڣ(��}�կ���K:��ƍ�ZE����K�`c�o���[�	Z[���ksz��U-< ޯ���#��ͻ�j:�8���+iMZ,TA�����s��xG.��6�~"wq#�C6�D~kEAAr����|���=���b[���6���#^�Z v��op0�r���v�=S�6Z�N�JP��Fj����D6(ugt4�A5 ����'���v[�&��,u#3!=�,;:�'t�ml[�����{2���)b��ʼi��<@��#��P�7f�D�v�2����gFS�=j���gX�0��u��*��.N(�D�F�h���#��i�����1�����[�;Y6�::^���&��Jl����z��8��<��S�#G�LI�k']�"g{�]g{22#^EP6O*Z~*d�u����ň���.p0�Y�t�i�0n�G�5~�(|x'}d��"�e�a�w��ډc��mL0wŵ�x(���)�(��muhO��9@������~JVabFQ2�������+r�^駻=��6+× 9E�9�ٿ5�_�?�Y��Yh��C�k�_?3>�f��m��)HE�6$��\�����3fWeh�2��L}F�k/~�4�����5�x<�}~�nѬKm�TplA~�H�@�B<��X1���H3k3�O����4^v�<a�ѣwp<_�
���e��k��+F+
�������:��"���zp���$|���!�uLf0��;5��]��4�Rʶ���~�u+�q,^W�0_�6fRg/3˭��.�����h�E��A}�n�:^@ ��}ʍ˻�V��U+���b�
*��&!���Y�����ytX�a>V �
͡gop��w�#��I���J��l�k/s!�K��I3�<3r+�:����������<=3��DW�R�lٓ��q-�Xe�}��2 h<N�҂����~3�Ǖ�!E��c7���#!�-��7B�Ჵ�J �Wd9cǅC,"95}�ͥ�+����%{v���8Tk�Ů���|i!{�o�0sS���	��������A@�Ip(�6���e%�<rP�j��h5WV-[��dE�͜`֞Ռ(Ԭ��|5"�����k:��6NV(���G^E/����mF��ݞ����ăxx���BTL}ӂUF7~��aUB#C�u�e��I,�zt��s8�88[�B=��c��^�z�����`�`k�*��R�Q�(�T���~���Un}A����Pr>�=�O%���*���rU��Ki;#����Q��C��02��1�{:D�e� F3���9*-���񿜏�@���$�OS����7���T�{[���UrN���D�z����(���A�(Aj�+Sn��8���%�)VK�=E�O���5�q���$��m��Z��$$>��!<�2B�,_�l������jj��3/bա+ ߿�mŎ������RA3��`n�?(���8�ͱ?����d�����+x�[%���f^wС�T4,is������º�%����fm:y��&�B�,L� pK=?�#;�5%�~�EL���?���\�>�aVS�lg�nEJAO������y�b,0~5�鞠V�Tݕa^�}Ƚ�8�#d�[���b����+�A��3�>��Q����2"����װn����M���#Pm���c���5Iƶ����N�w�����>��B�i���d.KZ��/ݏ�U��x(��H#�*�u�!�����*�{�iՔ���a;֊K�Q���i5h<� (�x�7����_H{t�o�����3¥Q*c��ne`O|R��D�H�ߥ; �٠V�^��,.�e��fdL�򴔃��
׽����k�ַ��'�^��?�5�
G��r
��o�`&[���(ş{�W�1 ��K�`��+�o�3z�Np�;�]�US�f��T~[b<�"	���<֌���l-9�F����v��3H"�n@:X4[���@(0��h�c}�.�6�Q�P��%	4�-<s�� z������k)=�Jy�"�^t9G�P����3��G��1�� �?3������	�E�ޖ���T��|3����K�w���;��G�$<<8�Llbl/�E��\v�*<�G��M]�Z;gԣ^�#p*dÖ��edZ0o������QV�X�Qh$��l�e>	��bO�b5�\�LLڤ�^����(.p�:�sw6�v�p���v�B���P����}��>��=W��#4ub���@W��d� 7.;2W��F�c:�=O��"�jm}#5&^��Cv]��ѱ�-�P�~[���V��y�ʰDq�å�˞R0],�xk�,��G���$)�Y��%�=^.�;����Q�r�:Ur�V�47� �d*}�}[�(X�\S��QdcB8F�}�)ΪY'�3(M�+r%�*+���y?W� �Tj����!UE
2D���V#�W#�4��(��u]��Jh�Q" {2�p���Rm��)s;M3�@��g��b|ɨ]�F�jk�����A���I/�e��JG�}��h=�}��,��&�����7�;'�ɼ~#�n��=�E�TCM���ר2">.+:U��x	�ޜ��S�(=��u��h�аK���#ݐAC:�tq%�Q�<�"��$�JP�P� "�߫�"{�g ���=��!�_�u:v�x@��I���pڕ,nRP|�w�1�|�x�$k�@sј���E�͆:���zT d�$i���B��8��J��"���|Z�s�˥����5ڍ����]��Mi2���o�t�f !%�qF�<%&vo�ғ��[�g�mP͙����-�%�G`�Y�9�B'�kP���@���0r�/dU��������x�@��fjCi�
�R����)�fP<1I#.졟��G��&J[P-�;B=#h�\}������J-Z4}�� ���s��֭j�N+,�$�ȿ�.�46��KT~�w� kM=04~�� ��&"�:��/����A�q_�.���T3B���	5�t��√ߟ6��ǻUt��B�ΣM�;����$V��Q6B[�5D�bg����q�GO�~E(�U�p�Od �v�;G�l�[�{��jݑ@tu
C$G~xL}~m^844��(b���Tԃ��Ja�;=8���t���$��W^�È��x߬�N��ܠ�$��A����@@H0V?DB
R�J�C�����q��p�J�;'�X׳�&��?�e#���m�T@�w���T�2�C9Z�- �8��e�U��s����N��\(�n ������@G����,q�ֳ���su�՘��#B#��:�C,(]k��i����C���.͸`(�Obli��\Gf���ժ~�}5�y�Rd�E?���!ZL� ���T�cS��5�
�q\��g,�Z?��"��eu���E�.���z�2F2F65iI��P�a�5���oX����L_T^h#�(�d�lMC"ɈW����'f���'n�sP�������Ӈ����p�oc�e!���q鮙,�� �L4�s)&� �kJTd���j���R�����}��*�_+��;KP h�p�����K�"��Lc����[��0=fh���+�o!� ����Оܺm�e'�T�4Y��1��ai��xc�ōZ%�?4\R���OH E��U���8!�@��G�*�mCW���騘t�_*����Y��k���/�Cd�P�6uە���ӈG��ZSB-��gV{X�v���^L�^�^�ߜ���̱Z��	��1n�
��������Yj�HfЯ�y�j����F_�_*n����=1x��?��+�3����h�oJa����3���7-)U���nYq���/S=�,ù�a�+�/��Z��ɸ�T�lk2��y]o�Ih#��C U����f5����O��"�'��|�O*�T�-��	�D�|�%�톜��P^a���{�K-ŖH��Ty�ah2c��}8Ks��l�ɏ-��w=dc���Mlc�AO�9*Ǹ��H��V�`"�Pw�����ω ��ݫ��ǆ?�ŊN˵��H�N��c&�'&�ND��U8�,�cw�عkF!lh^�1r��۰�y h63d��y���ΐlK���]ٮ~56���bq�z;/�d,�j���T�S�Ș��Xg���42w�(+���g%�o���Ԋk%$�l��?���+:�&n�W��!�L����A �I.`��0G�(���?!6��bw���W6�.{l�[x��Y��<��`1�i�^8Ns��[PD�E8�/�xX�0��$��i�+d���'Ї��ۅ�����4>��p�Qt>2����$���b���9�ٲ�D8�����6�ݫBR�����
��w2�:W
�ȕ��/�l�;�j��?�u���wQ��IB�|;�(�F8�~/7���#5��;��s'�a����v0���)v�EН�r��nb��c�9"e!���2`�]�����*K���-�==��:ry��F�?V��`9���0����>h����-#��c��"�{SW�F���w&wR��g��l8��-��M�!�� ���L|�6��|�<���eGB� r}�^U@�-=���|�= ����w�@�5�1P>����u�Q����(���X�\���<6�`.|.�I/Q��މ�k㜦�;=��Z_#=��/H��)�d�Ǝ
��6szB|Ud���G�#4��.�@�xs��zD��h�J�Ԭ��5K��&e<.qZ��Û
��.;&S��(l;�7C���D#��<11�tr� ��)(�ۯx��x�F|�%�MD�Z�2meD��	��#���k�K,�|��C)K=�_�/Aߵ7Z���X%7IPNk*�܊{��NY.,x�<�p2'	w}��v�.J�w ���m�n�mQ��z�0{A���(���j��o�$��3?�G���wz
��$S�#c������#�נ�{q�*8n8a�6A�Q�@x�|@���@��m�n�i��.�^�P�:I�ꐙ����ţ�o��ygrP�7�1��v1 ��cŘ��V�X0�����ޑVY���[N��T�ֆ�w���_��LD�ŁU��LD@o[!��F��U�y�w�����r��m���F�~��b��I�e2����$%�3�a�e���
��*��iz�dfc��#�B
!Z���#�hM}�\�x���t�X���&��sv��,�vk�8De�n�P�j5�ѩ��Β<���e����R�t��&��cە�TR	#�'J>��Zհ��lb��4�Z��i��ֶ��yd��.��������s�ؚ�|.[�F1ڶ�$=&b��F<m�L�{}���d5.��t)�G}��ԑ���%D�.dY�ڪq�G�d�������[�0����*j,�{F� {�����i�$����]Q���BrG9�#�+_�������3�T��@l�m�qd��S���'��/Τ���K�Σ�Sy E�Jſ�E�!����,�Ŝ�,�GɏZ;��C9)�o�2�W�{A�����t� ͒�h�y�L��s�$���R
\�ߺ����'��_Z_QW��8��v�UP��/�h����I�܂J��ՁI�x[r;ܦ��L�����-� Rm�\��)�B����?|����TE����E�J���ȤJ�^���)I����B33廚)��9�C��NB�d�Z`��D}*������s P�G���Al��~� �g}�$��T�����.��-K6�c���T�)����a��w�[@k{5�X&J���P��P�]{y��2Ή:��9� �@M�\,HB~��KX}���;8q@� �Ҭ"j�
�G�TKԜ�̴��f;��v(�m�h�^V_ 3G�Ǐ{1#N�A����í!��Qb~3W{��t3��D��&f�wK�&FN��7�dk�!��!��pg�~A<����$���Z�wt̂`�OZ2��c:�2Cu�+����AF�^�BϙN�'ˊ�T�!�E��W�26�2��#W�x{��k�P6��� �-�3=����q�r����*is!�J=3��f��5�̘���կ����eq� y�Wj�;�R�3I^�2)��i�ϭ�X�J����]�/�G�A�2.���:犌.auq�H���=���X�|�*tINJ}C�W4oӐ�'�\#V�[b#��;�?���ZGA'o�r�:���F:�g2�+�&���L�Ǐ��DoX�|���]6k@/ �>��H������i�pO���9|+��Cv���>in�(q��E��H�ɰc;؈�ѯ��N���Λo��uUK5�3���4x浝�LlC�}�8c�o�f;�ϧ8'Y�US�_��y=4I���l�����:|7�+�����k�A�~� ���B��|��HXݞL��n{���&�X��qb�.Chѳ�q!XV=4M�w��L�wͪ��C~���-�o0Qg�ˢ#�����d�mQ��5	�*�%�3���,�@��x�Ҟ�� ��c�lu���eq>�K��kws�ƙ��o�B#?]��n�������-����!�lD	�*r1gB�����s����W1Xʂ���^�g�i�5�R=݉�����.ժ��.2�Z�M��;?�S�/�P���t�O�V��:�ԟ���q����D�0-��I��)��^������N��I�D�}�Mx��@��0�[�����j��x�ڟ:��� �yA�q��n�3J�ns:�-3��_o�����m�y��q���pf�5FB޷&���
y�����<TL�z�ö�a�f?f//ed���J�tz��i�����E��*����.��ж)�&>��|P���i��e�6
|M1�^dodl9s{���Q�3oS�������OvB�?��ї�y��w&ˬ��)%}�\9a�9l|�˔?3L���k~�����PZ�˳�#���eQ�h0hl���*�Rx����>�`k�2n@:�x��]�X��k*	>�H�D!S]7�DmD��C���߻��-�,7�#T�Y�&ѼԪl�d�	9�z�b5��������y%��������@�ի���4���D�ai���=�S����6haS��4F$��DA�RB�m�i��߬69�_����ebu9c�[���*����7�\f�{�rL��g�n\b 7���o��u��W��6��d0�����@7���w����<"��9d��l�Ε��
�w���q�K�z̔&*�Eu�_S����rg������Mx�AW�)�c(%� ��h}Ɋ���Q�j�.�9|�PB��`}ώ�D������VN`�~��SE���W.��OP|d���3��c�Q�+F�JE/V�y���_q�j������@��Ȩ�;!]�7z�R&�]����K�-�|n��f�ay��J��ȋ�����͙a؄+m��>�	/���w;�W����B�nH)�q��z�oc; ��?�9��9~�ۊ��ɑ��o��ﾒ-�4���x��9�K�XSpD����f4/U������e�սG���1��PI2�,�
뜯�K�11cQx ��-�n�Sa�T8X(H&�8x�LG���	ק# ��O�]��˩��)fM��"��Vs�q�e���X��8̬gv,^ʁNT�{�iU��40��w��I[�q1��-���*�%[�x��+A�̱���"
#�¹�hz_ߝ0���؆�7��js�%JC�h�@�8#d�'7ˠ&j̗ml ?���fӞ��������
���n��fC�z����� 9[�
U�F"�#$Sg�i���*�K��z�AI�}1)\�,���*��;�?����8�}f10�����&9�Kޭ�W��k8�W.E��9�T����Qr�q3�+��<v�'ݵ"����t�6���������`%�_"�)�=�?�������7��\؝o��L=,�uyW�}6��xV��a?��}�0i9�4��@ljل�Bm��	aK'�e�颛����I�4�[S���$���`����
����o��URF'LK�����xO�0N�x��/�1e|Jas�d��%mg���^b�:��~���_~�P0.%I�F�-��&�X��]	��[��" �V�����-ѥ-}�����uqFC>�5�Z�[A��
m{�����4�uZ�@��R�y2���q쿓T�J�3���)M>�i����g�`��ӪW]�3�,����� �����[]��^x�g�g(b��2׊�M�ݙŉ��[K�2�X��0�*�>�U�Zma�`�%��
�R�6b�#jpIy� �Y���He*���E�ϻi�h���2�a�{���yT�v�{���)���h��u��
/�p�4!��7�.$�{��w�	Oj�&��H����q��p�D0�;	j���!��6)9�:�����M���ұ���.��S��%��
ċ�+MR��Μ�����WD5���A�)���ĹG��XVR���Dc��6錅�nr-^���/�]{��� �+��(a� �ki��o��(�֞��A�g�/�Kz�W5 m���,�h��ץ����G�_��_T�`s��YJ�>/w�B&�P���AF��?_��iOW<��&��.ȷs� �Ω:��>���g1�k �U��&�!���\�A���H�2?Yl�j��x�	�LL6h��z@�U_�@� �ύ�9�)���wS�f- �2خ����M���o�XI:���).�] ��BJ8����"N�Rx^|�ϡ_�/�6ف��0?�V��5�AJ'J�Q�Q2���+Z޽�\j:�� 13 ��Zڪ̼o���._=��(�<;{�qC��f�����X�$1.G�\�v?;��<S��Af�-j��ɏ?���[G�N[냸�JM�|Z��u��8j��"J��ȷ���F�a~6G%��ڙ]_d��ְ("[G�νB��-���{�s_ s�X��Z����5�񎞎��^�05J����$]Gu��X�����w!#5wz�;��������)��7���WS�͍ G
=�)"�7�[����/��=ّ?*F���1��2�Pluj���ȝ��]��έ�z�P�~mo�+��Z���;��ԥ!�1��I��K$I���*��l'�#����%�c��T5%E�S� 2�U5��r'�Яrա��um�
�S���o����WD�TW���=1�}�ϠߕNs����߁���/�I)� h�t�W֫��2�S:�+J��̵Db�!�0C����v�Ѳ�O�$��To~�F��yڇ>���pgqJ4���-��>r�m���u��p�m>�{͐w烯$u�ȧRk?�@��ڤ�H1���T��YH0b��٫Ĳ��˴�!I��/;9�Хb:������!/�SOa��i��]�a\j�5�*:X�N�U?�tS��� ��
�@��X&�Ӥ8�Y^�Ёq)��^E���6�n�*^p���r->��eK�_bkdHX
�1��E}ʡ��_�!;O�Ej ���	\���7���b2���^��4@��:e�S�2��+Er$:k����y+{�r5�A��f'B�e+��^%M�II�G�pԱKpA[T{Q_���<�����r	����a�^�?=~�C6Z
q�'31�dR1���z�8��1^$��	�b�$R�@�3���0P�(2�_�އ��vē��Wf�MAm�!�ۘ��v\���Q�nC*���W��X%��P;$���~�L�$��w���=�S��۷�f��f�5^<������mg[a��p8)�\��<%�� �����-�wm#5����K��B�!5�˒|��"�E�����[u��<�INБ7V���|@
X�k��Ǔ�O� g8U,������P�1KE�7.�Cp�rhFc��Ԉ>ciA�O�}����luAz���uVڠ�9���-�ԕ�F�A��	�P 44��d���L���t@��2��\�3��X�`}<��K��;"L���� ��eWu��v�m�ϋ�?%�9%@g{,�ރ��`/�-���R/�TG����r�����(W��<��dK�mz)q��2]�L���vg.��X���P���,� J%�����C������9�o�{��Y*n�ED "�Y^I���!�E�c_״Y�
mJ��'�$����\wύ?	Wj4ҶB�6�?s������屢�o³���{!�/3F�T�ݱ|Jo���H!9�j�W"����	������gQ�E��K�@��{(�5v�XPR�<%��(׭;��]19Hn���+:X��`����=3�+i���ۣ��<�W0 �2tp�i�mR���;�sl��W~��-�H��Ѕ`�p�ܘ���\�C<��t�Ӕ����u:0(��2K9s�]i��?9�;�4�!,��~�[dع޾y�z�����V�i����4�f��f������E��P�똂���mJ�N�q�Vz��2�T <�wѝ�,�������Kg8�'��*ˀ=0���r�@��'NXA�����r�*�*��~�"�#��P@��� ���W�A�M�
2��g�MG�]�i&$�&q��i�B�59�|�e7�8g
t%��aT�օS��$�������S�G\'ԟw�����{EWg7Z;�h�1��A���$�Xđ�̕�%�MЅ�
�;�:��u�)'���k�_k��C��w1ާ8�}�@��=oJJN�jj�)=߳W�y��;hT�W�T�d��O�j/��4��I݃)��Ψ���<��k Oh������}�B�[��<��uD��C�p��S-0Lf�j����Z�F��^_�^K�ɞ�����)\���&BĲ ��'1��ڬ~w>8���q�qX��In��.���i����U�ź�w�]��� CκC��ɡʘ�A��&a �[���+#ȣm�ϖ,v*��
u"�^ �(#�9��OI�d�^:P.a��޲��٧��id��.D.�n�nyA6N%���t7�/���aeoe���Eh���hGOa�p1_2<(MMY�]����8.������s�\G`UQ��8�8]`���]a}��DA�=K^��4R���+�6�˼�EyK�<Og����gƥ0q�͉$b��^�'s;��z��1p '��l̶�I�4���,Z?��8K�y=�B/��.���1���_�w��s��K��-���UAa�UZ+�������� �j��a�Jf����Ş�Px�����Si?&�����Y3�/�<����0V���O� ��DL]�
J�{ط�9d8�[p���*�v��(�sX��A
�X9�&���o�+�M��'}*��qI��L�(�(��8��e��s��ꒈ@�MbC"F�p��
����#%�)����%m��z��\��rK�wZ��L�l)���%���G���X�DU9kɅ������A
k��5�ʆĐ�R�ܘ�r��1�fkt��q(�ꏃ���/$����
[ApX3��y~A��_eJ}���&2��@,�;���j�*bO~h7���':ox��г�[���P�6�ͻ;��E���:jE���z�,-R'��E�N-��q��C�\�����	�Í�!�;D�߆�'�i�l<�;�5E4�֘׉�%��L�^ٺ(%���7f��sՐ	�l��5 �k6�-�y[5n���^H�8����܌x?`$��x��x��9 �RM���[ؖC��5��6���m�^
��b�'"Ù�b��h�=fV��?*�hM�}�����~���(ܾ��qkW<�:��U?�e�!����¾�9�q���zUd����U��b�6T��X+
�R�/��!<�?d�3XX��T��RW{/�~�LW�->.v �k��:��r����xX�B�hH�K�ܝ�o`��kA\wuclƾ�SN�aq_� ��v(ź]���;`B�f�U	�/��ú�}����H��`j˰B�ߪ�T'���jgt5T�Ω��9V?f� �&�h��B��� �˧:<2 2������3 �C�:lA-���0S���Z5����z>�ܟ�M���ϖ��n3�0Ĉ X%���1��2%���73ұZU�(؎�EI�塑���b�'�3Ad����`�#p��^^tp�BH#�	�[��y���@��{�|`	F����sp���32&j�D���T�Q��]'����sI>�P����.*�Α"����U>��px�젩Z$Z���?�}-+F{��)//���~�l�~?�{f��m��u�{r��.{�a��ÀX�57LɊC�/�?�A�mx����S�N����}��/Y%S�&���B��U,<tj��ae�s��V���b;Ft�]ի7O/����'E��ey��ˎ��8H\q4��{Lƥ	A�^�G #u@k��^�3��u�k�]�o`ƃ3^P��|ا+}t*�T���C��O����d۽�Zuv"I'��0+턲<��f�^�N��<�1=��K}YQ1��(8$��:yh5�"���;:��kis��:�Ӈ��:8���kh`��'I�\�ʡ��@y���3��;UNV��F��/P����	h���`�����?>��:<,jĘ�Ӄ:�꾬L��$��B���:����󖏞�مh3sօ��CW�ӜC�R9=�~)��z�ҭ�j:��@�$�*"u>j�>�[�VP*C���vzfԺKȜ�uJ��iЄW�b�M�.L�-��i^��җ耇�.�J��&N{*�Hp��_� �8<S�nA�w�>^��|�f��P��|ڒ�et�By�����>���^����Elp�($��d�?�+�dc����n mE��`u~�5�TkSۭ5U��u�ެ�7�p�T3�T�Ǳ妨��C�����V�:�����z+Q�A��E������Y�|bt�)d��'Kp�5H����3����e�"E�Fh�
qN���dxj�P!ߛ��^�9n3�oi^:�o{
&��	����Bl�Nv9�w~As:'�l�DO!�,xy��q`�ԂFxY�O����>��2����	�q�_��WB��@�}s�C�\��o#=���W)Db�j�^��2IKз�8��ە=}ߙ|�̙�{�r���x��~i�T�yk��"��F#���Ad@�W��0��9��6-I���'.`i�tf5�<�Z4c�[�S!o�p��k"��g���%�l�+l�
�Jס���/OT��hW������ }��A�p�mu{y==dGL�&̠��>!գ�m�&�8��ӽa�bo��v]{c��>lCj�=���j���c���a��,������δC<N��`�J�����Kc��_���yu� �����Nj9A�t���B�W�n@T��
<�-����G�e  �F#իu6�'�?FTL�?Qpw� #��&���ƥ���O��NK�>Tz�ں�q)g����"�i=���ZCޯ�ͦ`���`����Qx���%�i3/�/���hļ0P��l
�����;M�|��'��d�8	Jm����-f���J���V��#b|.�[�(�j����Mei!*���B5亭�!�Vݤ��9��2���t���è���O�+il���w2q�r�{:ٮ�4���`z��Si��x��{��8رUu"X���ڗ�x���d,��o�p��>01P�r#�d��;�����c��?6�O�㧞5mA��<�h
φ�>4kIp/ђ"����vb�ʥ�)��O��!��,�TN�1�'�S�EA`���܉���@�'�G��\z}�T(`c�GST�R~�x0p��j�������.�=Q��S0@$��V��y)����12{��h��J}������y�x�U�����-u���v��	�7 �IE��C����\���g=rU��M����wu�)���-�1ؤ�z��4�%�7-Es�G���}�ּ�Ƞe'`��͑��T�{�1,���/0��i'���3��/)ܯU��8��+r�<�^u��B ��j�Ǿ�c���ۗ�VT�u;�2��^Ǔ���M��Ϛ&�@�4{�I�j����aĄ]<��n㛶��5�s1�u����)9&ζ�a�A{��)��>�d%-�1�o�'�n$��A�0.r�=�p�$W�F�	黕ʙ�,}�h�Ţ�:X��jC?��q��#�PI���xi��r�26���W^$���t����N ��(8ST�s�j��eɎ>+�ח+E7�rϒ��ݩIb4ϵ}�	vh~$a����$g8Ye�yA���:,4�V�Ò���nH�:v=�.>N��E񐙲.썺Vp��Ӥ-��5k�*+rP�o�T���\�b�<�������|N{'��p*@I�(=*�� b����7��8})|�I�aJۮ,;yźZ�Q[�����p>L��H7�G�T����z��/�4U���Ĕ#`q����|�8z��Q�;�zd���{����5� 	s��C��ŕ��$f�^r;�UiX�J6z&#��q��m�䔈Pb�w�$��j��x�Ƚ��g�*YCL���P������� �3�ug蝜H�L�f��ҽ��@��P����$B�+��v�:U�at7��U�B���gAP'���O�޺J�]I�F���S�i���m��k��$���n)m��7�� ����y�t�׋�{�&��|;τ�_���(DnB�19�F?�qT8�}:����1�xd�7��T�T)�O��Wj�U"�'K�}�\.��댄M�����)�O* sO7�<y&7&v�Z��jw'��#�/�i�T�	��$E�����Z�����qYj�)����=�F}`�(K�n����,ʽ���i���M�pn$����T�����ue��-��n;�0-�<��;�����e�P�k�q֢`\�2r�;��VS�rP�6؃�H�K�_����/�6.���<K+�b Ġu�/�p$�Kwf�q�m����4bJ�G^|��F�Q�f~����[��x3�L4�6[����>�V�zy��\�M멑���� ��4v1���&�a�*ݚ?�_�l����kk�!J�*xk��;s�ep^X��� ]�t_�֎&ht��_��-z��Ng�?F����h���M12-�~5��S��H=�L�J�R�=<�z��%��/�K#����з엧����ߥ�]v-y� �4jYEA�8R�WJ�o	:u�O���=�s���dh_�PP�rY��y�I33^��s���78��9/z�PIQttZ5��
~1Iң���#�{�q7���]c!��f|��������/�	���j�̋7�q�P�j��7��m�\-�!�M��Q���M�%LfC�6��$<��Cw��+�RaДw�g�����*��7"w�^�����@�����|��W��Ƅ�Զ���Njcg���-5'W�~�;<�^tMޫ��O��8D�
1�?��D)�iD�{)}"^6m�V{�jE?�-2Ћ����n�`"ӻ��?��C@u}i�[dT���Ö�Ao�O�i�Up�}����Ѯ~0_��gxE�)�WL�b�#�7����,:l6�C����۞�'�j����$h�4ܚ$fB�	>*-?�[XtT�ߏ���g�p����B��,��6 G�
��!O��S��!��s @���I+E5·h�7HX���Vr����NC�ck#�JHެ�3��WR"�J�v�]�����#91���}�[�0�D6�7�]�0���*��R>�,��!qJ��#��`2���w���a����{����z���$&i������Zr�(4~��d�m�g�X�{:A$��N]������_u ?��|1Y�QC\�F[�Y�a�2	͋1�i��e�Q����wvr����&�e~W�>��r����]o��@}2�<���(�!j�9s��jD�7��xY�!�֠u%+�$`ϧ=.�Q-֯���%���Fԗ���`*@��X~�H���a��?7U��Y�W�����p�������L?���x�E&uU�\�S�Gy�3'���H�omh�A�Ymǲ��;y�(PL��	W�	q�X�(�C�w7w��f�r����I��X�Q�4�6_��,��j�'���3��N ,�Rf��w��x'e�+.��M7��6ַTh$��9�_(x�^x�!��Lq����p��2`rN��G��W�}���
��r�g(��M��'5	;�0�L�Q.w��le.t�{�8�Ǭ�(��o�@(��f�m�.=N��
<�����f�B�L�َ���
~u��ȂHN�I��/�	��ߕ������}����|� -�:�l͎6����0�+�Sŝ��$�v�/F'k��vG/�qb��0 ���E�G�B?���o��c�<9*���LPy���d;v�B�3z���ڃ��1[q�v�>�.�l>'�����!��k4$��t�� %���M/GA��nEd�� �~���P�x�pU�A�V<��&���+�@����h}���i,vO�l�OQ�"E�!��3�F�l�6�2�tJ{�����Z���׆`��.�HD��'S
����G�^�R���Ԝ�;;�h��C!�G�c��8�IbS����D��0�tՐH����7aM�-[V��/�O��~d���"m�
s�؄�g�|�Dm�}�~�1�;RF�\�(�M9��i}�8���}��B���n���1��v��yj>�4�*~����X�}�S�ß<,W���7Kh��r�h�p���1)���z��Z���>�[���I��-��&X�&���Q"�r:��������<�+�Lr�s&��{s*t����E�b��`b#)�.%�lw{.G4��"}���]��ڒQ������u ?���Z(A�H�CCxs�z��樏U���.	[e��D��U|!���.$g<���*�a�CT��W���Gf�r1F_�t���*P��XF�1��	Wԙa�xef�}]�:Yl�Ͼ(א��Q̷�[�����3gZ�:��,z��xڄ���aA�!W�y�f�ڣ�~��G�༒��W�%�X֋;]��nSrTs�DE����,é�%x]�Q�
Ǉ*Bb�8����i۱6�~���������+�W�ԱH�?��[�Q��&,���H�H�E!de��SK�5V�Z@��ʹ���[]�2��H�f�k������k�ϱ���4���U��Z(��t~�	�m?l�78�1����檸; ����ll��Т���i�Uk%��^V"=~h`�!$!T�Oc��Q��:H�ӒقN�m��L2����BG��;*��)=0wɔjr��J�6��-�K�l�LX~�B2:��}���k�Y5z�:S�rØ��"��=�1��AF;jeR��~4��.h�4�:�\h�����lF�+w���	]e��5�A�f'/a��L:ƞ���G�×�����v�c��v�O*AE�3{���	�~��	X�4��;�q���`�{W���E��� � T޹�j��)�w�D�t۲�X�3B@���.;V��
�9R�� A����Bg���_�9[z���+�*�Uo#��Z���(�
>k��c���� �|`蘒�A�?=��M�4Xl�W��{	�?%�� -'���x��5h��ݖ��I�@���橚YU|(<� �Y�r��"0�{�ӹc�Z?J1u�n �!�J�M��#��y�\b
�u��y"�D�$t�$>b�#�@l+$W꺶G��T8�@�R��5P��3�;�-Gw�zmx��'�R��|D��=�a��e�;JZ#�K{�~�l~��Ƨ8��e�M�ݹvH�L�W�^��m���y�e�-ڬ�ApG�W�k��;�3�&�$���5��C<f}�����(���2{Z���q�4�0K"?����RRc27 ����e|l���h+���H>�����=F�ڵ������q�S�So�
�5.��r(y���W< ���$Fi���=C�;p��s�Ƞv0���ƛu�v/#_�:(ZX�n��"!6ޱz?���5�U#!z`V��>�[��7c��e������B{X$ŏ���{�[�D�����131]��@q�H{�KU�$	ڮ��y�Ğ�#�B`���&࿥4�b�rO������ά��� �y$Ō��ɚHdc�L��H��Bn�M?I�2�y��eR,�A��4m�lܪ�%�*52�%W���$��S着�?I/Sj%�k��_icWw��cLb)�$�sc*[�@��|�;NL0�$r`�NV���G��K��������z��Ⱥ�>�8\��ŦJ'�a�cy1-b0�Y��&	m,/�JR�("��*�1���[�OX�Q��Ừ�`T�#���;�A�A�*�����k_1�N�>�*�7ڼ~�oo	<��Q��]e�[����J�m{8�Hn���A	}�8ޣw|% �S$����Mq\�I��ӗ?������T�Z*�W���)[!w��|�ʼ�e[��Wu͟S�H�wR��I�U��<��
��}��1��'�1̘���������Ƭt�c$C\�$#�����q)T�r���=5U�n�Gl��:�N);X b�Hm�%�m,˔���>&�ד��yjjN%;���ĩ��"	�9>�{=ܞ����:���J#��OZkŀ����W�G��tц��ىpR_4ES���7��D�S�������0���d:����:I����
���X�����9!���֬-�7 <�|���z�$B�苔"jX:V4�N뾥�N�Z=��@Τ���X�WXlX�|'�o�\"E�&Y
׶�q�$ܤ��N���T���LYd,yV(�M��@��G�A�W�oc%�n�n�b�������ʖQX���7#lD[��*7�)��s0)D�2�tZe�#g�WK��u:�w6�k c� w�_�������ݪ�L6�K@8r�k+
O�b^��T�z�\��g��7����<B
�Y��j���x/����~s �b=ACxDѹT��sv<쳙V�C�h�	q=�)"#��fҫC_n)xF�$b��8�1%��Q]F
�))��y�y�ʩd����,��#����c��s���K%6;��+�Y_E�Ȑ�'h�!A�ax�W����(uFB�`�h�&=K%���
 �7��Ǎl}�H���m>2{:��迠�7�x����^X�������@̔�BgD� g����{�3��V��P|�'G�P�o$}���l3��WH w�;f�ǀ˾h����3��N�BG��g ��3K
շM=xL�V�����ܬ9�\"�}��זEwa ��쭥�җ<,�,�̰�m�]�,>�e#�e�x���U'�rO�o�?j䙡������[~M#l�s��V�ﶉFoc��R�'��!�'��&$KnF�V�6����Z��ڛ���qa" w�P�]>�b[Hk��j�N5�eR��@T���=��wRJ47c[�Y�?;��h�o,p�Y��n�R ��^����:��3�NZ��Rp���_���ښ�x�}�ۗy�`�$Ժ�l�B�T�i��P{S75!�w�I�E=S���[�\�)�
ur3&�����������
�]Ny1n ��G_4�o�(��b�գ!2
�5⠴n�l�ѧ3��/L:1�Y��B���s̻ݪx;ʖ&��G�/�H5���.�  ��e���Rp9�c�	���9r�h���F;��0����$̲��G��=��T"��w	/��C�±��-�Dd<�r�𪠏ݷuh����bֲ?g�~�kt�MV��n�c�
ν�i��ENN���=I�q����҅r��!̵S�"�R���Ox���J���C������H�J#-�+@�yZӡJm��`��&Dв�+�zYg������K\�JύS�!c�MFǞ�hq��
��:�DN�q�e5��x2`���R��C�H,G8i��[auͧ���6�c���(L
��S$�>����p�>ă/�]h���G?�uX�~1Pݦ ���ywNa>��yYp&���ȸ���g�֝ r�N�������rA���L`%��йq��k.ҧ�t�Y����̮T��Op�ݶ�����k7RO��\�����҅׋	�b<
�
b���|^x���\��*�05���+h��!P^]I�.��oZYH)�����I��NW��'��7�Dܹr��*�όW�k��L$�����;��Ā�J;��Ж�����Gj	�B9tU7�ӓEs��lړRƿ���^yMyXqC25H��d,�]��nWdK�\Q`����.�Gű�����%�[���,_f�H�)������z��>�
ק�N�ƊT��rj\XӉ�9��VDI�e��i� %���t��p��ן����
|N�`�/5��E|�d<ұX�ǎ���_)��S���Q��dy���g�k��<g+0�{���?�����s�s�xx�g�����hJ��-r�=\s�U�rlPX�p�P'��n=�_������S��~q8��2�sY&mڂ�1�1Y������0���!-�ПR����G�K�BcІ�[��ﺊ�|QM8�q�s��DB蠹���	ޮ��)B�ݩ{Z@Z��v!y�i&YN���8ȏ��#>�mǵ2�␹����{��}���ꟗ�"W��~)���>.�~���"��KG3�3l-<�Vq}��>|����5�:�kټL�� wu%�?k_(:dG��iۢEX���4_����a�ӊ+�@�A妐<�1/4��n��"�}qؤ��9�3Z_Ts2frM�8C"�YRi�&�U;Q�{��F+Is�7�N鍟�ÙN� �Ƙn1����P��le�?g3�~�X:�5�dX<<��(i�i�	�@Eg�ϡ� �b<t�WQ&��xj9�r54�΅\t}�;#���u����oV�*�����/�Q�reu48�]�kBo��/QَZ+�:iB��/�;�YVbsދ���s\@�d�M[�@�2"s�ԇ��b{�^K�����F�·}���[�@M���>|#��W��K�7�b@|v }�D�v6I �h�T���7m�������g�A�V5�,���D�
Af����$��C���=��ʔ��˷R�:%�D�O8=��Z$F�P}�$/��9�mV%�8<���C|�z>���!9�9�4����.���pF:�T�|��'+�4��E	s��w�Ӧ`���$`��]���gb�{Ø�f�d�������_�q
��1q��|_�F0�G��jxFj��& �+]ɋ��M`�v�$����	w- &Cƣ�t��>����{a�����+��i�R<"��s��S��mZ��63&z?0�z�V|�$��R���O��W#�)��Z"�f���G��T���V���N�/d�E@ք�O�^� Y��ѕ�ʑ�=�(�{ΏrL�)�{Ǜ���J�M���Vh�X���^7	�N�( �����R���	���~�\}R�W��6)N�c�l��l��>���c`)��J�d����\�4��#Z�!&� �C��q-޷�.��N���z��Ǘ.j��Ѝ���Ե.Q�� I���K/�5�y�soկ��� ���1�w������<�zk��7�|@�e�d�M�,s�p�+љ	mT7�r�m� 6��N�c�8vUX'��l�r64��(��fN��C��9z�ݯj��a,�����F]�Pu�YNRbĤ�Z���O��>�>. c��C0ۧ��hζ��о+�L�U&{������5�%~��>�Ø;d�g�hg���F�<񜾿��,�6ݼ��׉j�L�-Do��o\xJu��q���#4k֕�|���:�{Y�c�1��/�0e�<z�HS�7Z�V�r@����'�ÐufZ�#��r�n��ͦ��C��x�aq;o�/�'�{�`��|�A���5���� ,�~�D%,8�K��ۧ� QӾ�E\�|��lTx'����<���ԣ��u�[?�,zr1�w"g/ə[�0�ԁ�U��s�t&\�!>��l˒�[���}??J�|vȂz`6�?�yݭ����
��m{w'�����!�iJV!0�RL�1�r�#���l{����5r� �V�
N:�=	1Ẃ^d��#�1!5g���Ji�g�`ɷ,� $�*6���8�Jm�.[?5�򱖂¨Ad��~B:C� ]����a��Aޓl�u�4;�_�9"N�z�ky�8���ouاDj�Ov�\Y�J�BW�/�\q%�rT�z��Zjƕsˉ
sBĸ�[�G*JƱ�|��yǅ�_ ���\_��F\�\�Ƣ���������C�µ�*�>
�H��`��J�^�Z_�R�:~*��WYL���<�-��&K��6*�10��2�ȏH\k�:�n�\� �%�Ⱦ��lNJ�.�>�$ﺓ"G|�3�Į���$|���V7�^�	P� �cR��mQ�{�NC�ۢ�pw�P���zh�8b�����n��0t9�a��������@}���~Ҩ!f��pk���fH�%�0.ޣ���{�"tٚQUA�紂��ɦ;N�>�*I��e>L��R��75���"�s�B�b@z��>P;]y�)A�a�� ��a��] �EJ�� ��)p�Ր[�ğd=N�}�4� ,XT�NuJ������ۈ�WR�%�ZlT5<�F�*��]c�"o{Bp�OSη��p�軆h$
�DYl�$j�W[��\�w�nw��Ke��}]���TK6��b���~����iP�R���#�$�&Ij�dBE�Vr�βN4�T+��4��~��aa�a�i���m�Y�:�5��)�������*G;J���9��F{����U�V͊p�-�����9­��PZ�;��2*�@
ĸ��!Wp������[CO��4�lH��ِ� ��|�QDlr�Ƕ�&�Ira�ہ�A��s4~���6\"�����6d���<H�8���G�l�J�+��#�B�>�Q�
� �m �τ"�z! � ;[�d \��(�٧+p�]��"�c��Cwf��70�Qe}�����wd�_j>Ca �����B��F��?ݭh)Z`�)ۇWK�&\eTG�N^ ���Hj�.�B��,�'�ϡ���"��XG�'r�$TT�ݮ�K��͢�����O��F��s�yj:x�ʟ���]��s����T���AP�d�f_D��� <����6,�B�״o��F���S�Z�0�����j��K��$ؚ<��x��>I���xi4����P�N�9t�&���d(~��=���A�o1����w���32H�a\��!3��Bī$ /��B�K��ho.}�b�?�\eƪr��.x�x���Z���ʅ\�g�M�%��&��h����z����?఍Sb�km�JW��t|4o�!�rb"�?��� V��K���:.�$^i:��K�V|��7�n��.�Ɍ�D��a�6�z��o*�Zm��]�a+�|�DmK�	!���.�uk.'�m�6`f��;��<�Ë�`s{YM�����\�oڶ��)��2T]
<ִE�L�X�c����h�����m�4lnK�'/A��z��Sk�94��#*��r���+t�5,Bw`�ێuNm� jW��d��Ε) ߊ)��l�{}N�*;�8zD���z�mCb!�0X򬵡0���K�����5H]�H5��d��:ڷP��v������!��沿����ܘk��~k�j�}��S!r��P�=�y�/�n�Sv�T����Pʉ6�FsA�O`+��cv��M���M�� ]�3k9"����YIB�GN�t�}�_��V�·y�ײm�Sk�ެ� hc�r�Y��bpF�zT�ޑTڰ�o��Nz)��{�E^_Ԝn�$B�!Wь�1�P�92�bD�����V?܄2�x<O���i*MA�����)�b6b�h.dD�^�������Q�Mu�������JW�Ƹ%Nb�����4L{�<L�
R��'U��r��Ă[7*�����P
����LY�O3|'�T_!s){P@D�|}WX|aZW���9��A�EP�����*@�$�h�v���诶���'�yO��b8���b5
LTN��O��B��0��n(8>����cF���!J�b�gx���;�}��i�ܻ$�֜Y%�����j^�bdD��U�ٶ ,]_�ޡe�5�m��3�Z����r�j�]��������QMպ	�q�8r� �IS�d���L�<V|�/2�s$�HD'��6�T��b�n��G�0'�4�󧻛l�~�{,2R�Ž� N�H!F������> ����/��q���M�������#}:1Y�K�=��#̷$�n>��)�Z�i�D���I��S%� ��Z��u������&~�����VbU������#���+:Y��n��⍪i�^f-��b*;�'�Xz#&�d�h�f��>��
�g4s�&O�<��~<�o����{�W:����c�Wn��M��@�-��#��t���}�i��=?r�0;�17�L'д���w���:?��~Į��8%�J��c?i���l�����gc.�UXq���;�#{UvW�ܗ��s�o���=�d;��]�+%����&%ہ�,�/�Y��{�"�+���� �	����b������g�W�wa�%������<K����w7g��%#w�=�n_ѵ7�JqrG��k��6�އҪ�*�B�ʮ %�y�V���$wBSq����&��L���R@�/�(�{�Sfb�>ʀ�#�����SfKuX�E(�9�(݀��n6)66=)�6�s�'!<�x~���LV�$��Bն�0���T��x7UZѸ��� �����w%�^��c��g���j)�����u|&��	�hw��K���NpW�^3y�$���m��N��9�;�#%muc�̒��[=���kWؕ��߻�v�R�I�uֱ[��$�H�5E�x��0�9샧�>�t�qti�{�o�gBu��5�d���o�U��/��,[�h`GN�_�e֫�s�`IɤG��2!��*{%*b�K������կ|%��I���r��Ub���`MR�e1� m���<gVX�l��V�_M��u���r喿�6��[uLv]�F��鸡�������K~x�mF�`u�@�.8����i���T�;r���}�*��E�ؖ ���Ytk���#F����y��������*� ��^�ᴹ�����rf
Q��RHt�����jZ�G�n�~����(T�+[0������;D5J����ǚ�k��m��p�q�~���t���o���<4�5�m%?<3��+�c\}�`���'�a�=K��R�c��Y�8���XHu��ȣ�a�� |��Dl�� ΰ_A<���F��/�����#!ZP3�n��6?*_��)��mZo��3FK	`�E��S�|4����7���Ը�����j�e�#i��| ;�hUql��6���-@��%��5����S)w<k����?5�۬@LRVW�g6���4.]<�O��0W^�RP8�� �Ȇ�s����s�z37��dU4�����&tuB{�l�r;��"���g[��Z~
u��BI�p7dK��zg�="�&�=�E�W94���D]�1�q�ҏ0��$�7}���=P<�,��Ǐ8g�(Z﯍'qm�mL�	�����G�u���H��$�(�	ۑ��7�D�:�k5̳Y�n�yd���Q�(�L����ص�«���E�������0|�"��~{��n�*,�S^C`:ji����)թ�6+�2�JH�r�4�U����ɶ���9����|B5C[č��Y��1�x�t�Ѩ� ��_\�i��V�H��M ��z��P�Q>�S��i�U�eݴ(W����*Uѹ���z!9)�0��96{\Y�y� �a�\� ��hu]鍻	嵐o��74�5}���~#�n�t6��jy�,��K4�]��-�ɭ���W�fT��5��u"�L}��SK���KT�� \cS5ޟ��X`Uɸ�v'��6],��r���D����\���um�9�OG|�%����6[�Χ�e��-579[��?#�UM��0{=ŢR9;�
N7��0��+���Ed��@�<g�b������ȷ0��8�Su�5��iy���Z���|��W~J�{xmW��B�{�}���zQ56��jޅ,R�������;��	D�l�}��ಆz]-PRZ7��'Y�YI�@p���]*�,����{�dI��Ǣ����]T��S�fsR+f%�ü�A[�_�o�3v�\,7Κ[ѣ��fIe����#�G����§��(��u�d�ղ]�|���˄G���p�\���2Ȕx���`3v�B�o]5����Z�x��<&���s���PKq�-Yhq��$r7m�].kV�NG�W+��)���� ��P=D�p[�?�����1Q�i�������0w�Q����͘`L��0�8�����as�m�;��V����۔�TG�,]*���$���W;���+��i
��,��$�K��<Y�25h���ɧ�*[O�Y�g�J%�0�=Z�n�)�=��+{���Z�y����1�#�s��zpv��	MV�s�%�D�f{Iq��ĝ)���1�vq[�^�!��ݗ�4X[�>+���gE��w?�\GyS4�^�Gh}b!u�2�>w�ɯʅ˓�����	�M�ȶuϼ��IHY�g�����T{��6�g�� ��8��2��[<`R�����~~���w|R-#�(��ۆ�m�Z6i��u��J+j�#G�Z�;=���!�{�j�������woV����W��o���@�L?�-����:%E��37D�2�t��h<
��6r��A�X����!
KQ=d1�R�D�U����̜`2��Na>�d�&v����պ�}���K��6zJ5��&�d��	�Z�����Ĉ������֠�0�M�D����n����%z�;���J�pR�P8�v���A	��^�C�膂�T��zy���[��Q���>z��8��Z���������]�6��a�4\Lb�D��D@��k�D4�k��z�Bmj@��UM�"���H����"$0����.WN$P5	�,�V�>�P�;D����Z�l�i�"EN�LYO�� 	}1�mUcdp��î����qsVq4��z�!N���w=��
������SF����+;ۨ�br�D�)�3���$H���^ >��Ձ���qq��Ht���'m�U�6I錣�k��K]�vo�pz���6h���2����e�ZM`4S�x{(K��nQ��#���L��w�7Z�"���@~s0lgU�R�+��Ɓ0��fV3�y��U(?.RV���Á�Si޹��	��T�kQ�C�{�*}s����"D�n��~���-'(�A�0Įǻ�,]DM"�EW�k]��m�򍾪S~2\ǔl�@d�̢g�����TM5H��\�7�[
��2��u*�I����x�1\��!�����S�a��Hpqn3�9���������`�5!��N����%wM=�8��yk<�_�JU��V��(p��r�V:��a�$�
�e�2�ƾ�B��-�U��H�0���]eڥ�Ҭ�'A8�����]��F�1WZ��9m-qY�
�>!�:<��bw*S5~ -��MO���@�3+�_;~�P�؀#g��'�뀦�=��`2?Rjd���7�̥����~�0�~(!8	���ĢG�<������biI�q���g�3�&�&��i���[4F[�n_�Ál�v0U�� ��h+P����ul��v�@�(�X�|�Ʈ'^�͔L�~nDƛ�K���8P�B��ֳr�������l��&��H8Ŗ���	�@v��iD��>�}o��!�M�=�xC��YAHcO1�=kH�	�כG�q��������S���u�ݣv�,�aԠ)TJ7� �A���b�NxR��9����&�����r���C��p�Ɂ��%�����gsِ% ���l��XڇAM�wL�凄SD}4�taͮ{��
�(������l�-A͚3$����s{#1��V&S�N Fp�%[L=��Cj�/T>���=���h��.����O�8`�tg��X
�R�%�;9��̤�����E΅)����p��\F���FS��Ǔ?���m����Pyk`���&������X��9�������r�����;^I�6��	�j�ٚߋ.i�
�Y�s�,v8T,pF���u��),3�u�E��쨧���w�!��Pl��)�(�� �*v�=��F�g�g��� O�4[J$2���KKiw�s�h�m~�T2G�y����I�g?�=ZQ��8O��m�Cy늮3s�M+1E$���%:h�����@��Զk뇿[༗�7i�b�M_^Jm�C��m����ݔ~��j�
���0U��&��ۏ�4�{Ɯн���N7�,K�	�Z�ǗUEk���4YF`O�E�E�)�˹b�{��Хئ9�� �pl�� wr�a����t�Ń�Sp-����X�]�����1���fA}�LO�����M��k.�v
�X�[���5LZ�����,T��M^�m�{�P[ɮ�oa���AP`?��Ч��Gb9�\�@S��m��?�
�\NU��������3�#�Ϙ�?}�5�����ֳ�@ع������7i�Pb�ځ{]"ʹ��`��!�~=���`K�e�v��j�uAl���Q�j�l�����o[0������{H��/z
6��a�^��'���宼��lE��g�C�Gg��lb�z�3\�L�pE�_q<9�NCm�F�a	M_���a7S*7!������Ğu(�E�@�<zI�G�ys*�n����D��:�����)�-D���V�{k�굹�@#�f.��z� !h:
�������'C�ƹ	�[��R��DF�y�PGܓS�_-�	��g}��s��
=)v�%�_ڋi(����c��WPHQ��:d���w�-�;���@a$��ф�2V^��2JM�=�3&�y���3i q-c��IJ�=J��ݢ��1����\kxi�y"��Վ���O\�7z~�p�ʀ��w��sj������k0�x�P�7"��l�+�>��208��R�H�!-�ݥ�j��y~?��lXe���;zW���{*��	H��\ɧR�z�4D8ǡW�7�'�2aJ��O���}Ƶ�zo���|(�|l���j>�ڇB�b�UC����Nn�Zrtk�:����ps�%u�-Qי�t7
F����]����9�~B�0��� �]��v��4g���(W��W:����H���<�y��%�˟�8���ve��K����B��!>V��.�%��#̉ͥ���_;���I�G�ӝ�K�%�z���3��nf����������mok�?��+%�t���hw�駞��R��� |�CSQ~���e�7T��t��(g��Kn��[Cm�~`���z���UT�3���W}������VO͓e�>O�i.�)���P���;���c��V�����S����_�vú4{�1c7��~	��E�3XW��(���uU�44zw]�Hg���*����7q�R�������+W&ԠOhb��s+k�ʯ��p�:&�O���?�+�����wD��q�6R�,Ac-���ӓ�|b���D�s^Rva�8۸n�v��{�Z�%X�y!Vĭ�(���I�^ӁI(��	3�G��2t�'<ӯ��`�i�����0c�tA�)��ŉӅ�^�ڋ1�1d[_�+~��[Zd:^��l��Md-�,��p������o� <����ް�C��C�/Z�P̓��MD���|]E�"���s���!È�#����T{�T�v� ��V�}N�rO�f�EU$z�p{9pV��	Ή1NTĥ��=�k��e2m�]��ÛE�^0���S�h( �[BA�m���EG�`�pӟ���^��d�{��*�~����A��3�D�+mF%u������	�N���?m(�:�N�:��Zʵ���,V��wҒ��ӞAdM���拟�b����߾�l2ȥ�� !��hń�����
�n����)�}lI��+��nlV�y�3���_����9��k��I|F���It�
`�xU������0'�� (�y�w�T�$���3��Ɍ��v�h�tƯ��P��I�]��F��+��4���^�ٗ�c���4R ������:rS���P�K+(��hLV�T��*LꎃF`��������Y��]��H���N��F���Y?��%��Zh��7SC+f)|���C�N��� �����eG��pb��!�o2ۘ��\-H"Ft���l��xEX�Ӓ��_~x��6��R�f�e��z��꫹����=ԔFjg-�͟��#�|	�o�[��[��z����(o��_��^;�>��;*�ʌ-R�_����J��B�]ji���w���v"[pO��1��oa	4��oR��E'7�N1����\���[��e�Q��t���W���#rI\�&�!u
?]I)�^�o��c��=+�_�YZڼ1�OmZeb|-���U�\[��_�Гhi������jp�V��מ�����cY�"V
��|]�"1���;1.:�Qֺ�(jK�?�[�KC��\�	T���}�1��)L�WT��Zgn/Bk� #�]1����9����K�$�b\"Ny� ����5���P��%j�Z���ʍ΅����q`2^Kj�+�ZLQX��8	uF�odmQQ�Ѕk�f~J<T��ţp��B1�l�����}8�"P3?$�k�1�9;UC�y����{ mq���[�,�zIy���(\�jQM���d��4��=B�.����b����
pa("��Lc˵ht�a�����: q`w:	!���1p����U]��j�I�0c|���9*@�Ō�(2=0`WՑ��hc������Q��<MS*�L�a�3�%so_�$���%l���FK2�lqm5�t�FE��|�ޥu͘k�{u�bJDzI�7�rq���a�eP��}�i;>���%�H�6d0T�?Yá�;�]nw��Q|����l�׾%��[�Ze�͹��Q��aK(��|�V����($�%�4�oA��A���4n�|�]:S�\�z�Zۅ���z�+I0 <��_�lܳ�Nʀ�>�&O�D �^n��������?�i�-Ⱥ�]�ˋ�m	�BHw�8�n����N	�E��	�"��/��N�o_ӘbنNV5az�>`��"��SE���	��V{"d�I�<����^ǡnr@ȳQ�8�j������굘b���IWF�|�Z��{`��=/�[��Ԇ.9�T$[B�zB��@i,c1�����0�쏼�c+q�V�b����]"�p�+V��rbs��+G؃�	5ؘ���:U��Yh�2�E�A'S�A%Y#���6SE����7�_D1"{5��:��[ԓ�񡾞.տֶ?25��Z2�/��N��$����D���8mOH�4|��_����Y��e���p�)�&
+�
s3�w7/CݞޏЖ�i�Ž�"��{�*��qU�96�����'�čTd)c� ~h�D��P��R-}��0��[2�}>�,�2y�g~ ��5H����*K��7�� �O�� �xHL�+Z!n���cMP#B���u�c�#O���_�jQ�p�
z��@�4y$
If`�(RG��B.8f�F�r�C8��%O���in8��>;���3~�ٷ��*#)"�BP�'s��2����`_���X�zAE��b���_��tH�Ɯ�����"�p\�y�v-����a*U?]�oc�ϙ#ꋇ�|߲$N�Jz;�+>�@.ʮ��`�4��#�r$Ic>ފ��ŗ�~��%*Q�Z2M�y!��q)=��������p�U�����Vҗqף��\A�O����!R��Ui����`�N�O1������>֏��g�W��~������	Q�ՠmI��Xsu2M(,gw��g�+[ 6�-`��=h��*Ewv���L].�Gɀ|���8�5\X�2� y������v`��Jv�S�k��y�@�.�}��WZX:��@�Jt��ʂ���f���5��.���^R��+`�&���KId��a�w��2�Z��;}uF�@�X���hPh�IQ�#���u��Pv=S8H��8�$�(�����v�bG�ٝ0w�7����,kr����H~���a�pT&���aװ<��0K�9k�R��I</�婆?[�Q���u	Pȁ�yi��E�XQ���<b?��Rؙgݚ��̱vw{�Jn��$\��($�W����S�v��8_�@���������%Ѥf�mIk�5�k?���	$�?w������`0�>H����l7�EO�~G�.SseK�|�J|0��>/�RZ)�@��{.��l��Hޣ\�����:τatE�8p���Ǐ�0�*y�����NC��š�d���`ԙ*������PV�<ʁj:�wQ�1�+��D.�Ѡy������P�	<�#O1ꌉ�J�ы�ˉu�)��8NgNǋ@z��2g��.�<�v����k=��EĄ����e�2Ȑ���\;�Zq��ytFw���y���tp�'�\�[|�����k#E�.��I���W}���}���� ��8��}ð�ơ����r���xXZИ�b�*5��'�.6mqh*&Z��?�����ĳd)���L8�-��d��_��#�K[�������
K�j
�䋏.��݌�fĢ��%��6!�k�	x������L�[磽��b�,k>�x%,{�M�rwd_���G��'����+y�d�fz�RV3�ͯ=T��K�n�7�Aqw��L鿡O5!�7چ
�]���W�i����bF3��w$�B��Yp5+D�'�|�N������ޖM�'�O�b�Ԋ�.5�[t8z�"z�e�:�vW!�@���DP��v�
oW���ܕ��Mm����A\�n��W!��*�c%��S�z�;̍�K[B�v���͋�ıZ����}���~�u"(7�N՜�4\̐F���l�E�T�m8#�v��x<�]�@��R��v��+ӨklQ���2ly
�E%\'�e��:KYB��	@L�C'~�j��)����Z�>Ֆ�x|ip��e1H9F�5��a��;�=Wq�`���A8>`���%�VˣX�<�H��`�6$�L<�BA��ə7վ=�z��O��)��G,sbi3��Ϯ)�=ďM�K�\�l�e?Tp�v݉�q���+��N�+�û��M�밳�R��ֺ3<���L�����ª�3�7xQd�mx�6<��@pw��B�� ��J���"��]�A7_��k���,I�yg��|�|�)O��'�u�o��JL]��1UE�3S#��ܨ�,���("X�,��f4�q:��V�KR������nq1�k.����D4�j0�o"O%t�o�6@�Pmdj�N8)}��oQ4�ӳ*y��f�̟�j\nn�Q�\R���9[*P���T�B�S$�2?J7�@�%��ģ5i�OKo��,�S�lr��.�-C�N�w/�+�e=���!�UL�"�AX�M���J�0@,�d�M��\������UQcW��n&S폍�e"�;��A�N�Z1sn�םz�nH�1;^�����m���P�q��ת�}��T1�
]�W��MIԼ+�s��,������W�����6]A�Ѻ��oF;7XOF�G�v��Z���ƋW6x�.���!�ߨ@����?^u;ū�C��,�)���T��qf�z����E��t:�#���.qY*�hj��?lY��,(a,�����^~��]m1v��j��rP���1� �'<.%�SU�ؔ�!��l?�&�L�t��o�Hݟ��qlG�Ĉ��5�3��ːi���	-|�͐�Np�S�<w��{(�eS''~�$os�`�]Nk�W�&�Tΰ��9/"�{C�n���[�XM�Ò��cQ��z������g�?g��דjHN�5�,YHu4���k3{@�|�(6��֬�s��A��7b���2K:�>ޓ�%�%�d�U�E�7�s��Af�L���zA�g�n3aX�?-Ļû��}utm�\� �� Z'�Y�jJ�; 6un%�.5�(�Ԅ�
����6X��y]��"H��źW�#z~�����j��ℙ�)Xou�{��'vEϢ�-���&�?[ʙLG��(�4b�Z"��B:,��Y�~���&h�*�=�wj��Qd=���~*���^��)�Twp������}L�ж�@���/�G��6#'�tI�7@�!�W�lrG@�@�+���O�$��2���H#
#�b��K��ً��uYZP�6�*�n����WR[��~�BR	�ƪ)���B��{���D<nq�u*�z-�z���۰�"��Utd���+RRzdxfja���������O�fg��lB��r���[.Zh1T��ͮ޼�:��&�-��?�M%��v$V�E
��A�h�-
�r���U$�J��2��ɹE��E�K��6��^*�#M�~ I�s�c�-�����2�#�ѯ�s��6�蟭�����<:}a�u�"�.��y�+�Iok;4ڽe��W~W�}:�sG�����
kI-�
f�C��YCw�no��ڧ�����.n�,�+x˜���%�Vְ�Z�n����!������%���6��TB8������5���{�(�eD�&�Z���a�_�����ھ}p�2FE�*�$$e�����[�{��R�[7E6Ig^%��Z�%��3�&Hy�u����^g˝��î�i�.I��ԗ���"��=]O\��5To���g'�q�^��&G��5.~�o��F�����Q>e��FP���O�E��Zu���F���j�ո.�åW���c��)xlX��$�ٵ\㿘>D}��ٜ)u�Z���,oZ3�<�����/�xRB��/hS�=��#�X��g"���٣�l�%:�KP��K�f��P��Ք=�n�#��.�Q����=�C����4V���~2����'P�:az�2pZ�"���r=B���a�5|M׻��b&`���QSkn�W<^�~��z�I�	$�2ϸ'_�?c]A`G�~8��e��-�p��hH����h�+�I%�!3���s5���pV��{�Ӑ�yF��lL��8�&��Lf�cyj.��e�|�iOTv|�Kq1�4�q�Wr|0F���nlﺞ,��Ϟ��M��7�����b�����H��B�xm$#��&��X���ryp��ѥ���^�uP<�>z��8~�N��U<��ǋaψ�kR�ºz��5'��;�Vf�qq��k5{�չ5o���Y@�u�"�(N3�s��C����?�t>y� �;(v�)qU�_м����۳tk�%9}C#�;̻��e�t���L�n��X}]��s�lX}]��xh>�ׂr}?\hSЫNm~�s�uuq�܏�`�tc�V�3̝�e��Xr�ĩ���B ��%��r	S[5�aXM$A�<nFB�1�{o�o@}�".����ƥ�A,qV=IDs�
P�P�~+�E+��Ch8j�/��9�r��CЂ)b�(�(�%���Y6%�CǄGC
`�2��W�&�A'c۩9�,
0�a����]/{���r+]E��2:|ǥD���xz$Yn
��@����w��bG�����ɖ��
��Ĉǂ���,���C%n���pwG�N>�l
>'�i��=/$~<�����۩W*]�1��I#:0�%�:��̾��,)נ�K�}�Zj��y& ��r*d>Sm�T-h0�r$n�<2do�3��<gu`,�S����L��3�R�m3�����W'	~#��0;���n���bK������]�V�uB;���zqN���n��a˟'m8�U|��b�=#��Q�a�`�A�+��>����J��`�B\�����k�/Q�'tzݾ��:p�d���Ϫ����^�sܤX��C	+;ǿc�<|�wp���I�q.9_fF��"^yk�YhV�.�d�
�\�w`�oM\�47���LUD_^Y�肱���ԯ{�s�+��3�~�� l'�	��y"�v�u7� _J�%7�T��Q���p2(�q��d�Pz��v�菦bQ�9���O�ݤ�|�`ƕ0���*�y-�%�t}��A��e�n��M]=mS�>��)в�4�p��/Z�����t����Ϡ����`���9��F�l��R K��7<�������¦���7��h����#��+��	�N0��_�wEն�c�b�/�$q�Q�d��hT��F2�+L���~S�
Z �@�妷j��q��dj��@�_�[V�C�,��8��P{�����+Eq�4�)�Ki�9�[��>�k��FI��ӡ�ZwT�ױP����5��v! �6����� �ex8�y�rk ��k3�A�j�~�÷3��.�ұ���������z
����X���OB��W</]�Ӈ��TG�3f�S���r�Md7��)W&���3\��0�9���8R3�\Ӏ��;Fԩ�Ď@��LAmb��R�'�'-�yճ'6ֶ@��\�DdV^CO�D��n"W����s�1�W1W���ĥ��=B㵖�`�R��t����U*W� �念����A�(X�D�`�vRVlr"*���
�3X񮡥O�v�p�g�o���9���ha�
{u\(�o=V�F�A�Nh�I3\Q����<��d�թ����dǒY����S��	�L�@j7[�����7�>��C�cSN'��9�n��i�Y@�M_^�I�Y���IBm7�:����{�i�J��ׁ�q�˸�YL����7	����[b���p�ew�������e�����ͽ;�5�4)�5 ��۪����vFD�Pm[Upy�������~���
��\x&\����6д7��_�����{�H~/�03��4r�S��1��y��͸���*̈́Q�_��7�K�%-e3x:/ʂ�*`iʾ���xƞ�g<	7[��m~<���0���r��.�>������C����N������zWd�C/<��5�X4�����b�4Se1}|�`ɗ�û�CP��"�u�׽��Y������@O��>�1ly���f ��v��O}.3���Q��kf��y��pd�!$�V8����L%�샃&���}ֶ���١i��N:~uSt���#,�Ƴk�����*j<��m�Z���Q�-7��J�Z2�5�눱N�������~>}��v��d��l�q�-f���,�L��P�`��\��T\���E�\Gp
z��W���v��x�suX��m��Ȣ~*�E��޴����KS#1*3�陼��K�W\��֝k�[���o���20��';9դ��ƌ�6�Y����v����R���F�nV�I�M����%X[)��-}f�>�U��%C��V��0&�P* �� �(kݏ��{S��fZۃ�d���D"HR�
��QDG�ȢJ�X�HK�G��#�J�pƹ2�F|��;l�~ry��o��V(�$#!Ը��@2^��fI�ͷ�k�>��b�늲X�͋����f����t�J���j��K��Oq��Z�����DGu�-b����3�C^�|\�)ld��Tq��{��&�\�b�W
�M��@f"Z�E �s�1��j}Rͯ
�F��A�mx�Ϫ/�pK5s�0�z(~�<�Oy�1�Z`�#�T����Rh�J��L&���D�� Sg��_�V��V\�9{N�ϻ���zMƌƎ�����%H~~t~������a�\��Y�
9-��/�|�&>h O]@����W���O@�a��-=�nu^��{J�Zv��6�BzvC�5�~4&ع �v$Ed���LJ>�aͷr47�$���g��Aar�@��ܦH�8����y�&�6�߿�!��"��FqGA��뭏�]C@�o��zg��PGy�h# ��/���%\ge���$&<����6%O_����ܪD��1�u5����;j�8�� O��a��Y.��z�M�G�y~e�-��ӕ'G� xڐ�E��;aJ�}�q.>�\�_�$�7�� ]g��+�VI
Ӵ7�Mw~���A�����,�*���� �g�INwr�zq�#h�kq�v��4���������/��ujB����9�h��Tr�L�\��x���j���M�.T`"[���D���0�~���.ayI{�V��r�^��IIʸ5��&�6�dLۻ��`�~� اNh|=�{]�b�'O�d� �@ȭ�����n�|4��S��i����MC������Jʪ�X�	v�!� t�<(t���bd/�e.k�B����b+��"�I����Z�	\����L .�<.�������^��(W���᪁h�ݦ)���Ĵm�f�(�@��u�y���хZ���
���V�yoi?f�I���w������Z���0��f+[T�Q�ba��h�.�~G(L�lc��Kg�yx ��"�s�K��8Z7�=�1l.?SN?����8 �U�Uf��{͇;�p�]�z��	2#����e=�`��M��,ZJH� v��`��ӽ�3��Cp���M
���Y���}��
c���ML]��N}�
���#�`���¾ɿ�˷�Y�9�4�=��X��t��)n^~	���Z]3,�CCt����Jd� ������](G��ڪ��������긘���yu�l�㡬��|��I�~��:�)6����(MAR���&��\��
�S�>p�_�����$��6����N��T� ��+&�v��:9�@��9d�F ��j05"L�p��)�e��*e�s���fnvKp�<�*@C���9�����8� �xP�	=�
����^yֹ��FzXQ�E���"�C�w]o �z	`K0���f05�. �ݵ��:I%B>���-��m�FhB��n�HE�Q�˘�}U`D�O�����B%�z߶M)n��L*���c���^��e;y @j�$�yq_�N�<�*l�oh3*�dg��E%Gx�h�R�u�Td����gl� z���m����
OA�S�L{h�tFt��f��ynH�	�����_�A{u<���@��ks��7�֏�MDQ[*6����l9��]	RB�,�H�̑}��}Yw��C���b�����3���9�� $���&{56ko��s��x�c��	� o<���'�O���c#Nh��JԐ�t�ǈ�mf���Xβ�|^�c\`�J�҉R3/�N�[����c%��!��2�UЬ����X�ة�Q�j�3Ho`nI�ߠ��S�$�j)o�%%��:��3	����B�W5��E���,��c�r�"���i|�#}��3��yK����hX9f1�ql�x�l:��Q��^t׏	0��S{���iF� �=C�"��Ԫa& u�j�$V��m����O�Տj�'e�����ځ�7��tϞ�<n'̷$�;�_F���N��J��Au��֭xɎ]ܠ�1��bv�>�d�����~ij�Ck���H���Y��;v��?��I��}{��-��6���7��m�W��>piѳ�N�o�I����K�!5ә2Ǒr;am� G�ǒ�S��EQ7�7*�?i"6�ʁ?�4+.�����V�)��y������6�jԾ�FL���G�����9B<Sл���}҇ >�� ���3��OKش�F�55�}N�<pg�"J�S�v���%-;P=����Y���7�W��j�,CB1�P�zǱ�����o�b��@'�`�H��F�I�>}~����R���H*W�`���C,�k)(hM◻#B�cցo��"�v��щ)`¢_wmvg�LW}�ley�kV���6�؁~j�����Y�2G\����:ݸk ��%���J�v姕j� �)�-� ��se�?0yA�G��Zr@�:���bunόPx����_Fu_7�" ��,�"�Xt �{^E=�]��p����k(N��p�k�_�Գ����A!n珺!�)[�=�a����!��O�e�t<�H��3\MRD"K�R ByO�Z��0��@���O�|s��g��F�������e��.� �K�#dvg�_�+~q=*�ߕ����Ȥv-^Y|�X ��LR`�`Dq�����t�/h�vGU�P�%X�R�ܲ.f��x��^~j,Y���ʠ4�@Zz�D'�c�$2n�qa����O��S�i��t�]d9�.7r=�-�,��0Z	Mj��������4����k0�����~��p�~
��J���ԁ8��:V$�H���-��*h.�\{]�����	��f5 ��P��g��Q���s�(/�ظ]�7+1Ѓ4�C��S�.NTfCy�v�����������Eo����t,(R�$8/꿢F�l.�տK0B e��(f� Ͷ��N�3KG0����j�z�N��nf���Z��ަ�F����{m�Q�&��{}�-C�*�xC�*k�ͺ���=M���Q XDV�h��m���7дu@��u�2��?�FN�R%�=���aD��i�jIB�X6��2�����#��a�Y����O�d���+,RA��8A_��g���+����Y�Kd�`��kS#]�<�j*�G������A�N�w�����P�x���"��~��[�.�(�D�L���t_Nz��5�a�?n��y|*-^�n�#QHR����^A)=�K[�&�:�z DF��.�й�r�c��^_%��1ֻE��������CǕ����-c��x�C��-�^��"�;1��r���VD���6�1����܏�ΰ���>�����e�a�ǿ�G�n���Bs��7���rI�C�d�F}�'�%�Ը@>���f�ob#�A)Y�w(	T���zo8`��{�p�*ǵ	�A���E��~��n3	U���i�ۘ����fF���0����t��2�N
�Ȅ�'�~�I�w#��ܤ�4A�[@>5�M���ҾI1��s���
#2�Zڞ��m��@5@`+��_յjvw_x(F�$ڽxP�vd1XZ��i�kP
�e�@��|;75J�z�i���>K�<gK��dFY�r�O��a�Y�W?'Mzbѧ&���B�S!<p�)u�`������-�¹�Q/��T�ɉ�:��Bm6���ù���l�R���f����v-`�d���pt�f�}�9���UV_���6WB�5sB�
�B°��:϶��@���q!IH��񜋡��~�GJ�����9v�&W���He~���Q��h��H/VmCu)S7�-�YJ�C�:D0rGsMJ�����]l&�=�/8�P�R���,D���s��ȁC�t� e��AV0K��	F>�'�5�h�ý��?N}���ܬj�L.(��J�v1ޟ����u�m�&�\oyk;��L����L�	���@@$ڭu1to���9J���y���Z(NJ����u��|�C�VZ�u�Оpc������'pA�"���^�c�l�D	Q���T��:	�0-Bo�G"��#cB��`���Jܧ=}�:U��ܸ���R5:;g��M�d�;(�� �[�(m�Q�a��^F:@`����1�2-�L72+;�Ӟ��؜���<gas?�c �	
�\M�&o9}a��_�9�l�1S�D�����6�Tr$�����z�� if�V���2��y�",!���x�p
���Cְ7M�r�Z������jN�qlV��� �<٣._�h�ٰ|��VV,FD�%;��[��I�~�@C[E�MV�{��3/��B��c;����2�*{15���b���ǎJu�.D�C���#kM�'����hv��=rQ��$rq�S�Y~m�6��1�<��י��y��AA���c"$∐�6��ğQh��bD>��l�J���f�YЙ�㴩��k���ѩ>��+������Eomt�(��-?��aD~PxC��|�Sp�!��Pb%3���h:؟���-�\_H�����#<�Wc��D�q���2�b����F��8��2V ����\ bR��S�Z�	{l+\�W� $�3�Rvvl_�=�Ř��O��Sq:%u�fN���������^dj�ő���>WHV�Yěn�!�2����!�3HU��m-�i��g�ܠ1�~݄�Z[�6/�[16��@o����^�s��p!�C���ڹB0��]����X�cQt����^���/3hIC�PP7t0�a���ջ�xQta���%'�\OF=�Bh�ѰG\��5�h�m�+~�Y�q}�Q�Xgl�7v7I�]��<��aV�B͔��V���
(=R�WZ����3*v����=����N�>t����1j�����k**P�b�0��
DXj�`�;W���Թn��c�ik[���/_MV}��,p���ޛЄ�XB�\�4����h � m��N�>���x�h���������"�i�C@҄-�^%Ԍi�$I�㏵������X�����.��zI�������ݒU�Uz�]Tt���-ٍ��\i����j��Lx3�p�L?��`=-������s����)����]ӭM�M�&�fo;�]��1}P���at'�
K�������]E6Z7�~�f�^mF�Pз&r�БZ�FV�p��b����N{e��fv�U����u�5Y�I���k-;([�8!�p_X�n	����4)ۘv�����T1�⥇1ϽG�P�P�����
�}�S�ǝ�Q�T"a֧��m���krf��F~Zh����{F�J�F����K�G�2�x�'-xȗ�2Q�
U.�s����+9n{}N�0a[��cL��:�g�n� ��l<�Z�P��]��$���T*���G�n<wUl����J(�:���c�Ԍ��\��`q��`�#=��°��TCXT�c������)��[m4�:�'�947�����Y�t�R�u�f�S��ڗ����&�����=�ZQrzD�uKɅ��9̠����\S(i�]L29N�8��J�k�/�殃ڒv5\.�R�eݪC�x<נ%�_=
-��=Y��%��ⷣ�а���r$0y3�AlľjyC2j�Z[�Q;E�,��>4�	�M�%#��	أ�r��������S�������g����(}�9��[
7!-�n~�>Y`��3V�@�1.�FEL�n&�~ހ�-l�ã�V:6p�n���n����3�mc�)��܁f>�k��$�BT�� ���z�T��ڻ���Ş����9s�p�H�m�1UD�h�*IMJx��P[��¿���Č+��{Z�W��{YM���֭:� �?��˳*B���I�.Ѻ��m(�6�ժ����Fڳ�B�M��1����"�*�0Ff��[��~c�R�85�S�1Cg]
��EHMה0�Dt�R�l�5V�m�AS�AlNd�JT&(1W|��H=�º��i��kLd�q�m��D����$�0hu�<����V/�UC.M	�v N��#�t�'��hR(�S]z��u6S��S�ڳo)��FE!�(bM�_Ү
�1�,ٰ��??n�^仃y�w��F�q�a;'�C�T��Qx�����G�5)(�O`_�vᮕ\����|�NP;�D��7�j��!���ϣ��{�Jݲs[�|(�*d.$q1�c��{�ޠź���x���.�����&$k��G�]���^��q9#�	���ə��5��>��WV�ƈ���xM�(S��.H;4C�?5�
B.�cC��|���Fr�y
�f�8����9�v(������=?����p�M��.��AP��N��!8O�� r�F_�󑫲Gg{�#�`����WX҈'3�6�biK�v�-i�3k�yZ��S/�ԧ�Y
�?�Y���8�Kd:�繻_՜��q�5�s��@7��u;A	���4��=��֥���,6O��r2��)�J������1�sP-�^P�V�fO7U��<����å��p��w��gWI<��Kd8����l���*"�s��2�'��4Y.W��`���W�|����E>��*�\�D����2�)�tR�H�,5\ʣ85����fY�vz#���^��3V�=�er��:Jڂe&���Ea��;go��x�) jl�hb} �����ţ�b�g��� [�i�����,�{��P����b[]�)�6y|�G P�i�a�D*!�|��ӧkK�l5uic��d:����Z���(�Pʦ�5_>�`�!��^z������#��	��ϵ��{�	@E��t��q����&�u.�rGgXG�~�&�:ÅmM*E�*P�[x*��ګ2��������)�X�}�s��;��_2v�@�A�5K�eQd������i\f����\�<-�V *T㲢��-�̹��l�$՟�b��l�Ʀ������OR
IpFa�:I(6Ӛ�������xX&y��A�V�!�%�Q��_�]�r2�4�N[�(�+u�7�HUs9��ބ1��u#I�����'�p/}<�8x���bUR��`+���3�E�Ƚ��t���8܎�����"7r�o��:e���8�8^�VP8uV���Úk�<V���,�X8s׳	&FS6"�5��gT%`,>���)�qIIh�|���l��OVs�ܑ�z5E����]��i��Bp���b9C3lϥl��^t�Ao��QU��$�E�}H���{�\^l9���  ֗ߍw����=Q����A<h�\���p��3�A�γ[h�����W:�4�/~r�Kr���Ǭ�C͍�!dH�@�R�$�]T-�73
:U�x�Щi�"�k������Zk�6$��O�J��+5?��y��:�|el��S$�'#�S4�����.����EX׋�+6>��)BU�W�.�s?3Z>��g�Wb'������)�O��e'�~$gb:Y��Q�}�6ؿce&���]����q�w��}��&p2^��!X������ �,_��&�"��������r��,DL��Sn���+!�}-��DQMoYv}�d���`	���͂��(�P���M���Tf>�8���v3͍f1�ie�t7T���9��t줦c�)�]�#!/��fy
���!&��X" ���	����3�e�p$ŭ#}V�W&������v��v�����~kݚh���&4R��)4�N��Ԫ�8�'T��Օk�����a���?����DP�ݧ>�]���(�� �u�ᘑY`ЅIe���f+���u��;%����P�s��}�Q�������CMï�6bM�zo�J��N-� ڮ�{�b�� ApY�0�$џ�{��2`c��#��{���]j�ITj��	%��3W�����l�\���,��%�5�+a۶���
��Xg�S� �p�Ƚ�ܲ��#����b9�j�[����˨_��-���u�=l�4̟2�O9��rN����m/	���˻�-����?�~�ގ���lMᬐ��nF�&�9��3sQ���Ef�W����Ȯ�}f��S�kH1�Y*&>�	��m��Nd���/ޣ���8�x^*�:x�a�*�ħ�V&�?o�I�F��-�G��뼈V!�\j�&lƭ��8SsA^�qy'�����v$H?c�G��z��3���=�����kE���s��Y��,H^?������!NC�A����a����/�u�qH6�����T�(���~w
ӑ2:矑�V�k��>6�a
7�/�bR[�����"樑̖��0�D���� ��."�1t���b�g6.�jң��������b�������M:����Z���J��LL�_�rg�3BTm�������]��qb�6-�c�#��:���R�e��?�Xɸ�|��������UK�hV4�\�8�SVe��a�k20�w+���x�L��"�w'���Z$��DG3�w��pL$/����H���+,��[�M�Z�����6p�5:�E,+�=�C�4Ǯ��W ˟������-�al(��u+�F~�����W\�+'C��,�����qF���n��E^<�W��~tNC-����Kӣü�?�D<_�^�>�4.qSj��D���h�mgm 	��{G�"�B01����g�qc�/�G��H����z��[��b<ʭ�/�*F�^p/�e ����^^�XE� ��K��7�������}�s;.4
ݖ�TѬ�arr�#,�H�n����z���Ȋj��.�j��sr~��b4O�e;pBi�.�]���"^��`�#Y.*[��b:��<��C_`�!��nJ&�9y_c���#�!��J=d����qi(�\I�j���1���V�����T>�����j�����\/�SE�����9�ӗ⋚P_�>'b���My��%��'y���ƹ����2޽�ze��!5Ci@K�Ux���Q���}|�O(̤=�5`��!�nk��I�IA�q�Q"���'��}��|R��D�t��N��� �k�!�r�B����WjK2�9A�Ϸ���N�'bC��=��~Rȵ���Sf�7�x���C_WE�yu$���_G�C�H�mIZ�a��O�c�D�H�� yI�!�oyu�8��C�����77H��"���ō�GgW�5yJNs~\�'M��ƺO�W0XC\����d#�9�Y�� /�V��ذmVj�L8��HS�Њ�P7#<�Xw�ǨXev:}��▧m&M�EXN����>��eI}�ӣdE����֕��Z��"�i}S�O�p���u���ۇ�i�Y	�3}�T�no��	qu4��2�~w����I?s��k�ŋ�K2lԫSF�� T�����|��tS"�K��6y�"���!ճf��H4[W������Z�8�cE�B��e��O�F��U&���h�K]�,:��Y=Y�}7������Y����%�f�2!�8	�q�XV��7ȆbIS|�׹�<.�20�V���j�3KtEV
��+g�_Y)��zX�SK�G�U��q� ��1ډ�$�}y�'Y�79��`�\���F����.�a���F _0��a�h�C5u�P^�ڍ���u%eC�Hxp�En�3flp�`i�7[X�:"��7�C'x�jm����d=��2�ާu����u_������,A����Y12b��$9�/,��(���o�t�JǸ�6KާXb�R>椘�祰���D�@3Mo^k����.�Ԗ���Q��U{��޴�Lנ~�NV�p ��u��ƿ�3���|!:��[�
��mmR8ѩ��D���]<W�?]恢�d�gV�?u���G������Ԏ�_��bhU
�����r$j���M�4	Iz�%�i>�2T�ď홅e�S� r�Rf]�Mh�j�a!6�\�(��/8<uf�,!����)��G�09xͬ�s^C^'�q[�h+#�:1M�<V�

�e.�B�7�_�	c�S�T 7㑠<x�R?��y�;C�&/�f-	z��z��>̑7�J�bXA>�NS븘qG��?w�sr�������)��u�CEE���u���L�f��m.��a�S�v�s���2+w��Q�C��yӸa�-'�]ͯ�e�tq֙��b��O���3,�"��{�k����-V��������7cM��S�ltd����oh0�c�����#�^����]I�R0yʬBQ���Ƃ����p���!���>�c��cU/���k(\e��:��l;l`M���r��ƥ
��L)��Q����&�f�Pu��#SoQc����|~M��(�Q_��G��~j�f������A�tt��>�r���97M�I_��:H�H���gZ����} ����+�Z�[��Q��`^bgKpj�,Y�m~~��s�q����"� o%(���������m+ SW⬛��hVORg�]i�	��%iO�\�J[m�?�;���Tp�0}��ve�ɉ�8����gu򄝋� ����j��n�V���v�Ѩ `����X�~[Q��EE�"$F�{�4�s�wrn�
^��2�г���X��gI�@<�'{�
u���0.`��q�КI ć=�I���F�B[�z�z~��32ٶ���gt�&��1��@�ɄRYm���1�W���F͖��~e�S���nw�4l��mNn��~ܺ�f07��7����<��ń.Y�j�&��#?*8�+HۗG�9U�Nb�T��A*�#kE�?)�(�Υ�@͚x��G/Jn��0r�o���Pd�k{�[`Ԍ4�����:��CDYt��2�gG�X%&VU�Н/���'}����Y��)��lG�qU�30V��*�Ĵ� �BC��DjK?�U�?b��h.6�2�;܍�nF��}^�)���(����/�I؊׫�>��F�F��H���0�*�`�����(�W�L��(�r�ퟭ�e3 �����4�a��H���8ѨR�������*`���K�$�(��nw�JԢ��P����5Y�D�QeX`��e��4�R���IiRP�MG�{8QQ�6�uU��)w��ܶ&��>���9F@���Fm	G�p*n�PPg�����8��@�D���I��``��]E��/4�r����<�>�����`�|21���̳�u�0�~���6�ʴ���5�#�<��c*k�lt䃧�5�J�S`�
�A��x�.0f ��x�ܟ�N;Ǒ����S�~^�|M�rr�{��1��YY2?��I�[{I���ä�0B\����M5���&1��і|o�8P� �^����$o����u��W�<�ߣ�Lܥ@&bܾq!$g��s��h�n-��3���!$��_��n[f�aY��4�j{��HZ�O�����D7x�&	Z�b���1>z�I\�S֤%�2+�^��&`k�t�Z�5����ܣ������-B���!��i��Z�1f{����G+�(��n��c�̤NfϞS:����Y��
��;��	4X�$p=�ؿ'��m�눩�����ܢUa���c9\�8	+
���:��e\�Y]&u�k��'�:����u�[0�g�Zw��1���ҫ�f�6���\h�{���M�3�T.�2Y�8w�C\��}�b�a�l?W\�Sy���z�^��^,�t�f_Ph���Ouɇ�d�� o������"t�`�� ���T��o9@ٓ(4�YE2"���y�ncǫgM�\^�=�-�.���wW��r��Xʻ ҟF9�l��$�A�=�W��X��0ɶc�I�]�ф����q{e�D@�XS@��Z���J��V�.-��;��D,U>����/\���4|w � �.]�ɥ7��:��	xͭh	|6�bfR�}���W*�N@�FƯ�/����|�EH2���{4t[���+Kp����G5"����7�*T8p�Qj�}���0����տ������G5�����aޚ��U��&���?�r=�S�H��J���H��\r���Ʈ=�Im<#5GZ���jC�ɌjMb,��
??ex�:ߖ;5��Ŀ�ߚ�G�+{n����G�����i	�b�/'tw==q���oNH1�F{��&7�G���V��������J$�\Z;NJ�(!m�/���%��K��;�W%�IPI���bQ�Q6��k�Pۧ/?��߄�4��l�!���>_cC�%�j�G�̈́�m�	P���M��ٟ���&���sN 򊰀��ё�3	�P��i�p2�hfo'1)����quk�c}Rw��*]���
�H����
��D?|��S���b����Lp��w����0iOj �
�!Ivˠ��գC�.��3̴��EN���;���ˏzYj�PN{��¡V\��C��$z[����hG7y��Ǯ��%nlb�����0���h��&qM��9����a�[�_�üX�M������}�s���sYB$=W�?L�r�� �u)1�6�6�����������u��P[��?�t�`|��I��������^~K(Q`�m`�zj;[��?77pOeTQ����g��ӗ��R����V:�\K�p��kq �i�����
+�I�P�6h�0mqh������Q�c�)@���v�;!T�\bK�{��A�u7K�;��~/3��{6�o��K�a��1�{��j*�hJ?J�{#���@f{RLNW8�|�+K���Y.�����^'��&��nd�$��[���x�m,�1�=�Ɇ���ߪ�'��Rw��nlP[B��d�ڸF�����o�]�}n���.���9�3/�8��_F���ڳ���O<�`�'�5Ng�m`_� ����G��t(2��c��X��K�Gg���f������dy,��'6?Xj���=�,�#�9���V�H)oV�����:ǤC��P��Wy���w��3�#�#V.C��Ό�&�ƥ��lIತ%U)
��Jȓ�1�\hg烷(Y��÷u.�8�K�h�"&�t&�`s�h*�[��r��/�u��xU�0�ٹ����@��3����1}��\B,C��pDcw�*�nM�V��A�S�O�&K�o\jV�Y�Eh$4���]�GJ���ʳ���%�z�n��lS��g3�B��Ҕ ��r&�F�;r=s��G�]Gr�֘k��7�,W�Јnܦ���f�Ǩ�뚝�x�3���`��YQr h2�r}�8�.�x�J�2WA)MR�E>=r�
�G��zO5�r��Ѷ�۔8p� ~����/]�0�7�b�x�Ip&��TTU����٬�_�")b`Ր��Etx���B.u�J$"�f7��ET�/L�*�a.��!�p�QH!�{;qv�F�'O~ ��~rM�:[�:5L�K0]@�-�ُdp^�P,騝T��.L��-�d��vc�?�.�/���ts2�?7H�r�E��k��Z�B��suU��k~C�dm���1?m!��;__�y ��8��5�b<�J��` `[�>���ڸ�e���D�8'���х�Z,?�K���Lſ���W�8�����f����:���J���Br�_��"ҒP�̹�:�,⣿��Ն0
C^
��2#q&,��3Թ0���WVk�n�-�I�y�\D��_O�����b����B�J,�Iy��D8�|���'WWc!3t��P�n�
��J͗F�C��7�/���B����@�~|�R��=�μ����6y���l�����Р|DܷS�M}DE�ӯ	�C��� ��ڢIRw�$�EzB�k:<�:b-N0�0�;��q�ѝ��ֱv�P�[�w�u���?�(�0�[���Z��!�5��G����5����!o�."�#·�Z�N�:fd
vQ�<+���%�`�n�.�|�V^;�����kő��h��;2�aYSO�8#�V���2U�Ku�	"_tz� qgo��n�]��G>�=�V�=*f�ʮ�� �6e�X�Z�uI*�8����2�m+|�vj����pӵn��A���`^4��Sd�����*��Ë!�?)3{k�%ܭ��;��:�7�[�Ӥ�/�,�Hvު֤���i� }o�+�v���:�,�����[E�_�aH:�
��c��%��7\e��)-s-��y�&I:����n%����l ��\�>"�	�����^�Q&R�8���cűZ�#�^�Wl��{�}2�Hq�2R-=ue[����Q����.��а9��sk�In��1u�d�����T�ʳ�p��Y��<:��`v���lX�J���gih�"A�,䁂��������H0�d羑�6�fi@o�0e��smc�\�Qf�����e#�� ���84�BX�ܬ:&'��,E�76з CXo��i޽ �$Btֿ!,���(��qWXb��k��T(�lzA�J���P���7wTz�t .���1��<o�VE��ę�K�����
68vI�P��W��	+U"%�Jcy���f6�>Ō�|���&�VmX�S��8\�l�M�Ԋ?�r|��D�W�9^z%����y�S<Ra�3��N�]�c]���*9N�u��S�Զ����0�A�֕lÑ:�p����}�u�������48���c5�H���L�lvW�*7+�Q�HT~ zb���ۨm���σn���וD�Q��rU�6V��M ��n}y�*�Ig.h�*�<¿������?�(���l���dY!���q�=��6<�$���ox	�;xP�l�yM{���|������ÆNܪ�O���D^,E��ó�@eUO4zO�RS��[o�U��'�p|�=��d�L�x����D�A���s�o���xJ9���v�77:�*�˝ ��i�aG��iaŭ�D%?/�C��9�	O
��0�[B8uH]ߜҔ�tOʲ�`�M���69/�l9*DE�Mb�Ǣ	
Z0�m`K����7y_�+�m���_�ب"t��CP�����mM�ķQ�5]vB뢧���)8���%�<(��0�3yL�����������C舻9�'¢Z�?ʺ�Vk�0M��>��?]<h0�4��=��ݚgҀ�v����� �FSb@���b(�� ��"�e�~yM���G��0ҽOa��G��K)m<g��b�kRf�(� �2瓴���']���j���I@���HJ_��͍�U'�@4gz*�`4&��>v��#q!��A��aKf��:��
�Q�Z ��/��C'�8}���:�BH�����D�Ca��>��R��|�`�=�9q��!ڻ
y->O�)}~��=�6�P�wi��_��ٳ��|H�_i��׏��q-� 0PU�W�H�/B�� C,���\�b֐C���}����g�,�Z.�n�E�9c0�sf!�6H^�V,�$����^�;�#'u|�b�{:���@f�vA���`�}}fR8T��߲;��O)����~ٱ, �!~�M}�_�J�TY�`_� �(���K;�NW,�E���jHE���r�b��C~$���ƃ���騽��z%˘?Q��~��*�)��m=�Q�Ⱦ+P��ّA�pI+�cU�BV���8����-��NGsP��ў�9��� �l�x=�I`��1TV�=Ѹ�)=;8b�s�E���
�'14�C�y)�l0�,#�i|
���J��}�O�C���= :��ܦ*1[��M���+f�b0�q�"��%i��CW��v�5:bpe��)AX �4霟'��_?7��bЄ�q��q�@V���>I2?�H3P�i�RI$�IO����v�KWADO�Bn��X��v(wt��&\�����j��a�� �%�	%�FD� �MU��جZXl]$ �i����Tnd]Į>qv���7x"���xR��wH�b��S������u��6�41�1�����4o.U�6$�׆����V-�_��,Ԫ�5L�׭�� f�IX���?tM"����ʘ�����l����Q���E�� d�$�����Ot�:��p�����K�aa8�' ��\�<Г<�$T�+�!���ST(irl'�G�IJ^��-�ȡ�pG�?ӱ��&_g��q�{%~b��E?�4�w-�$>7�
R��gΥ+[7�,tʏY�L�%w��a$��5�xn9<y�X -��O��<u����oɁ�S��\�Ń.dMm�e)~	8>���q#��B*M���h��~O$6�����iH������°� 	�ԓ�&�5F����j��3�$!��)����:��*��U%�x����ս���)H��� �րM�ȴ��=c䔌p�� ��wˠ|��F-R�#�������I��t��P~G���H�:gF�sߗ8�~c�xa��<(PàEH�dp�p7���o���_�LGh�c?����qŐ�pm�N�/Z8?��n�-j���d��Dlk�Ȇ�*�_�C���	�x\�C^�$��M��J`�Z՝�$�������
�r�IL?c�C*�bG?�Հ���V;\i�Nr��.12k�D^'�"���'l!d��^ZPf�R�ʿ�n��'l�αop�n�QI��-�uI%-�as��S��l_�JJ�_�2B�E�B&87^XA���ʰ��x�I
6I���l�"�'����Lm��R��SKy:vi, �]8XV�r�'��3s�Ԡ Wo�(M�������ĮS#�>	K.��"�x�������� 3f	;�A�lv��k�F�]kb�?w���xC͚$(U.�"-(ge���*K �Ildh&R�9��
�����f邑MTA��M,Y���s[�Ze��o��66Ȕ?%	�-�<�r�?4
��tlU��q �3�\��t)��k�)2���4"Z��YЪN��e�`�F�w��a�#-a̖�kJ��9�`B�|�;aBֺ�����2�mC�s��\O�x��v�yn��Y��a�A��pp%B�����ђ�7�,��˜)�������!s�:���s*�Τ]m����j����8
�!b3�'�l�Ʃ�7B�����̔�8"�p[�H^�Ϋ6�c����q�`�y�"�<"x�t��ka�N�k�a��N�E����0�x�R��kFs,s����3��
��tb��\6��y �`�(N���L�ì���Ǟ�l��G�!�Y�(����<� $����?d������ۭFI���Fq-�춤xE���6V�[=�Xc�T$�N7�g��|�Ώ��Y ���7�ٴ����E��gō�+(bDx�t�T��p�6+����4!��>���$�)�%NU�J����ŗ.�����H���4��9�z�e�h�u�F瑼��v�PȚZ� e^aYYr�۫��g^���	%�5�W�U�̻����&X�QBӽb�[��% �0�o��<�)��S���fɯ��ԑ;Owm7)��U��R��*�c����Aώ�g·��j@��R5����آĔ�P��}nu��G�a�*�*��\pzM�"_|$'�o�P�W`X���j3/mj�`*��d��Ƹ
?�q��j=�}$�81z�D�c}%{}����Z�.��簼�������°����a/��r�����.�&���4��.kp��E�BG�t�dd�,��?��{6& �u�O����.}��:lh}q�P�lѩ�ŋ���Zx����Jv�ڴ�#G?�ۼ:׆�h	,����U
�Ϙo�@~v|���:B��:��|����ڃ���]�%�BEAHܮF8A��=�w�S�ʻ�h���|E��=UA����� `���%IWgݴd^Mwj�JB�)4U;��'�C�S��^P�Hӥy��@S6�����=E{K��Evn ��w��v8ij %�='e<�o��n{�ف�S���P�D�`V��G�@4�3K4a���4 ����o�O5d��W�Bz���EcTյ�|$/=Ժ�}�!]�e��x<J��ޟ�4B_���x.N�X=��l�Ʌ�}�F<a��ŏ9�\w4I_]��w_��g�`��gtG�� ;��n��#�C�s�	��$<�`? l�~���^e��
��	]Nr�������@h����[^��̮ưt�C{��ЗVZ��J�{��he��"�$NmZ1�j<�ݬ7��^��J�z�Ռʗ�ϒd���N��N�S��=�`��䕥 ����lS3&�$��.�v�ik$�dG��0P��cLs�Y�EY��II��9�l����m���R�`o��.�z���Y�۫�V��Ab ��W]έ�ye���N����9=���Eł���Q�\�����C�l`n]�ù�2�}�{�oa�|r�� @����p�q0�Gv�hv*�7�0�� �ƭ�'����}�m�]�$�FĴ�)��.�K��p'�����A���٢mKy�c�8Eh|�H�=cb\���}���B#)�|��	��,~"���S1�����/�A1x�R>��;˧����t�{]����AU!>µ�r�U�������ˏA����	 nK���q�Or��/�#�GZJE����Z���l7�::�a�)C�����O�qZM��'��� ~����z�0��?6�fu��-�2]Q%4�狕m ��#(�Ϋ�_rJ?�U��Aҳ�&W�iG�=���	����J������3�����־�N}�mg����(�u�4V�H�5�A��Ab�)Q��3ж�Uzm���t�E�g	HQ��l�hjD��H�Ȼ�����b{-�jMf|~u'!.�2��=�����G���O��3��������w�%'٩T�P��p?$:�3N���Dʩ������J�g�;���`�_뛓��}����N�8r��؛��B}��cc�J�<%̴�W�d�IG��S�¸� k�� � ���<O��K*�]�a0*o�#��4lA�#�q�ϻ�]X�5خ`�h��Ȋ��
ӭ�Ab��.|dwl)��uO�3�s6�?�6(v��*����V�q��Pi�q*����fT���|)��"��KV�N�)��s��/�(�9	�:��T�唟y�F�$�
��.����n�K42>�{a���9�2h�;��O,���9�� ���1ތ�S��]6���w4�ÖR��W�hE�EI�AM�$�[�?8��D��bS�.��>kO�v/AOդE��{����/."��u
�n��OK�JA+ xV��q[�}U6�a��O$��r���r�"5��C}��qG�c�9:N��` ����v<c�m�Ȉ\}�4���RF#�F���ݽ\��'V�d@�D�/�����6�b��^x�zJӾ��7��։A)&�^�q�
>F�!��� �:O�pñ�v�����t^`�xЧ^dl�5Y�W5*_�'�����D���QR>p@�Hw��%-ve(q�Ʀ�w#1�!A��:�X@�4�}�'��um��3��-�t�2�2T�Fi���gyh-�~�|��g���D�a��	�u�$��Z��j��EPc&�n �/F���vW���	��T,gX�]7jE|�6�8�=�T�� �
�B=i�~Hldnj�� +A��q:������o�V�ed���!A�J~a��b�ܟ�H�8y���D�vt ��sg��}Uk(�pU������U�9�08����F�#�#p�������=uQ�TGO��N���E2,р�b�)��[VQWQ��]�y��ǡG��Bc������N��sh��̐�uׁ�P��v��|����3�^t'>�G��v�K���~/'O��mcx����镌�3�i���r]�=�}�G*%��.��J�)�)O�1h����yz<
M|�R:D��H�m�����(WҜ�#T�}��|��L�V���o������8��c@���E���O��i7VH�~�T���+�����H�O���%�Odi�>���0��CJRς�F�<V���p���Q^���Z`rJ�BI͒#T��6"H��7�˻��d���@������T��<':a�!Y��S�ȻFw'�
�i�t�4`��g ��4���-���vQW`�~�����?(���`~��8y�G��7�yl�[2�;�v��ʞ�8F�V�#R��!P���kK���9��M� ��"sS��H\s�#�E�}5#6�\�̓�fn�2�����5�;�ۃ�1�c���:"u�r�,��^S|�^BD�gl����A��8�a��?�1t�w#!�H������J��W1��!ؘd@�RSO �f
B�{�,���`1�@v���Lu������묟�*Z����QF24��%a���\����B6T�����,# .�&�3��+��N�`�8Z�<L�k&%m�_W���(u���r��s�������|[rn;���$g�4���L�������G:����-�U�e/��x��pg=\*,}�\j��w
f�Y�e��W�6g�4����A��Ѡ��nÅ�?���� �C3�ڥBC%�/1I�(��j5EX���r>G}����j�D@���N��y�X�Ni�s�F��0�K�
��lN�E������V958����j�˖�0���(���"���ˆ!�g{5�|^Ț�b!�;w&�6]tt����G��g�1\�����P�j<������=����$�&��ò�)켫f����C~j����d�y����vo���ׂ7
�_�@� �׿���e3��ě��W�I��[�y�OLc�X�������wP<$�p�	���\(��*>��ظ��������#��A|�'	\S1��bv<?��@,w�4�c9c��_"�AHS��M��W��
PnIV�)R�Z�����^�kPұ��<v;N��~q]b��a�Z2���4�����z'�v[]�N�Џŧ�U#�m�{�p�#OHt���aj&3�3mDJy�槀1���m6��~�׬"�����a����H����0vh7�y�֌�ک����W�f?�;��j��sE���#L y�^����y���;���,=��[V�/�/��$�0�����e�y=����߮}�B�o"�Q�t`��\)�� $G(���jI�
b/�����bGb�Y�)���A�ְ�ͧD"+�s#	6).:��א���? �D��۲��ؗ���<jRHU��̻��5�H��y#�Fu��Aa���#K0�P��������tG�*�IyM��v�b	W�RLOp�,)`tc"enͮ	 (��%E�;��e�AF��Mϴ!� �US�b5���`lQ�f�'�Onf�`H��SN����`4C�G�F�v�Β�BtPΤ�0{��q��i�L���""S����?w�g��Z�2�#
+�cUU�E�ٹ������~jES�x�W<��x�Ү���:�Q��y8�!�#�Fe�,�h�؎)���E]����T�7a��K9�����ylQ!���wJ����M�:l�k���k�ް4:�}��Q�����¼{"��?ɇwO *��+�݈D��u��E�̫җ�˕��MX"�bzf��θ{a[?EA�������Ԅ�GOM&~4 )%(=���m���M�?�:/���ſ13_��w1�R����7�[�=�&��ҷ3��o���֮�nc����x�X�����X�0��DoU�X��J7��2I�Ș���|ɰx �f���o���a�}q��0�n�%������u�K0��n�B��X��4�0pzqe����&�R2�_!;Ʋ�X��-�Z9�t\1/����fr���E������~���~^�>�J�-2D�Ѡ�ȑ�
�J���Tj��+�X &س2 �6C49ĝWJf!)�^S�kY����ٜ�����R���Z��E��E���Rcz�K�;z҆��"$��;�/�'�4�.�  m՚�h�{"5g!ڞ{[� v���1�2���0z�]�
?�T�΃PȌ4�%��\u/h>����!?�?��Z��O�:�j�0m��{�'�h'������9�͍;�T�,����b�ﾻ�˂�V�8�Y)�Bg�q=#�Rh���bqB+4�EYԞ�1/�-�;���`8b��x8��JѮ�����+	���⣂��po�����%*�{�w �!���:	�h�6R)� ·PôJ>�yEz��v��I����Ί2�Mv��y��
Go���-�h����������V"�d(i}�ڕC� ]��/_�U�!��Bq��d��"��N��r6a
��E��h���$≔5F�.�Hp��9/�S;J���ؼ���8CV0@��*7}�M[q����]{S�P���-%��ћp��J����Z���@�LA��y�`����TY�E��ho��E�SQ��?2k�CN�)!
*M"�Eu䍉-����Q7��&d�  ����ѯ�dՔq�[�Ӈ�!�'�n<$�5H�턧K�&۳�<՝�<���G���`�: F�	5`��/XJd�C���Zէ�V
HTj�V+�+x~�<�R���{�l��K��خo�6Ҽiӈp�n�یdd� 
&��[��kҨK� E&5�H44��o�0W���+שN�jPH  B4���E�����#1��Xэ"�����`=u�z������mp��n7�s
CM�}r�(���yl�;�!��(�%��-�ڄ:������G��2�?Zf�O1�^,?�G��{I��$��c[@KN嶰��a�l�!���zn�jw�.�B��Y{Y&�W�˷��c��E#�6����=Ú�e��&D���������V�&�����G�.�C�����O0t]�׀�Z�>�2J略�����ɥ���`6¨i1o���E��
���u%��
r,�-����b���mŃ�]�����)�s�\i�(��R2>$UH�/d��x�9����[j0.R�P���S2�b̷9�4<���o�ن2y��1������9������~/k;~p�c�'��/:�7ϰR/O��W�Q����l>��� ��$��_�*�'��ح-]����&'���;xG{�g�|T&�  �@Q"�{X?�/Y>*]7Ux��V���r�/rb�2fjt�Ld�>1��f�w�m9qvy0[?2��h��/�fZ��f"N�4�/24�zA����8��$�>yO`A)0Zz@�0/�'�w�oz]疔�G	�H=�yg��G)0�Z�`
WX��V�-���6[n��t�}�G��Æ�a2d����6>e�W�#ax��'�q�ear7iz��ҜE���le�������Ɲ��xn�$��,:��"��Z�W���)�2";E���7��3W؊��,�q<��&;?ї�9A�"ҤX�qbE���C�8E��d��,w3����y��eG�a�Sv�;9��T����f��(S�)x�	&!mR���?�Bh����2[��vcu,�o�,&�f��wB�˼`��w�0�l�6	;���͊��J=��&m�;����3�`j(�����F�����ƛ)�ɇWĹ<d��
K~�e�ͼ��yx��\׷���<�����SG��m�#7$�������8:n?�{!.;�|l��l�xȳ���}�z�:!���+A[�"
2�ނ��{�8���ѐ$�hň�1����ވ�O�I$N�
�`u�
&"rP4\�;S8@�J���A����M7_Q�L�2M�Ɵ��6��'���8�����n�������/��>ۉ��1�M �U>����v�D��+�2���t�����?�\ztp�W�È��	ⶳ��.x"�~�qH��4�3ă{x�up��}3l����� ]��v2<:���WD�Q�O���f�:�'��8�Xఄ��s��ޘk��B�s��Phz���B�'��d���=�s���\�����>���1<��rO�bN��4=@���f8���5�1BF ��Q��{za�l�];�Ϭ��w�v3�;?{{�iB��|���j��?"��i�P�5�j�ߢSro8��e?��\���Q���H�o0��l�H�U���d�]j���Dt���N�_�[{$�&8a�j��������+Z<��>����d�G8[=����y
�P��&�H�۹�23��ܺ���5�)���gd�psԋj�g0�B]���
��}�)V���W�S�ރ��n����4�[ڐ-�r�L�0��s���e,�jG�'�r7i���G�]��9�o1��[W$f�z#�;615�B���;��*�z�McQ�3��ط�&F�[�Oa�M����OS��pB �_�.���N#�v�]}���;�^=I���p��c� ���,�kE�����\?�����(�8�R�Y���4"���@�D�p��)U�e���㮩�voMa��^�pr5$J�A���6��I���E���,+��� ʹ8��;�?E#���d>ga�*ݬ�yz�����O�BpR��Fq�@g�
��.o����B��%_z"s�'N�?-4�$�i��s!��#Z��S͖����m�ܖ���d��YC��\|xcW�l�C���%�'�K:��ㄶ0�ԁ"�YP��+(��R��g�̬M
i�	O�
�Y�M['�JI@j��:|�Oބ�Ž�u:�*?k�M@U������ir��(��uR��:��JEp+RND���0چ$)��O��ss	Z7�[ς�3"���C�o�	�D���'��I�~�!�?�@rQ�'��~D��AMj%�C�u�f�o��f����%hB���!Ԏ�=�JE݅\�Ҷn���nU����M�+ ��gʒR���f��͂t�����OR1%��ާ)�v��WL��T�"R?���-� �hUa��t6�����e8��IzV��
4��f(]�����>q�c���Yj:Y�C��L�� �I� ٪	{&�'�U�Lo�tW������6���� 	��y�	*�)���#|��K���AN8��`���~��}'��J;e��Q��b�<�٤*+�7O�k����%�0����Eoh�Pz`���5z@N�5��ʖ���c�b�*)�G`�'ݖ�ez�K����҅+�FY�p-/\�x>gҳ���ǽ�� ���؄�ֈh��^[:%�M�9�	g?���	FX��BW]*��0Qx]�"h��f�̳�(�/������1��ܘWe�t���*/: �
��4�Sˡ?���z�v��y��?gDJ[yk}���	+Ύ2�cIl4l����ħdE�������13%���iQ#�s��w�#�l%M,k�
I�o�j�{��n&��(X��qx2��P���C�d�fWB������h��h��*zQ�+�W3Q�Ѷh� Mv�����2kئ2y(8�����_�SQ�Zܢ|JM$��[�L*�`>��v<02�|D�H����FG��P������*��*�:)�	�S|ޕz��Ģ9�������o�x�o����f�O��<��:��vԟ��cG+*���I�(�gbABZ�5a]�:a��C�e�R�nY�2�\�O���_@l1��*:BO.R�P��Q �����`�hJHgwR=�Y�O�3��ЯM�y�J��mᗸ�^Dt{Ӿ� 2_�_�9I�j�N���Ҳ'��m�|qt�:+�'T<�����u"h��{�U���;>�t_0���"g9H�(��˄��aS��A��[{�{9�ۍ�#��,�N��vC�P\���\ �����M=�l��#��?v��!C�
�C�S�V���ʿӂ6@����q]h�H�M�ii�ٺ�m��-$ArmjS��I�U�×}�)�x� �Cy�)�;݈z�!H�]��&Sz�%���#8j�m�(��@nB&��mF�m�b������J�(͈�H��b�6���zv��;�[ɉ�K��E�5���Eh2���p9Ca���n���9�D�
Gs�qxS�~0~��=�8
�}n�rT�_Xe�Y���ŕ{�։��9�]�o��9�ٽ�עS�B��j�,s����Ld��0؆'�j	[�+�ӳ��11�00+����s�v.G���Fǜ&P���VI��m?�Z��8�&}�܎�Ɛ�D�I��/_�}&����-�9�9!�Z)��C�S�*,x#�U>;8w��T,����{Z�g%�� `_�����]L]�r�x2_� d��~D��}v a�2w�p��Hk,C���y��AP^�����]�og)��POpǃ]�m�ٺl�M+Q:��T����S 6�z��K@[��$ǅ*:pP��+�^3�Te+��"�j3C���v�x�����5F���֫�L�M�Jd��Ѥ삭�}<���(jƞ��d˅]������Q�5w��.�n[�a7n�l��� ��s>#�w=�v{M��@��°��]�C�UU��j�������y^;�'�4b�!*~�r���;Hߴ�H-�D?�������-b��#����M�5̢�����w��E�b�Ѡ�:[%��,�W��*/�4"�V����Y��-:��z&���x��?�b4JE�8���#�+h;t8�Q�k���H�^���;N!��1퀝�8�ˏ�yj^���T���e�>F �g
z]�N���e�V�.�ܖo!H5)R^Z�R�Q�䌥�P�>j��Q���^<V�RF���6y�j�'J �k0�v�M"�2�QB�[k@���F^�OgR��c:e�.Е���FQ~pȚ���|xi}��A"V��ӇZ:�`b���󬸉۞>lh�O�%���V6K�a�g¼lg_�%��y��C�j6{��78��r����%�������_��|�8sǳ���Q����w��T���������y���V��SP��T	s�,S����Y�hZ���l�/Ljw�L뷖����e^pyQț3Y��e��mA�e�o8�+Ƃ!��:�ȯK��j>WO�#���גK�yzpMEA-Vy�}l��U����=!�GT����*U8��{"�z�r�=��lp��e|j�ц�}�����pc6TU6�������3�6��ݜ�X�
��P��hQ�wl�ŗ�ٖ�x�'��K׫)$��-�.{ӛ6*I(���r�����$uFj��-�B{'�⬚�s��fT�k�m�acҏN$���B�ۿ�N�}W���Ѵ]���;�+�Lk}������.c���-��Rm^�~���e��+R�K�K������	
���M��{�x�?U���ثbx"GJ�V9��B�艔|�ȗudT��7�#@�V�\�FN���rI 0�l��Vj<5��*�|P~F�li/}�bI�*\k���#+�����Q�����n�9р��{Q�LIׅ��}�	�4�z,�sA��.>���ٍ4S����ew�!@���TG>_o��{;!y.]��=j�WF��	�@M���b���:�ǟ�UEP?�7��  �{N��� ��W*Y� A�n9�o��L���v�!Ee�خ,3}���C�Z�r#�7uo瘮z�0$$00�vu�U��LV�����݇!��ԗ}}��J?��<C��>����N|�&Q)�=��l�~ir�͵��ƺq�K0��0�19�8��%!|��镼���^����A��5��L-�A����O�A����7��R���U�vW	_�0���Oz�-�șrb��qGYHT�lW�i��(��D�\k�Y��*PF��*��~o�X���,!�mR�MGOj�}N���)=���TS(���M�r"4@/CA7}���Yޥ ���c��N��#-e�Ž2�<~���YB�C���8�2�/�R�>�	,� %�#��J1��j����4�ݴ�e�31�����m��Y�)Բmc�$�:�*��6��#�Lkj�]�j�I+Ud�^��X��A,Е�,�:Xΰ �>,j6|�,��+So�c�͢���[���đBT��Rt�(��>�˝Qp��Iܗ�9���pH���b����f�?d�<%a�Y�MpHɐXh���pݟ���ª�旝h��^Ꜽ�Ϻ֠�aWI��6�y-���y4:ﵰ7�u]�δ{�r^��eT�؈���W�X[�Q�M�� �����K���
Ilk��@<#�����C>��m�������Sؼ��d[e`c�і>G9kc��)�TC$�N�;=�.Г���J����d�U�Q+	�#�H%�}�m���w���$7R��Yc�jH��_�s�[bU��ΣB3RQ�<���h�9� �R�Lsb#V|ܓB��Mf�����������ۋwp��u:�":"�BI�c[!LQ��_B���ff��-/���
�GY�ȧ�z%$Ɓ6�Ċ[
F�^։5�1c����Q�N��E*
R d:�6��P��;: �o�Tǲn��`}A�
����]jf�.Ig��^8bn�2��
�	>���CfTۭ�J����<"2��#�^j�L��Rk��0|���+ӰJ)��r��NT����tV��5�*�isᤷp��a�a��͏I���n�8o������v���WG�ѻ���y�W��V��j�eޘ��UK9:��ޝ^9�:Ϋ�d�rE��ƈ=4�����}Oz%%�F.��+x��F���(��F</�!;�?��l\yB�� ;�[T�M��|�Ck���l��m+u+������Z\��H#K���՘-�lBd�A���,� ~�/X��I�M
��8��ѦtCD!a��{��ȸ�J.�H�.�ܰ�w�~�񴣳c�U��,��N1~$j'K� >�E\ߍ��)S6��]Z��g;� ��m�m����l��\���t ���/2��~<�s)�(KMc��xA��([$7XM��WfL'�{�ɕP�a�O�Y-e�h��ua�_�8J�nm� q��vX���^~Y/T�*����<[��2>)����a~4vO�դ��F��vv�S�`�{��l^�h�y�Z�����7e�8�{ХxP��j��u{V��)�_nW9��X��P&&o��ߋ�P�q,ʲ�*�wDU�e*�3^8�؈
Ff�5c�N�;�_���M,�F��ۧ��-��tS�yX�����V���6l��(��^5���%����4E�b�ݺ�{�`ĉ�Q/~��1k��|���?(l��}��̾b�!g`�4T�8������!����&���1���蘍�x�| r1�p�S4�6o:n�TZ�. ���k~��i� �r)E����k������O�{\��'Ӝ��Z�f�6�0_�h����)r�D��.�g(�z��g�@�؛5��4Q�3��]G�S�AR�Yk�2����u�K�A�4�D�r{�&�q�1�D��}b�ʧ�ZK�E�5 �lxә��n���<2ǳi�2"�;��-�X�_@��m���F�W�Z�H���~L��77��վ��2�l�nr��m��[�a�m����"���X�V5T�*�a�O���z���bι9J�C�8��=���zK�jB���ZYBνX9>ZW� U�/�<�_X���V疮�q��g����������=a���&f�uo���=�^��]7�L�D��N�ԠR�����;G�3 3�/	P
ŮLD����"h���'�v�3ޫ���-g��;�����u��f�e��X��CU�"0��C~�̉��x []�<�m*k����7pb
���v%������n��\V�$t飡46�8��1n��.�\msd����3W��÷���u�oC������"ƒ\�YLR��K�.ď�c����)j'C���me�թ�g��3Go^W�/->ͽ�f����e�$��t
�eY`OD?��U�mɢ����PN�76�R�qB#>�C����J&&�1Y7*�l�HH����B� -�>ޯĭ��9"��d�����^Gȕ1����K����w���c����?�י
!�/�Ɨ��\�c_jŤW��D5�������u���d�F-���2	o��j俕�h��,��#��V@!��̫A������3%\s�T�.��zw���$,�l{�Y
M�}��Yg���un,Cx�� �s=��#{N��J�9Y�����b���:�.b���[>�K�fD�Bn}���6q��4eq�-%�iKB/r�V�U3J�B0r�j���pX$?�+�/�4���n{����4�����x����a3)?.� ٳHҳ�wU`j�	�S����7��2�h��/r�L�o��ƒ����AU���o���[izA�����k�' �^�U"�%� ��������5�3}�O�t��T7>C��?������jm�������~]�-ߵ/�mԏ���j�,D�ԅ��SX���N��m鹏��TE7��l��h#�,�w�&���GUiӋ���a�S^Ԟ5�U�,V�)�|PI���HO���q�6��@hT���v\�C���q����@Zo2r� �:`)�o�J�Z
끁k��W�Dp����<L����k�X��k�B��
�:^�o�f����q��A��ѳMvHڲ+s����F$3��C�=L��fm�b����T�Kz�8�B��*D�1�h:�I+
u����煜�Ӛh�m�K�)z<U�MPt2�h=�:.)p�nA6&6��ꞧ-��^l	�`�
���,�4���٭����XT������ Q���c[�h.�tO.�*zWY�*Bf�J�2�4#�C�J/�Dg�oh�L�c��o�D D�� ��Du!�Ɨ�E��C��/6�8;u�^� 糝G ��i����z�F�$���	w�>0-ǶF���8#�Ų�s�RD�S��v˪_ץ�?$ç~�b���"ī���,y�'��0e�E����6q�O�r���g��-9��;4�'��hg��7��zM%X"�ԍ4ml�<����s	��(o�������}!�@����}���w�^`r�];ߴb9D�;xտ�� md%K#�X^�H����D�F�[���zBa��;�r6�y�Ȁ��M�Y�#>��Oh3I�P����o�k�����	�vw5_�Z���i>������&K�L?k��
���P�}-�o%�P*C�����l�A���&0 '����H"t�1/�a+Ťqzc۽@Ҍ�2'�4D@�ʪ��ֽ�a�T�[;�D�����s�h�%�����,�jv�e��@����ae��B���C�~�^������2��D����O��Yz��V�@V�݈�Hi��e�����Ț�6q�#�����zԢ:t�,�Ȋʃ�Q�:�G�n'=fb͊}F0�&�`0A�\h�wۘ����1��L]�d�8��,'��Ͻ�*�OwN���^�Jg�n_)ف����f�&�a�JYe���!�X�����w<��E��X�{ �+��&?u^��H�U�یp�(��Bϖ^�d�8{��+���Ӳ U2��G��]��
T��g<O>�-;Lys�7cj���(<0~�V j���M�E�dMC,ɍ��ޔ�����'�Q��	����g��6�1�+U6�U�>ٓ����Qp�gr�Fr2�6�o6g�l�D�:�v�̃t6�ؤ��c��k΋�6��[Y`�z�|�i)
>��D���J~|[�Y���\'���"�I)�R�
�ҩ�xM^�Z{�T<'q�界%�Ǯқ1@8��?\��'L�F��M]���lW��W]��qd��"��M�W%��k�a�gC-08�t���Dм��PڦoK����n��-�/2/9��V�#�Ec���/^4%�qP��KJ�O^�8WB5�
d��`xI��������i�PH�~�����~��6b)k�V/�T3#�
��r��>Zk��I��v����=
���hW�
�a��	���Q{n�����eA���`�zfhm\#�-P�!��������5l?W|P��k���@{?��O0�d���
!/���z*h�ǓC7�z2��)l�`}�a�$h{X�W3������,���8��`T�#�_�� �����=���Ġ�H�3����Mu���$��k%�{´�y�g��>�I���x�NFB�Oo���h/	�F�XN�ʚL,}c��%��ϰ�`t�1��ڝ>9B��2����tHo���J�.���Cl�8���g��cn|����`��//�	+��?�4.�%�<<h�>�Z@{hv�dX� �����*�����MY;�H���GW�Ƽ7���Fk�B?K��z�`b��a��mjI��0��؎�!Bp0�h�� �X��z����rk7MS�]�A�g�Q+�W��,_a\~V|/>���Ǝ"%CM,��1e=H�-j<J@�a����W���r�6<N��ǅ��Hq"�ؠs+2R%��3?�Sd ��~���ۭl�^T�[���\Y/�5����7i8���|�k��ߥ�rY�Ѓo�a���D�d�
'\{�;�s��I�#�6'��R��� �,��$[��%�!ں��Ln,/ܙ(��d��<\���(P�+���\�$��QJ�Q'z;�#L��mct/7����7/*X�hO�����tK��U�G��(�������Q�����_�u�n�askW�ͼ9�l�q/��`�ϥ�C�s];MXha�S����{�U���
���II<O�����ޡO�M񅠣=B27�3}rG�`d��A^��8l����'�t�f`��;O�N�%$���k��N�*��v.n�ӷ���$�K^X��/>��8�X�u��*�T��R�z���݀�ݒi�+����P���a��S���@(X3���L4ې��:��Y����\�����k{�"/��������Y*K5Ćʍ���ͿN7n{j*8a��K�ي��V���).�������g�t����uX��ƭ���{�h�	�Լc�3=���H��.�Ug+<��4��b���GI��g�5|[��ּ�99M�~�U����+�ۑ=:3�st��<٘?u�<��toi�
�{@�9�8������J!0�E� L�܂7KZ?G�����B�a���tp��f�~��6�6��f,ml	c9�~)3���O�i wi���j� �!�/����(^+ռ�ţ�h��p�(>͞�gc�s��K ���U�xi�>Z���������h֏�Ee�~���eXҙC׸���&�K{�)�$�k�7�>!K�m�k��p�R��޷�-$�/a�5���W/)l�z�:�{&�W���.ݔx��=6mQ2��H�ѳ=��Qm_�6#k�-�&���#2@�K�3�� O�qX����p+E�a����yb�0�����%�Js䋀t������)���J�܏B��w�k�q�[�Gp�_���@��'�vm{�zLbIQ)��rP�gKb��+а��(�i�s>�[��ì�񩝥ʍ=�������!D���!��[Ģ��U#�?�>ʬ:��p�(�@���������6�����c���3�VkOI�smp�<���h�=��om�8�!�5�G�N�F} z¾e#<�5
^28D������H��Z�x�x�+$���	(��������ܝ,&zN0#G�5�f�����=Q�׿(g����Q�kPD�f�&���c�5��(�2s�`��>3��	 ���b
+�a�(N�zSi�(f��:�;�TwJ�)��7������dw�#�8�u�#��Ͻ�q
��B+"_j&gY�@�t�&�����Z�Z�l��ùa�~�����C�"��x[(��������
�*$��"ҧ�k���H��3�x� M�%�5Ϳ~9t��^��좋]"+���`?�������2I9�l���މ	p�ڢ~��ɱ��C}�rK�a��ka�����1:���o����z�$�H����$��ݍ�1����{�Z�e�:��v�I'�]��%��m&���/��3�f&eׂ/���t�GuR��x�,_$-
R{��G�� �n�����Bg�g�Ǉϒ#7304���Dx��m�K�Ӌ�):	��Si=��i��D�Q|t�N���
p����u�m�k"�Ta�Z�s"�&�d�0�!B�3�Q��A}`�p�[{��+o��Rc�gĤP�U�i�ر�9��?��Rᾙ������Ϸ\�$b����
��/|��n�{���%|\r\��老�q��ګu��~�f����Lz=4�o-��b9�`��*�.K���#4�[I^�Q>쌐��U�;~����L.�W�ïpq�a�"@�>�4��^��ζ���͒����'�#?��(���Jڄ6!�b�j5�S��lZ]_%�6�>Ž?
D̢kO��3h�8��z��4$�4��g_B2�P���2�����D��ٚ��TB���P��J���n�嶬�ޤ�����u�5])���+$���q��VY�x���S�z`V�V��E4���]s�h��:[��Ęǥ,6��s�X~��Q���]4��VsW�[�̈́���>���#��?OtT���y~F0C��eL�w���֍��hD4�#�5BV��2�~�%(/�Wt�G�cΧ�D���C�A��Ҋ~|��	V����t9�<6�VT���'���?�Z�W�B��9���0��G�ꊆ�e��������o�?sO��w��.&h��8X�)�:
���'N�FoʋmJ�BXÎ�p�ه�(O����+6X+�9�)��7ca����Jy��2Ώ���PA�OL�|�0J��K�V@t1�ޕ+���h-WoGD�g�x�XN�B�+��H���?�n���8\�*�ÿ�?�<q�b7�h0\��7"�zw���N�K�6��wh��|���N��Ⱥ��L�̯����[�D��e~�f����5,��| ᵥ0vj���.&i�3��*����Z��}��Qoئ�(:>��n�/%YD���"����Y_��S�|�ڙ��FŲ�(�XS���_��� -Q�,��ٕ�`'l�:v���mAa�)��15	��B�|`��F����G�q�D��:��vř����������*��l+�ҪT�W1�o�,�E�¿;Hp~)����)SD䯐��E����:q�G�W����vPR�c�t��]��Y4��Cj'�aKj�+R$�Ǔ ���<�$��9�6\��F��v�_P�nz�R��牐����%���A������q�#�t����;�:p~uy�>�s�	;<��C�0+�~�}%PߋL��Y��:����=�>!=�����`>^F|��9C�׻����
nq���_���X��I6��ۃ�ش��o����e]�E�Ym�=
��!��B��f���"����5�,�L�}�r��N��%]N��[�Aw�* u������q���Π���e�*��b�x�b�� �X�9���{
�\�� ���J���?V�vQ@4�8t�&ۚȌBG�QTH��b��w��J���������9J�_A�]ʅRʥ,a/7t?W��-���u��FK�跹��V��M��Q�ڃ�R �up,�R��W���|�&K���@s1]��U�N�4�8��/:�^��s�۲�Eb��D�;q�I������W�
�|JU;����s��cl!��EB�o����R��2�p���?CQG7l~�a�1(����VR�Y��ZḔh:�{1�y���{D���>#�]�Y?/��r���Tַ��]}ǥXa� �o_�B��_-x�xG��5���� s�ugNY�}��E�	� �_p]�?��u��ˆώ��$�}VJ����%�H�p< ��ۢ�P'm����n��]��&�b��sx&q.��!% �"+� .��"|��{|���mJ6)t7Q�V)�kΛ�2Ϩ�LR�_���򋯫�:ϧ�?g���!���i�&?����y�m���7|����e�L�Bu�l�֏���sX�!�/���#]!����J�-�9m��.�E���l��V_I�q.�����@��3���k��J�n-����-�P���
�X2jK�"( ?��h��Z�NMK��Ɩ�NA��������5�D��'ř�kP<�6])VihDV�WV���O61SvQ-�X2�_m���o�ĵҟU�T"�2 u\�r�7<J�K�0n1�ܤiZ���j3�O2Y�++��l��%J��u��Ik�^A��Ŀ�i<�A��q�Q��*�D���^HQM]@�1:W���l��^��P\���m�V�e𗫕ڪ�צ�bV)����w�4��eٿ�g*���7tXD���Z|F:�k���	��h�,S��Wrum�r�� 9Luv.`��_z"�m�8�u��(<���Z_���i�r�����·������>�"t��1R�(��c���5�H���a1�ʛ��Z�(V�IC�[�����\}��T;L��D���8��ua�CH����GW{5�rҲ�����?F%����׆ �ZѧU�&p3��ٗcZ�d�Da�E�Җ�&s�-���`r�Gc��Ϛ�X"p�؛����6p��U_�j�a#��;�3?�w&��9�fL�0¼����PCkVl��<��2��?����T��?[��%�2�r<������z$�-X�j�x�\�lw3Ȧ�=s��$ſF�F��0�B��Ӿo.�=&���-ʴ�H���}�Ĥ�iv�t�]�N���+%�3�14j�)��F�?�]�̍&`�W�V��¹�e�^eGX| ��K�+�k~i�KJH�PԵ��L�̌:W�A���| e�h����kn����q������-c�jU;D��ȠZȕ��i}������8\���R%�1�~�33����!�3�v���3u

<�iZ�,���K!�V�s���M>�&�y�h2�BPhZ#cȍP�����t*~�|�Pp����Ip��|�(����l�e(&4�������x^��L��zl�]!�xA⬋���56	B��u�E�Ua�鲪��hHN\y�]�F,{�u��b�cj��`tLm"���Bha�=(�����\��B��1b�o�tTB�Sxba�[C�x����K�g�GO����/�8n�-d@S�}�E��U5=^�/Z���^�^|��"�+g~�]��"�I��r��VK��\IX��;ۇ�hĩN�xc�	"w5z���c]n�Mz�x��aC��J?�2޹�V.�E�1k���I���Pu߲ ���;����$�t�R/o��� +|%<�?���&{�:fqW�rP�g"/JD��lIzB��Xk \@偐d0> ���ܲ�nRo�Q�.v����gL���!gL��:\��f[��n��׺�6�*�?l����RåbM�[J8q��7$�C�ͤ�)��l�X�gy�K�U�:�QÛ#��D�0mq���ꩼ?�p	�Yل�^�ڌ���:ۡ�
1�t�XT�oEr=�RL�����_�C
4�&�ڧ��?p->���Y8�DNċ�
���Kc���L(�-,�Kx�ʁ_���=/KB�S�*�7��4���KF��hK�&��a�>uj$���/N�ٶ��
��ǒ,�ݱ�w��Iا5�Ѐ�+Z�������Ldg6��t7��������^�'���uY��8�78t�i�"wg�8h��O���~����$c�o��s�0�s�ߙ0�E^@j�5��_�J�+��K�R�^��S�M����L����nՐ�`����吪7&�aty�"�tG�L���e6�G��h��_P#�� �j6ޙ�ᚎ5���;i:�yJ�'���II�<S�ңW@>�g>i�-�w�?	H�Mz�W�^��r����Ws�����
@ ��B;QG��:���8���z���O��ZDR�Aǰ��B�M:?�v��)n&�
����˟u8����.���Ȍ� a��҃w�U`�@�&N�C�[|3�FǺ��+�_W�����	m��B~�$`3>LЌ,Xת�Iu񁗒|ܖ�����~?ܹȯ�&KC�Wu���,|'���2	���U�^��;�u����er�]�L���ve!fϧ�P8��,	,-�{U��ńj�)7:p�V>�G�畬+�Kj�|��Z �t
�W�����~�r�/R���K9���e~F}�{�+9�^�Q.Ov(��jdB�)
���i�V�!p{&T4��Z�ݎC��"u��s1ݻJw0�zmy硯��,^�{?,�b���+����5���~x5.�\;�j�`0��?��1Zr�[HJ���v.���X��?�y��%���g��C�V4-	�?3�ڳ6yE/T� ���T�W�FjU����u���X��U1~���>���;P74%��9���h�<�@H8�h�x�^�_�4J,sY��1���\�ukZ�c5*��lg�u����2�JVL^C�n�[�Z�n�Ŵ��qG��5���`Oё�in
�����
s4��$���6eA�x��&А�@�0����?���S]�٩*�xo?�������1t:ii\��{xP��\�t��o�ʫ&�Gv����4ns��2�9-�9��?:�NQ�@0m�+q(�S���ތ&o,TH��@���l��<в����S�9.�%��iE*x���^,�v�g��oaĩe��FL�������c��^L��ھ������i��I2)�ڈjFX�T$�B�Q'0a�HC���A��%Fߝ���ej{���ǘաh�Ҕ6���+�xY;��ji�����á�-�;)M�� ) u��;l�[E��b��|	X�x��D?�=c
�ؖ]����Z��>r@�:h�$���}]Ï;���4so��$)��iw0��//���7r$n�R��H���sHa�6�Ãk��Q�>PT�¥+�s�(8�E�e�oU�6�+�Q �zCB~�/�I�n�����љA���X��L�VM�����sbo'�e_��]��5�����u�����T+a����A
�*�[>me�y&b$���1��cX��(��+��':K�pyx!{�
z�ʾ�0�q�?sÔ��H�ƽFQ��f��C��R����N�8����4jK���rJ|���<��ZK���<���R��6�4���24Y@WO�pu;����No������'��/��`���X�<�C.I�@�W�p����Q�Fӏ��Q{���ԾxR�FDN�lp�	ɡť�P�b��_�)�=|1L܁JO�;�o���$�xcsTNiPe�V	���(B_7� rv _�����܎����-����+� �;��T���GdM�9��Kk�U|�V�v��.��	"�NMh$Kk10Ҩ}L�ԾA��}�g���m��D�ͷ��Bԗ�뒷��Mt`hW�e*[�>����'���?��������;c�$U'��2�8�����x�sߴv�Y� �Y0��c��P������4xGz��`0���BT���t���Pϋ:��8iQ=������Iܙ@�!���L1��dR�z��g
-;!h��|��ei�1$)��CɗRLŴ�#��]�@A��"e��,*��-9Y����|`���ُ}+;���.��z�W_�����i��[��0�qQ*���OP�[��Y�)�X�CX�f��0�!Km��w�D�	���ٵN�����P����#�pt;�S��T��o�DC?�gMer.^�O	�YT�V�ϔ�h������-�o*!*�Y�</��*l�!T{��Da��R�]�6���)W�ED�t��[$Zs��G&T���Ue+0y��p�9+�<E��݄ۨ���xO��_��F_Z��<����O/��KM�+���{�yk����֯v���$�o�~w�F�N�.�J��谒fs�3��`�#:��Ʋ��؊߻���CI J�~LK�y_���@ɘ�)�_���mGZ}"G| lrI[�%Y6f�%���{��U�n�z�/���9O����m<:��׋�;������������5���R3�4�	�:f5�t�
%�(��	u:�T�Q� 
�t�OT�!5��%��D#-ة��NP���JH��O��G���ɞ���n܃S�D���2Ҥ}˭�����;q��1e{��?_���'پ}uh-9�m=���%�t����h>�Q'� S�Ϭ�C{ٳ�/M�%&����-�GI;鹿��¢�4�G������To�z^��c���M��0���=���e_)�:L��P�_8c�3Zr;y��~��lV�����o�|�ȡ��s�[y��Ÿ����b+�c�f���9�"[�N-lÂ.U�qE�����+5��F]�=
*Z'o.���dݼ�%N�H3�6;�g�kG��p��ۺ��yA���D?��!R e�y�q7��K�̶B�@�dЕl����jIw�L���9oU!�� ���#�1��=��	n��a�|~qC�����0��އo��O�#`�yuꅁ��ف�T,� ��MST$9�WTϣӺ�G8W��Ch����a�!N�$"��Q8Pg]�;�ɸVI3�
ߕ$*��4���>�O�aڌ*�N�ܱ{7��:��I[q4Ok�
�Mwљ������l	m� �L����j�1�u�E��ԆxU�����T>,A,��>��7�n�2��S�`��WJ蔍�]����S��!WyוD���ȴ<^�@]����Ja(��9��F�����w�����L�#��	B��#G`�N�Ur�]9�9�c�υ�� ��|�y���,�H*A]�b�k����W��F�5ǀ���U@���'0!���"^y��V�@��?I�
Ǫ݅s�#��(nS���iw?���������@�7������B�[棩	�uoP��"��C�5�VQ,�.Ebi��Rz���a��?�3y5�z���H{�,B����(kkrW�:��.�ܾ��ؘ0��l�W]D�Y�5�F�%��}m�\��$W�`�^�FU�Ag4�*�_��^T��Cn��iO͖����߸麕-�����ޝ���D¿AL��`]�� /gݐO�b"���*F4�n0�|M��;�*Q��M��y5�Mv*S�J9��?&%q� ,n�B��C7h�;�,�m�apt�+S�B��{�]R����kq�p&y�����K��2Fj���WÙ*2l��Mj�e).�ݰY,�d���O)�k`��gj�FJ:��}\C�T���jbbo	]&u/g����n��D�p�Y-9�Q`~x ��.j�[kwWW�ګѰ��Z6�;<�����0�%�޻�|��WY]����[}S��C�6�p�l���"��eQ]�@�y�"6��_kO�d)����n�(ll�N��h>�I�q�W��-��S��
�*J���bC�u��:��y:ACȑ>�bt���da)�ކ�y�T��s����*�)�"���T@�p�V@"��X��ψ�T�(�<����h�\i�RR�V��IX��n��~��
��&H��`���ܖL�N�
�jcu�IR�s��Y�*��0q��Z��t$�U�̛���_��w@��fp�B�u���zP�M�R�I�_�Ob�*p��E3Ps�hjVH���~��bw��${�����ɧ�W��s�8}�e����y,�raJ @��9�5��#����؟�0VըXh�)ۻ��q8@֭%�.��[�� G���T��. i��c6��dZ)W������M�@�+��f�s���0P��x��6�_B�$�%�>�g�vMŦۦT�{��ay
o��R�o���y�T�U?(� ̬��#O=~m��7�i����j�Ƶ�EE:�N|�˝`W<�R9?�L$~��&'OpqV�o/�������RJk75����'[A�E�0�fʏ�S��ǿ}�Q�Kr�����+�����<'͈㜮� �7~:k��c���ϵ�����:�8;lP"E'Cݨ/kxnC�u��]v�@Z�uG�Ǜ9���O2��i�e���;'QZa<�Q�'c��®���KK�n[��*q��ly�;���(�� 
�tU,u>��x�n.��K�U�%�CEYM>I#�v|G�urTKiJDNk�z��9Z�VK@���W���n�j9,�H�u0�[˭z�#�6�b�[k���0��k�f���f,�?�ohX�Վ��!VF�r��IoyKX�M�T�x� N��Y���(��LM�$��_�Q� OT=�,��2����{M���!�[���1�ob�Pv�����2����YG��컏�UM�A�@Z�ֳ�����=�V��:�F�	����"D����S��++on�����zLfV����-ϰ?�.Hy�\�
�d�Ťjg��F�����T�ʬ̝k�ؐ f����u'�љ��9�'}kV��i���K�a%y&��ɲ}k��rRe_2Fp��)\�k��W�š}�2wx-�Y��������E���2ϴ ���b�8
�j�E��pe"��x0ɋK��œ��yz��A�Y���~��� 8���b�ɡ���D�g�^���Z��K��US)�X�X��Β�18""�4|�
׏�.��#�B�'��"�S�$�������x.��	�
H'���=^�k<t�蠾�mC����%ة��yG�T>)�V��w��uӳ��\�*�K8�Vc8��/�:ǽ#h�8Da��-y%�=�-a'�Z�Y�����(��a�Ht0�� �������ZEMb��s��ĳ��*,�c���+��e���GG����$��� հ0�1���x�MVea�gB8dIt@W���Q�E�jy+�����[��=m��<Z�K�]�!g�¬�KwQ���,�N���L��m�;� �`[)����cjrƆ��u��+���c�ZXW�w(��o�ф9�ӊp�l̉Wm�/'�ٙn	iS�7p�g�a��S�-�I�O`�m̈́�� }o2Xq!�s\�:�q�g�&D.�0-M��R���H�z=q�R���?��#o|��h"k#1yU݋đe�2��]�Z�1�b՚d-G��7�eM�i��*PxS�{S
l�d��<0ȷ��c�|s
LCm�s�kͧ4��-'�{�X��-8��Z��S��1oF�>J�j��h��	@�����Aá8J4��0��F���6��q���B��Pk�V���GTa�O�b!
M�4}.���tY)�_Ǯ�D��D�v�0�i��F/cz���:��ϵ!���m���u noj+��w'��>Q�!^����-�VZ�&����`C�וCkI��hj'Jm�\�W�y��匿�/ŏc��c��T"�㗍�K4�H���d�Ԭ;���2XE���0� ���^�0vW�4�r������v��d��:�t!u-�ێ �U�n]�4u�B�	�&G{?FB�O�E�s-��>r[�H2{������Zد#��DtF�e.�^�/>��	���:�X��=�ԧҠz#:}��\�C6���
�y��e� $����G�o}�%=e���G2�>�J.^�����ت�{��q�������uJ$/���\���TcC�7�����eI]�N'[�*�#�ќ��Ygz����
������:��)�x���آd�X���es�?���%�깯
4�q��?p���C�j��Sx^��N���%@y��*�k�	�аx^�4�QƝ;���k��X���XZzT[-�;��)��Zd(^��<�1	�7�����|�lh�o�J��d.n��c-k�A�=TW�:3V�ҡ��r�I$�9'B2��پu��7�ϰ��3	"bǁY�����
��wz��DT�
�����F�cE���c�gn���y�9O.�
n�i��b�$X+ �8�RV`A�Ɩ�o� ���2Hkq1�	ٿ?wK���y��G';�+��C=������ǳ���E����Y|�S C�`o	o���e)�)y&R���ޢ[n�$�����gMY�no�s��%�a��{ɕ�N&,@LcL9]/�l�M��4�v���V:�P5t�$�}���NpE@+�A�~�U�$>���XBw�Z�c��P�q��Gq��D�Me��$���Q�Wy�����o�#����Fw���*�ڕ!�lG0;R�'>C�j��B�ħ��B�%�����Z�v�-��"����"�2'nӑ��B��:��q,�u���"�P��*0/.$m�H<$�WF�Pq�R9ᯜP�uC�K79�{|]܏�q��|M�I�bc����� �΄o^{K��B�L��"����7=/�+eu��*J�f�~����L�㭲�e_m)��+�ơA<'���C,�&��K�G�	�1~P�3.C���$�\�7O�Jb�e�ƹD��>��j(�>;��sK����we��)���_�]i��΋�s�(Nx�| Ĝ2±����ÌEbT2f ���T��n�$3i�,h˴�㫹I�p\(9b�)�K��T��q��<�5��;�/�r´�.	=Z���Z������V��եr�I��7Q���%C.	�2���8]b��iDzD�Jkֻ�J�狑�����7��}j�y�Y�#�)9Fp2yEwAHa����٭�1Q�����O�Ȫ��;�@�C�֊A�-I�3�EqG��SL���h�?l�P��+��b�H6pr�bW��`�j�N�M�R�C��r�Jy��A'섵���c-Ƴ�(	vHS�V���<��@��G��Q׻1����&K�|4Gq�A;�f���}\���O㵗�U��ɕz� iBg&Fr�0�~7Ol*5�I_尲h4G���n��tꌯ:�����8���/`�s�u�G
����(���M^-�+�$�y%.7 �;]SY+:���}��c�t
����đF�=�c��e<�����c ���K�5�@t�������K*�f*�MB��[#z��f���KH��39q���#�#��z�K^ʀn��`�5��V��Y�e��%}똛�.@n~dI�a�=�ϯpz�{N��#�EY�*����*�AXД��f$.�R��R��H�s���Va��9�F��-��nO�����VC�p���角<]-+��}��?��+�a	�����h�C��pk(w̸�]�8��q)w�aw�"�ab_��Ɗ�|$O�pS �<s�s��h����j��@Ɲ��D�=��>z[i�>����&2�=���}�Z};�j�6:��J &�l� C&���Z��xY�H�d��1d�Vr#�˥T��B�o�+��E
���܂�^oS^��kT�.�韔��۟��
��J�Fc*��o�w^��DN����V�m!w���%T�?M�Xģ�9���/�&sIƓ]tO�v�nT|c�H���A2&��?�%n�k�\� �ը]������ ��]�����!ŚO��w�\p���������u[��D@�W���w���O'ᯄ+
�
?�R�@�o���w�ǥ7B^������%j⃙?9�!H}����bl�RI�d�"3+@]��8wȬ����%0ɰ��ޢ�m����H�
��WTQ��VG�(���tQ�co֕/Y�$���,�)��������"`���>2��￵����x���D���ޭ�ͰQL��0� %�랡lxī�C�O���ah�/'{	fք����_�x!W���G��F��I~������#_m0�x��(���h����Y�ɬ�b؎B,?y�\�0�����X�������W�m	�,�3s������s���3�zx�d�np��xF�F[�gȞ��3ф��QYɠ��7��l��]J�?��7$���QB!�|$�ۀ�a�lh�PqG���`�̑2�r���H�܀���X�)�ש�^��V>�~Vq�82��.'[�2���zp���aM:јo5��_8��J� �������C���v���]���a���]o���' �m�n��fh�QK�'��������\��9]�K%�������rM�ʂU�h����"$Z?�ِ�T4�B�g�w,NcU��Q�#�r�{�ʡ�~P���R�&�[�t�����V&.I�s=EQJ M� ��G��/���w4��(�Ax����!}�j��˸��>������q��Nd&v�3�HX��h�|���� U�e�)��Rr~FNv~�n��w�wS�["�c�1�!�?�VL�D���R�V-����q��v�s!b#)�����S�6�uZd	ڴ��쑌�H-��.͏�¾����Aˊ��+�Y��q8�{x2RC}�Z@P��Xd,�N�}�@��ؙ���[�0�4h�&ׄ_y�6+��Z-/�`�z�16�����Ё�]H�9���fx§<��b��,�QjY���<z���Zͩ|��w!�ڳ��>scB�E�����|TM�����J_�$��"��{��dp[��/�-�Ǻ�d�A+��(EG*)J|	�![D:��7���;�c���,�t�r���Sˁ����p��0�1^�w\ m��.TGP#�9�X%9_��>:��{�"\t"Y�+�K���*��(�h.��s��ڋ=�
+fϓ_�3-Z���+z��ޛ����"=N�dnbX��,U�vQS.y��ꊖ3�YuO�⶚���z����mi ���]\O���;u����T]L��1�,�I�w�<�g�s8y��)Q���I��;�L�>�0O����e�K��v�f���SQ�<�qvgx���U�)��d����/����-�m��G����X������+?i��U���6;8���PRG���~Vi�&*����S���-�1z��ˣ`fv c�-�1��(��@e�7�Я[M���ͭPH�R&h'e��|��+�>�D)��i����P��(�?��>vѹ��(V�(eY��Ѷ�>~��qz3A�EB�Ҟ-E�@
�R���g}��sH��E$G���G��>pM��O�ޠ�E���Qj3��I��yn�r(�$!�'�b:17o	Ÿ�}B�%��~���U[��ꮃ��f�Fi "��e;��gKr1`RPW0��9���
���c�D;���]��#�WkͰ���s�uT��-��������pO�d¾�S��g
o?z�C����X�^��wu���㑝����?����{�G�����%��ڱ���H��F�/�7>�
�����0b
wMc�*�Z%i��>�l�T+U�R$��]v�y4���%�Js����G���w�ϴ;b��JKͨ�/��7��$qi� b�}MG�i��[N�trm(H1�u@���M���pȪ\�VM��kf��G�B�����ݶ�#�a���g71�7�۶�ܱ�h��ky(��S����0���n8�K����k���u?'ЇY� !�I	�E�!���}�B�����i|�DX�{����t�,�<Kc����\��(��Ie���/���~��MTw\��'sC�E�d��NA��Vz�9̑8��iu� ��<��<E����+�>"�P����S�0�{��z�l�l.�����e�L6g�^��<��,̜�h��B�=�n=�?HR��e�ڝ�����U�h�\5w�rE�� �����b�Q	z`dv�Y4�#/'u*d�nfD���Nt^����-��"� �b@
�x�}I;�Էy� �'���@����c��i�F�Z$�|Ü����ڟK$![��U��?$`!��R�h�3����=H8���}Z�9��r����n/��fw�F$>̄�ٝ|�_ws~VV�k����5�:�I\�E�}XJV�M0p��S6�H���x�&`~�Zθ#�J��Z�iN�f��Q`0_��u
��4���s�ў]Ԣy@U"d8��#d+R���X+j0I��W���)�J"�e���{���?�Y�h����Z�$�ރJ�zg�~��i�?uf�/�Q�4^Y�N/Ƹ��|(	d�%7*h��1]���j��C&�J8�CE;7�I��
ބ��a��8�5�d.O�.}6��Z&���J7Kmu=��1':�`|���;��o��B�+��p�2��$y�V1uق:Nӓ'�H^���[��s{>a6 �����r����H��r�K�����bM�pv����-�Ki�+��w��bѯ�э��u��_wm��'n�c�\������0	�G��E&�\�gk �Sb5��6{_�ݮ&`��9XH
'�m�3ST�����+��|�׋���~�AU���N���������D�.dBeUR��e���G[���)��vWD8�G���D�2��Y�;k��%�W�MH\����><��j0�kz��fe�C�~�1��-و�.q_#�����%怣Ů���܋�\7~�s�q��֧Mq�Y!�h��J�Ͼ!�ѫ� �郟yg�Oh�]�0���n��\P��U��`IS��uQ荧�[n7:��4Bz������yL�w�E$��&�8���r��S%m�n	!&���&��T�[�O��j�6��˃3�D�~β�v�������t��EY ���l�\��ċm^�K֨����=$$�����pW99]6���	�A1o$Hn��),��sn�ӵ ƥ�Gz�;�6�%�'[�j�e4E����t���_ry|�eJß�A^������+�b�nnI��I�S�x��W�r���JNZ�Ҫ��Z	J
;+���dS�����h6��$��/0�ڞ�Ұ�'�PdA��+�'�L� �$�6">zkxĢF���:�r�:֥���Ʃ���
l�P��[��/R�	L�)�={J�	��`#�j!��`�R�!�rf���ԓ�'W��SAg�pu]�ms7��qi�?�#f���D�[���j��"J��j�5Ux!i������!���L�I�L/՚<����'������Ѧq1CZ���i�]-I�|�a��Sl�����vo����T㎾�ƫɷ=/�#��ٷ 0|�������#�3����n���K&��{��-��I�����_Psq	��Ϣ�h��)[eEqw%����r��V�H��X��/J�FC�L�	< �y��G��_�*P��ud��eA�)WfK��������A�ɟ�^)��ѡ����wy�&>���'*Ηd�5c?�^o�^3�P��ٶw�8�B�3�TE�=�ʃ��G��7�>I��M���K�	�i�r	�'ʺUм)��Q�ì�͞PZ��+�
��<=�j�$���J��>���*���Ŝ �W1�A�Ǘ������kl0*���4ُ�L�����w��.���c�3/<��a¥X��y�ꋓT��֥o8X��
+�����NOM�E><E�q�z�=�O��΄�q�wáG�<��L�;���l*:r?Į,��j.ǵ5\�G�.�Ѩ��C�C� ܬ��<��3k#$���@��"��W�/v�c�^f������U��s��Bk}����D:�eAr��9t4�*�i�ψ��t��o4�Q����:�C�/{��*�ej9����n}m�'�A���I��d�7�lUcj�b_k���OοC�UF4�Lp؅'q��$4�kA�����rg\M���*Ή�ޏ��aJ�����4u5�.�.�) 94�H�D�_cG�VC�0��OzU�>om���c8L�C��[f �/�'s��}�
�thb�<+�����J`y;B �YC�)�:���X�&�w��-i�����˿L-<]�����KyJҿ�[�/yV��I���w�`6_Oܡ�|53���<T!Հ����&�{|�0 �B��Ӛ�R�[�b�5����̖�"��]Z܋��I��嬠�r���4���r�1�b۬�qn�&ͮ=�Ɇ�E�4n�W$�u3���B���B�����T� ˪���q{�<RW���hf�e���Z$O�'�&�^�K�/�U�A�~�:�D�Pl����{~�E�0�iu5��\�!M\���ΡBQghQ�I5.ݠ#|�}E=���nj�$�"�F�&��T���KS�����e���T�12�z���a&׬`4J��'Ȍ�u�.1`�oTq���]��[n��Iu�۾���e�{�~��a0g	��87�}�����Dt����ցt�HP�ZY���l�U2��'�п�E
-;����IZ�����Y;ʶh���4?�x�8�`��]����},K\�~$��i>�LQ��=a�[!l�ɩ�7:��+��`���Ar�D���FE��pv��2|]�(%�\�unYj�eNI%�
~J:��b� �mJ˞h�" ���`GS}���L��ċ�W��{����c�R9i�.��̖�v����cx6�w�)\��=ҾUe#Ř�UePauY�
��N=����t_Dm쁥5v��J&��U3pb^ &���W�W�D_���T�	ص[�мsY�!���s�!���j��^h>0�?�XQAt b�%�b��0Jn��������j���)�̷�%1;N�D��� OjmP��ϓ�s*��3D��G`#)g�S�+����L"TV����ཆb~@�5?,S�!�A$P~502 �?�^�~0g�8*�	�^�7`��J�S�Z�����V�n��5EP4WɱQ�Q�q�x��ح���v��w%��8����r�	r稀���p0�儗05sB�|�q�/� �m��lU���NA����o�u�~έ����s8��7n-��d"�b\�i�-%�B�SX���� ,�g�r�wz�N�/�cG�7��� x�ד5g;�`�dY~Ij�-}4��{UI�~fh�Wq`�nc�{\�4R���ȳ=X�?��+��U�� 0�}9��1������M� 1�� �-t�I�)LA��~�������h�~u���̄ӛ�1�<�gCKJ��%R�q}�\�E��^jؐ�'b��,�X;����=�m��|�q�ܓ�"�0�W]AAN ��q�!�YH����ғ��E�V��8�uE��E݉�$�n�ݨ܍���0�'�Q�w�ӧ�#8+�*���M�9?�n��í���+mnBG��w�|��}�t�;�e��}2�}8@��a��fA��B�-�E-HE���-��"�SuO����K3��3M�`�J�k�|�Z�Y6�ȁ�i]�TS���οO���+�Im2��e�"����6
��X�r`-3|�����N\i��f �P����I0�o�H)�d7��s��u�̡	z�uc"�,!nΝ���ǋ�|*t<����O�?{^�#h5���n	0�#1HV*r[hJ��u���Z:bX5Z-k�_��(����m]���}:���-1�i�8�	��\�}���4=��E�	h��2�H?C7c���o�t���˶���������Ay�M�Ô��w���f�d1�������W���偻�=5�sΏ?g�K'���YF~�4�ղS��֚��y	��4�e5.����-t� 
NVi�R���@��\rb��P}�8���d��W>�K}pU�;�S6$�E3XW=Cԇz)8R_`���"J4��3��\tu�=���/G�3l���+�u�#�l�8�d*�fB�����hg��r�!^~Q]��K3o=ȃ{O���q~З+��h��x��[Wft��l� ��3�)��'����	����d�����} �G�ј���nQ��}�f�K�D� ��uP�+4��ï,���Թj��0���k)���M_��<r�>ʍ��u��}a)�eY*�c��]3��{^z������k���|N�k��\B����0]���%�����˟w:"��A(Q]z��r ���DR\�T�I�X٧L��y�\ų�=���Pe81�����_6y��D!�5��*`o}c�Uqx�}��m�J��B!
�K��)��1g�"n̓���"�kJR�g����UR��d(�!C­H���1�+��Tk7e��_��q�b�>�NOXl���זN�������\�AV ��	����R�%;�V�`3�d��%Iw�J�/��P�'�GZ�[���@�aeᒧz����^��˞p�֑��@Х(#���u���p��ݞJ_�C Ý;i��6�-���e�o�u�*HԹ&�h�l�Ĉo�����hԝ������F֭M4Lu�k��m35���ߵ�o�y� �AY�z�S�Ր�6J.��4���[M
����7���BWDP~`����sT�^��q#���C'���h�zP�!`߂�����uHwp	�i9��+^L&8�#�Pr[dߏ�T���b��2bg�b��"����WwX@�
�ť��c��ʯ���?wK�Ǵ��t���.�[�^��QU���&��/~z�|�S-���d�	I��G�3�Ql������ey̾##V�(?��G�ܩ�b~���ȃ����f�,/1�DC�~5ۺ�T��g�\W��U�>�Ȍ_k�ْe�1D_$��V	u}[�1R��m�c����{Z�u��rl�]��xȞ4���9�.��聢�����������_ �k �K�_�ސ�T�wJ�x��+�pPd�e��fYvkD���4���&�ɝ �CYeJ"�#�r��X�bM�QyRmM��~�hC=�%��@�Ք�f�x����Q�k� �^	��OT[|��͘a��0���7Ц��Vk�ߦ�mݥm}f�q���J�Y���ܷԍi/��čس�$Ks�5H#�k�`Ӄ���!4�=H]�O���a4�ˮQ݈���0|���7(z���
�?���T"�� �X�!�Nw��t[��Å���`�s� '޾�o�x�n�e��]�n��$Rn�>� w�)AC:,,tu�T�}HR���5q3$7��~ͼ,+�NF��:*�h�;R"��;�^"�r P}�����h�c�~fc��0�?x�8�`XgY�{6�_�����u���e����][v�����a�G �'cv�*�p�e�����6�+��(�X�ɟ[�ZM����8�E�R����6s�lT�&p_ɻ%K!��Ć�K��n@'�\�|/nZ����j�q��.�̞1�"���R_�!~���[��:ȟ��T/��-�Vh��$�wU���e�^���ik޹�j|�#r�47R5��Y��^��(��w}��`��wG��0�T14��� q�ldA*�B#Kn����lZ��>�J�����~x�9��[��G-�9�)�5��}���/���[��a֚+���R	�d��@�:7�����r1���!~)xrۆ�L���񾒡�تc�:�j�rP�R3Z��TG����W��:�ۅ�����-ؖw#p;�XMmI���R�hk�J乤{7xYM��0lB���_�a}�F̠r�)�� ��8 �AمԴe����W�!'��\l�Q��o^.·Nuy�/��b��_{�$ڑ�sOǸ]@�����~�Se�L��}�<T.��tZ��l�J>�v+��;R�p��1�c����kQ>&��:u�(,�_�t>p�^Jw[t�[i��x�R�% �����3S�x�����܊���&!+��ZW"����z������2����c߿�v�d�JOP�k�i�(/�Һ�tΕ_�����2��7:;jN<�#	�!b�>�ҽE��^v���y,X��\��Q�|��tă�!�����D8($�K��;4Qhڸ��i?}����������34��cU��?X|0��8%��%����z�V�h|�Mw<8� �+m�N�3	��$.��&;C�{�ڀ|�4:z��b�1.�����`��%�{�m�\������R$�<�Bѵ+��O������k8����ǍH
���(CD��t��iz�x����!����:`�L���ލ�W�|��
W�9�hA<W���.��5�H�_���AO�7/�I*���
%!�-�6.n�EP`��Q�f�z1�:��P�i�<W!���ꌘ|Ì��-��=z�1���k�9�VV�TtH?�����d i��>g�!%f<�ґ�,���:T#F�3�����](�#n}���yܺ��o�>3���ܓ�+�����E�%�� N�bd6���&2�A�T��[HH�t���LM��{}/�D�9ǀ��D�ae��R�W�R���Gb�vJI��T���wy�����9��xv1��s�QYhi�$^��N��B���1��ZBv̽�B�1�b�,3��Ğ%�kj�s�np{�}^�7z1�9� M+��04'l
`A�xj� Mg�#p��z[\�j��gќ�U.���@��
 X�F䌃�w�R3Z�;q���z��2�"r~��#�r��?<Ψ�v{%.��a��dT��(,@��~] ?�0z���L����"��;ֆ܏Mkq����	Bڎuo^�ndMarZ�k�b�hz�9"�i��9����O�E�W( ��o �@��JV !�V�5���=ȿz�
4�ϻ��rE�F��$#͢�p�lG������� `��`n��*�������2)��-E���@���x>�Hb�>�h�z!�a���G�6�ݐ�I^��6Q�w����l[�j�I����Ssf*b��{|���o6@(���<לlɇ�5�B�,�׵�nZQ��寵�XXH���?����y��������l��<}�&l���a
�G֬;_����>�AE�g�j���;���S���
&��i1.�Zht��Y	����N�6z�4�_$V�q����u�m{S��RP�k�J��4,�v��,����g�ӈv@��^s:�l��v����u<�����Xi������l�4�Nʏh�\�1�No�o�V|,(� �sF��?�KLx�C��G!��c����>	'�*+G�[,A��¥�0;��.����]ڀE�w����"��{���p���?3�]�S�*";T�vI�[����%�]�	��@2;UZ �A��>x���������!�1�8{�aaG޵@\�u{	��]�m����	����� L[�i*�B�&D�3}S�������SD�!{�  ݲ����:6�-�t��Q�z�����۬C[tW1w6A�����v�ựPh)��h�~%]�LT_���@۵��n�}�W�羏�#�����T���5�� �zl,pu���~K����V��Vl���o�AU!��_ՐF�!�iS8L3��>�Q�z-5�Bp��R��#�>"�4π����.�$��Uc��&�)���@m%�`�n����><����m�xú�nuç_�z88���$�)n��p]��ق��	В��`��.�a7,�!�\Y�����!�S��G[:�gd/�!V������R.G'��c�P ׺��>Ξ&]�GW����M���D�>����J/�v�{BMU5�b�R��F�(�g!��+|�Bryq,�w�R:��%�Z�� �mw�q9�댔W�o�1'�%լ84)	����f[�f��f�(�βDY'�&(Χ�(����h6u�-���^��o��R�����p�W����	j���0��"�����ض�X�Fj	�)h�d��ڞ�W�G蟮��s�}�Z��`����#h��)k���j��2��	�H�"�N�Pt<7�H��p|�.�?�<�@'?��Eӽ�P�vmJ/��6ن���'�zm|�B��IZ�	�]���q��>g��X�j�?�ϵQXo�D�g��n��T��i_�x�6�Ңa�i[r�e�-+���C�X`�E
�Z���}��J��Yp�6�г��	X �T���D�����)��8����r�k�ꝲ��<?!�q��e���O�90>a����Տ����q��QD��.�`�T)��6�6N\����%�̄g�/�?[
��w߈��߄`�*V��0X~@0�������t�7r>�]�+ZE�t�1j��VԐfU}��`���$X���2:���jÂ�6�sb��y�=�>ab���X�R�ϭ?aȒ
$���0����P�6 �xb-00[تP,ڰ�:�Dn�5 �ʞ5�FA@{j30TF!����Ջ�f�
��l:�]�k)�r*��9��[��$� 9��&�˥��;��Jz�L'c~?e�U�/�!$��cPt)h�W��xG���UJ6�o_1reeڼb��Ou��-Q������e�M�XgNO����'��8�Ƒӆ�O,j���e.�z�iv�b+9Fso*��h��:�q���@Fe���"�h�2Y�>;)]%��~m	��Ҵ=��[�@���-/~\��:�Dpqp��/WS�,s��mBQ�������'�ǭ#s�t��Az����t�Wo?VH+r�7.����Yl��V��V-�t�֖���[Et������꿹����VQe54�v��a�V02f{�[jh� ���Ϋ�D�����V/�ʸJ6Z�af���~�h���p���.,�s���JӶ";�Qn"���������[�N��3� ��϶�'s���G��)Ɍ�;k�iX�gLb�U�Z����.9i�.DV���O��6�?��6U|����A��>�M�e�����=�t���/�[G�(p��o7�V[3�mb/¢S�7{΢�Y[�乱�](}�8,�\�2>�CJ�;%I��4�hb���s�W�ˣ��mWL�a�m��U8t
H�Y�R/5�H5��5��BU�:.��c�&���z��s�������1���[��e�T�z�Ye��z1��Y	u]0H�TSpC�π9.[`���N����<��-�UW6EF���l�ʝ�{��C��IYť���!P��q}#��^��0�i,�G�ea�fY㲷[dp�����ZӧS���#�j�.Ŵ��^�)Y��ڋ�YF.����ӏ�6@;_��Uo�SmQ��f�YUT#����;���ݘ���l@d� 9ru�f5�;MEUܳ^�^���8��i����v�K5��//���IZ��a��X���".�h���
�6�v��|#�&�}@��ř�&�Uй&��O�W��ϛX�>����߲B
!M��Qm�u䮟/�~4�?x��WX7�E\
O%	�$�?��O�\I��P�R�E�d��h*�I�uJN���|���	�|�Vyp�F�򩹨,��1��
T_���G��C֨j~���{j�vf��c�?����C�I��e����;�+o���Y��E��oH�|������Ɩ)�<��x�XYh
��G7V#ѱ
�R�@�q\׽E���~]�zM��!�].�+��+|��?�g�X��^
��v�n��fs$-A���=!Ix{ctnKA��I��M
�����Wm~���c��P^R�w?d��%���0�5��eD��?!�N{�:6oD�*�Ar���@*Ҍ���}�wc�\��} �W;��D�]yi��}�3e��=��`�^�Έ�B�v�&�E�׈�)�TN�u��9ckE�-���{���^���pU��>]� �6�U�y�/�m�?c�R^��3�D�����\�X�$9Cf�Y���[k�G�����M�@LЉ&���]��8�ԝ	�����pzY�M�ƍR4�v�"C%�J�;�����V|�u��&UQ ��/4G�I
/H����-[�\���W��P��[�ǻV=�</�Qܶ^h�
l�T��&�H�EL�U���׏�]sm�w��QM�T�����{Y]� HASQ�e/��5������j���u��T� �L���:~.�?W�V%�+�%��v�(ǒT���Z�ړTY7A�d:�ۙz�E�g�B��O!��	�1�f]��7��%��%���=.��?�~�b��D ��l����:oUUN�X|%a;�0P\�L~66f�g����B��|*��I}>2y�̜���r��T@ǘ�۹��n��ABH�\XRQ��á�.��;�̶	��,��n^��0�����Rm��A���ͻ��F����Cj���HiU�&~��jۡ2l2q��f�b7� 4aoO�V��Ȍ�?`�Up�������"��h܀HPՃ�/��%�l���ٝ��+u&�(��9��J:yT��1+����<����N�tQ{(5����Ǎ,p�E�o���D��}3K�ՖnZW҈ȶ9QN�W�j�EY�X�i�6-s\� �[�M���BaT"�nG'���ӭf�29mA�es��;-@��-̱�
��~�
T�x��,6T�E�8�@����(��;�55l��Y��5-���z�\��g��q�`�O��de�+�1W=�6�E,L���iB���3(�̜ii���Z��,��'��e���V�C����=��e ny�u�Q�=�֙:��t������8��<�}a���c�	kZ��u��2���54|,g�76L�5�v��F��:�|>�Ӟ?I�h0�LCx\�:l�=F/5[�<��7ZfBq6�2
b�G�^���ݳR�X��Pb��f�y���GJ��Fސ�)�Y̲�&�*�g�p����L̒�343��MEO��h(z�A`���J�8��|��Wbt�I�����k�k���<�@j"HZ}�})7�q��/e�޵y֛]~�_R\�n��T�G�� �|����E6��U@�E{��i�Kĥ�S���j{^y��4����'�Q�o��q��U��#�4�LS��֏�'ˀ� %eM���D�,G�Iy�e8eԑ��h��Tz;�6{��߅&[��O���er=)�yc��l<De�s�@gq�2�5�������mS���;��-�y��'��w��w���rf�b��z��>���s�߉�5�䒧�((�D�����qh����uط���2u�nF7en��c��~Fg�&c�UM��#Oqdr�63D�Oˈ����!T	�yIe'�r�P�W_�j�X@s�J�}mLE�n]�PH�@���z����k��W�Y~#��x�|0[6��X�O���ş�m��1Y�:�D^J�2�sύ�!X���{�YIܒ����l^�D���<��<^	%��x0��h�/T� �Y���t�ͭ������`�h6zWH$�����w�ϲ���Y&<��Λ���
Q���qB�)�����)�"1��ǀ��_�#`�XS ���j,��j����5c���s^NFr����?}�C�Fr�]E���tB�%���+��Ĉ�s�'K	ɪ�����M��O���v2X���=�]��/�Q�%��L�\ ��#²���k]�L�""��{?��}ΡȊѿR��'��������"�]�m�Ԉ�0f2Ol"Ai^	jۺ�~�c�m���=|�N2��� �����D�44+�DvZ�j���Sh;�� 	����|�� '�E�=�$�3V���4��~E��U�t#��4�C;S�:ZJf����x�"����v�{���m�,�����@܋X��d>}��Zr��ֻ��=����� �F�D�*��M�x�38\y���=��b�ҙ�]̤�Қ~�#�T~0oE�J�uanw��4ᛮ��B�k����P�Ώ�`W��׳Į)\����ԳKO�n��� ���B�;D̷�h+�qg���d����a��1�v��e����O�)t�W�<�{P)��!�� �6����'N��H�P$��M���Y�S^�F�T ���%��m�#8h9f��4&+���^��~wYRF�b^���?0�c��"I+�6d��h�|��<Jw/�n�Z�g0���7b�R�����v��L�n}��{��0��;Z��>��Ew.�z�ck9����v�� e2<,�	/���U�}����Q��d���HP��߫;_v������d�"6��2���r7��sD�v�I`ăYO�uZ�4�6�rF����@�-����3�14����o�$��K�,�&f�$h���P1�e�����X-�_Fz�{�D����|���e��l�\���5������:� Ӹ%���q`:)C��M�O�30��Sg:���!r�o�S@�Rm.��K���fK�퉏WU+��������˱c*tL�>�qO���:�2镛+������둍T���=�)�����'@-���X+%���y�-��`��Eo �JZ�y��.wL�Wld4����|��Gl�� T�����A�`�Pw�eޯ�VD!�sm��`͗��`]NyL~O�lm����[����>,���e���u��y_݊{�/��"r�7����J�=��aT�{�<��&�z���������*�S��ӷ\���k�c�/ǿ�ˆ��*�
Sɲ5n�N�\�*[�H��eR�z�n,+d�������0����"L�e�&�Oq�hk�b(�(>2�~�x��{N�PM
p�Z;�9889f�n)�*��ϭ^ye6U��2����ۑ��j(�.D8��-�_�}x�P��m=tԳ@5p|rH~Ӌ�٤�6z��1�l�μ,Y���V�� X5��)��2s��!y~��L�a;�ɗ�;�÷S�;D�;E|����K��T�ײ=7�@xAx�Y�>��
�0���y�p���?�f\kGj�k[�/fq#�e�5�ƉA\P.�B�7��/'#���d(֚��P1�	�4���@�� o��Z^��H+�.�����f���0��D�Zj�;d���?ݑ�*�j��Wr�ƯY|&����}�?u�n��l��],[�#��51Ո^-dmT�弞��!����4Ō�!ˈ�LMM�����a�2vV��#z�񘳲�������?vw���9����Pȱڥ|���L�� �)B��Z}��ܮ����Iмq�t�Gu��~��9�� M��FK;<!� ���o��mO{�0����wۥF+뷤����++R{S���1X�P^�x���OF��X����Em���>}�{�l!q,R��t���@�?��[����K�ϻMƒ{����6�Һ�����Z�Ԭ����o�増�|�ݢ�}�Ӆ� e����J&��7��l*�ZQ8��~�~��e����Q�n��)�(�ha����U!+�J
����i��_f0/��q{}%
��D�))�M��!���c�ȁ/p�{��,��w�"W����Ÿ͛�	�
s��_��OL�sS`��m9X�C�W��P�OH*?2�~�z@�9���-�bӺ�N3��#��Is��2&�b��\s��XEE@c"Y�Td>��[FlR��D����>F�1�X��kQz �4Է3��0�+����;��Q7�j)��)�Ems��غVC�q$�Y��\�5�OK������ �2��~�^�a���ܓ Y/��$8cCks��t�uZp`F
ג��[z��[+X��' �b7+��D�P�������ܢ�.>#%G(w(� ��c�7.��azچ�!PIތ���Bڭ���C��IdI�<蹗�]>ӏJ�ԟ�	�r9e6��;q>Ϟĕt��2��%!��Ū�T����m�n�_��#�"\)�yۘ�2�����ؐ��zX����©�;]���Y(fg2�Zh*(�h������d �j+�r���{�r\_�a�ҙc0;E��#��<i$A<�u�r�}�{Te��؇v2�~1�!"�a�9��_���D���37S&k�geK���:S݊��m��=�dQ��huq~jB�,�{�Տ�Is�y0B�֩ T���fN�\Nu�{G�O�THEy3R�V��L���Q���������J��;�e���Q�њE5�q �w��CU���Дcә*�%��Y�GI����N7f���K�mI�-m�8�@�&!����ϛ�n҆��ݎE�Έ}!�K<������*��r��L�%���y�xIZ�0�)H�@�.	�� ��1=���\�%ˬU\�/��W��;��'��]}�(�����;�;�T�n�{c��q�;A�TRq9_0��sǢ��������)1��﫻��[��'��|���I���^?���o��į�g���6��ޡi%�����F?P�oL��B�����W���: ���P�]�Tp���⋕��o꽼qN��o➂����m~����IL�ʺ�}��t��)1%f����-��MM�@��)�ķ]���U�����ͩY�υ��9�4+��Qr	�*f�&�f��M�uxdi4�(3S4`�x�D
0K;�l�yHڣf�9qoG�\�:.9?�& �1�Dxt5o�oDqW���=�1���Oki�(vZ{��h,���
�w	�f��٤�鿑o�,�x�����L�/p�,��E���� E�A� T���Q6��d� m2`�V�V�F��q��ʑ��O[Sj H��#%h�O���W���=�.ѪP�,��o���s�S����_*�p˭�{c�O���.|P��z�bx�L��^)Yh�'>򭓺a7�h B���@8[����ٝ xnmOZ��3d����!��bi���G�]�dgyX��_C�����dQ`��y}?_�J��b���	�gvwB�"qӟ�32aF
�p^��z^��hMj�fé��,��V����V�ҭQjۆ��д�9�R���S��6�Ч���m�Z1�\�W_Q��k�ݯ��55]Wy�F�Iwhb;��p����.��Gc�N��cmf%0Sb���V�szgPK(O����<*�_0>��Rb���:1{\�6�ӽ��1��~I��t9��������B�%2�A-����4��ø%f�#9�|��ߌ�dX��K98�=ڗ�8��CԀ�c�a LN^ 4,:���8�Fy�{��V�Tlc�W�בUs،���H��_�}����o��E���ˠ���Y�Q6�E@,�w�p��$f�A}*��yEÚ\�
A�"��� .ڼO��,
�=na}����~'�H&t<��Ik[{ԖU��� ЄP�o�U�M�G>�C����|߃���o^���/�R ��o_!���N6�� [*[�<�L�D�0:H�V�f��<�ǀ%Ǳ׵`��G�b�(��Ɯ�e�YE�آ��CO�(������m��$^/<r����t''�Vi<��I=��� ��c�û��3 &��W����G_L����w��ִ�(�t�.��ݭ1 Y��iS�8c˚�R��Q��H�_ �GZ���u�Rq�Ċ�5��HĄO����Հ2䥆�EJ�T7Zv�J�H,%-��g�_=Q$4y����hw����0��r2���/?+����X��`���R�"�:�����NG��*�m��#�4SvKP6,[�U~�^�Ͼ�a:�򻉗q`�~L�5�aw��o�ƴ`�{u,���@�?Uj_�Qǭ�����ۡ�]��[8�\n` 7��������u*�J��9n���u�e�}��׉O�rN�S .	��tz��ڹ��� 9	�	�0��O�){�T>r����v�=1�_N��w�� �-��&$��K/_/�5p����	ӚK���؄;�7�L@̶����t���ss�n����R��0���fv�d���+��]�J��V�jWkl��$��p�2����[`/?�-����v?z��Ж����~2�u8�@[��c��`ިp^�?���'�2%��J$)�fG ��:e􁽪�#L�͛�b�0��oo?����63>C�xq
���S��������T�tٯt(��*c}�2�WI�g<e�R�l��U���sw/�&�7p�k��or����8\<�m��F2� ��2/�=7b�}��&[8
*��ȽG:c����S�b�&v����w��I���j;��G�ŗn����
�ZyRr�Vd����qHċfUQ�M0>�%~w���OO8r�sl�ml�.�{}�T���?�����!|��V?v��b���6,��z�ɋ$�g�z�U�3�e�+�&Vl}!�l�<eN��8q�AO:c��C�2+��he���O�sf�۽�x	YXmM�������,���������+���3f�C��5CX�FY#J�Ls��/t~,���>������T}�Tm��4h���^�����wLS�<�V
U9HT��� �̚&m�E�<$�LG�4���Ea8�K�a��Ry�@����;y���βMbm��Cu�EWf6�u�V"#�|'�*�4�'���o�)H��T܉6C%����Ȭ>�&J�zd��x®Ws&t�C�kߖ$��VӨ7Tv\J��xn�wA�����_�DTy�%�e8�5}���dP��۰�a�o��Ļ��&��fh�9�b������޷7q`%��c�!'���r�7>0��+� ��O�����W4�L�����:T����x���j���$7Q�)N�W�����n6�	�l�g�-�V�}�?�_��8kڶM=��J��_�O����\�:}�q�$B�*��=��:jP�ʆ�>qj�*i]a�Zr��z/�aE�W��D2r�(W�Z���2�|;6��� ����e�Ҥp�0�����E��8��z��Gֻ�u>K�:N���}N$�����6��^YT��)q#���oM�e棿�]@��L��;Y֐E��
&#���&���d���S���1޷�nw�|�LؑgA+���s 蜂W1%J2V�`n�[��b��+T�"F�[Vn 6SO��&K�xr�#�H���va@8;�6����iTIw���<S+<�o�:*c�-萘Gx�m��&�� #����`ƫ��6
�>aO��-���cQ&6!ī�Qs������w]����)��y�,'�5�=��� F��L�]���_�iؔ!m��F� � �y �é�l��r�b_����$Y�t��$�o˩�5p��2ĺ�o�;��e�,x6��97�F,�@q��@����.e��.O�����L������	3��@J#S.��u6���먕)����e������
eA��s��z �RН�C�E&5ѿN)۾�*�ױ��kǼV["����	T&u�*y~Vu29v�|a@�)hP�����,ŀ���)	�%]����q���/W
Y
�3���i�*�ઈ7��ԕ#"z�3it��U���T����l��/�++�w�f�`(r��M|�ܕ�H�iS�o�2�C3��ǖ�sMj%z���>x�FF��Rf���қ�w�&��@k�U���@ze���i���p���H+r矞�B��U���i$pU;�tqp�ML�ErP���`��ije���0����{u%��l�Ĵ��t��éz!������ړ�Y�}q}�%j�gb���`I�,�
dR��� ��m�?x�!�?���^�|A������+���Po��A��U7ͽ��$`%���L=�]�P�`���J.͏��]ajfc��E�ud��f�5�7�;<�ϒ�#�|��,��ŬM��r340�$�� F��#�M�w�K񜲗5x��=�̝��嶖��3��M�B4�9��$����z�;@�>�=$.�H$
X�֭U��2=�"�|A&N?D0,�Q�71o��;C��;�Օ�U+Zy�����Gg�]�xѷ���<���ԜW��
�9�����*l'E�#3w$�?VD�'\���Rl؊L�V�v�l&+�YJ��DR�T6��9�V��^��Ԇ�
�b�u�6�O�q�E.����B_+�3���+�5���5ۂ ����eW�@ή``w^ּ�뜍���W�����)���2a�̦���Ġ��]��(5�Vc2�?4&f����=�?u�6�ɚ�v��0ѫ�(?��$sL�VU�@\����b���ٛ����C`���׌�6��V[���wb�5f�ת뛗���B�O��;��;�ю��^^�bu�, ����	��#WO�'D��E��F`�"��G��͏���WV�K�`����g��Y�*u�z�(S�o��}  _6�: ����W�k�S� �Soҳ��[�<x�P!l�)��R�����%6��d��Z�,n��6�T� �⁨���9���B2���ʨ��2��ϗ���-\a�B�ۧ��MK�&��):��������{h�r4Ƹk�$�8�tZJ��Cx���Bd�*��uP��m��2&"�F;@��0ֲ�[U+V����a�8���S5�:�
x�z���f����z����k��e��N�$w3o�5P~e�׃��!����q��㵊v�������Ao��$�~gC�B!�1)zY�O�����4F�)�UW���@3�4�Xc��;�� &ٍ����1`��d
�	ė\n��[�Y�h��t�]+:IL�>����B�d=��x`��"B��Y�ڞ`8vM6l�X\��QTTl	�U�g8-�R��6�r[f����G!�5U<����
���;�2���ٺ��6�Wtv�Of6��� b�X#�u�b ��X��T�b�&��aЬ�#S��n}��Q�����,p�)�Z�V7<��F,��ۧ�lJ��Z(��=��#A�h'oc��G�(��DB��5eBU6�
� ���e��k�*�;S:�(R���`^�%�7��<Vs�f�		�w���3��@H�`$��V=�I�v����_rH�H������@h���uJC�x�!��0O�k���-��?��uy��^C� �]�
��9#�*�tDM�/2WV�{�Ikْ����?�jb$�1�3��A�oMQ`�ƣi��lhF��'�)q����EI�mYY��Ou�$RY��y��9A��Ӫ�4�{54�֝>u'�$�3&Sv��ٴ�V'��?��ϪxKK��9n����}v ���I}�_�v&n���TŠY`�i.��;��1�u��2����TdR�S��ؚ�&	�3+dB�$�>���Gx����Vb"魿����Kws���0�m��j8������_H����6<��F���%b�C=��V�o�[��5E0�>��m )�����R'}v��>bY����@mK��e��Sŗ�U���]���.f�A1��h���>�H���ٚ����y({7�)K1�6&����ٸ��Bz�V6�Ư�}zqz�X7yF5���1#�J�[]:�>O�0�E�<W�'�ZgN]�'M�Ґ3�����N��%\'�J���A��*Q�G�#1�K����XA4e+�$��xӜE�׼�Q�R8 }8G�My��XƤ�h��9{��!u�`M�4�g�3,庋�:�����l�FV�lr�}/���49a���l����G:N�U��3'�2��2K��rA�s�
؋�p�{JEҊ�jo#0hy��A�Ԭ� K�UX8��?��]����{zpv�k�����Z�x�gpXW#���I<D�9��u}�΂��,���n�Wb���nk3;J^\��mat tF�B7M8Ļe&���sؓ�p�*�]��%3ǯ�"Ҕ\�MmC�kfa�3��
���}=��Ś�ǖ_8En�Dc�6�r3�jB���.D���$��$i3J�����{�mi5`�������ȧd�k�Dz1��C��yqh��X�
�Z���ԕ'�\%9����"�S����1q���\��r���f鍆�V�\���1��y�T�*�>k��(�3���Yΐ6�:_դ��u�7���"��Ә5C'=:�d��5J�r�q�� �j}v��"��������T�n�X���S�4��1z�#���\wecH}k�I�NK]�Vr��Y���e�/˧���>B��U��1����:�l���I�쯯*�(��;����'�g��}�t�L���Dd��NV�c�����Jړ�h������sY�Lb�8Jh۪��],L%ҙ�����K�g���ߡDN�Xخ3b�*�yxRCa�6�n"~��2�t��Ԣ�������b�2��WC�eaߥV����L�ȫ���ixNv�5�j#�8|"<�YA�t��Y򗎭�Ȉ��jxԞ!���h�*빣�7�� ^�t ���t�o�׶lC�$^卺���К����r�Ӑ���§����+ƿk�Π������fV���嬶�k2C��9���}���C�?f^V�y`F��ީ���<܃4�bx$Kø���
���H�n!?^��H*w4O�&�g��=j�
��MWՑ۳%�j\-,<�M��Sa��}�h��#e�B)D)C��l�7XPy_(I��a��&����5Uz���e��k��'��O�,N�����[ CH͌X���U���� [�C�����;�AE0LK�h#(���֐ϔ���#�����N��aN}=��ho���:WP�n�YE�]�����@$�u"�l�!T4S��6,kNI��X�M�Ÿ��g��i���3#�Ճ��&�yo��h �z8���[Hds6R��1'�K2�����>_�p����(oP�Pťк5���?�7=�+4�H����`+{��Z�@?ID��Ǐ��v�f�}�k7f"����pC0x7��(`3���]P��/���	Ȟau�����|��$�M�4��AxW���W�5���,����G$�e@�ŁL�v��NO���W���k˰���~���e��c����/����7��K>��$l�f�M��)y0S�������"�J�Lbw2anPT��O��6���Yq,�/�9cw<����,;�1��N.a���e�S�B�i��W�Kf�\v{����;�Z����C��~���5n���b��1�A�wp�s�+�yYW�M�Z�]ܭ��!�8<1k��W�ݛ��dV��a��B9�M��+��	�����I�2���	�?U��qG����Qjb^Y�Ё�2;fZn;L�./������0�i����yB�!��@=�x�^��F��	��.0��%�v���y*9m�F�	� ��p8u��4T��TX�H��E(8���W��O[q�����u ��P��#�.Φr}�_�:C	�A{Q�E����~1�w�����^Z��� �:�Krm��U�� �������kSM; `t6�`sF��LrĖd�f�*�L-mZ���딶�b��2xC[���G���751ĺ}�VY�����5�He�<��?��g�gS����:N��-	��p)s�.�L:$z�.00챩ѲƓ�I��*C9(핞�����\+� ���e�8O��zQ
���Ǡ��@���S�Һox���"W�!�,�>k�[�T]�����7�h"�j_�i8���q��FS[�����7S&���8����!1QZR��x�̇�F�*��f�O"�{S�EY��m���(�Mj�h�i90�۵bdb�u���=�<��A��u�J��׉7js솼�Q�{��R�W$�;%�j�5Z������Ҕb+�	�DH�ONo���q�h��fVq��#�@�Q��b	]x�y	#��8mю�i�}y�G�@��>��k�Ն3��K�"|Q�L�c�^b�l�XC4K�x6�`��6�1�N!C�qk�<UJ��=��J-��H�RE�h"��E�l�7Bp�(aEK��X���UUIWX����x��t#�wy�\���ھ\)�3H��=����)����,�$�I���$E
�y	\�.7�_h���9̵���%���7+]��~�6K�s�ǟ�*(k'�Ӿ���\�ظr�lq���1i��G� _� �ܽ�M�3E��8H��p(I��g�I�q;	�8�=���}0f�*�.A^���j�`1Xp�>�d�',i�0E9�ο���w��i����:י�t\#���V����S*�ߢ�˺�ꤤ��&Cs���]'�^g{A� �֘K��3@n�aZ�Eĭ�N6� nڬ;/��U1r�JZ:0�{r?�/S�F
��G�0���/�*���� х,q�-)��<v�fP��(�튈��������?!��6�w�k@����U[Q�=����[p<���4�2��B��y���`\��jT]
y2�	jx'�$z�,�t�rXd=D]�Zy^?3[6).�<%s}���Xl:���1J�;�,I� ��><	K�o��S�v�ѳĞ^��q��'T�y��՞<��;*��c�q��~�R����������X��(��,ѢΠ���$��
{�XXj��6�;x�n�����)�
 �Ի�,îʏ|߽�gWk�c((.�wVE�{�H2���1X���"Gt���rà�!'<5d>.�X�68l<��qEd֘�-���]cZ#�}���(�#ҏ���g�Qy�i�b2<x�G8fi����`�੧��^�j�|Sb��F<�������_N��JL钪
#e��fy�F4�#�����!���b��W��fE����r�#�r�o�)�ޕt���^"�
?��@���W��gyME�_Pb/�L CB5��|G��$A`��`e���g8��H��3�(]'{p2.w$'.��1[ Cj��&�ި"���8���w�'�ǌ;)$Y
|�\(zy�=��_�>�.kb�����RR�l'�*�c��T��I��J�_68��_�\��9u�X:�5��`�FU�Gmo��T<�X����a�>I#��TB�X�5��b�T�Oʬv��ep����| ���OC_��M$�c]?qu�X���645egkK��ѿ��ߦ����|�y8d���!
���P���q4��p���i����lq\�ۚ�[l��T&�{a��ċ��N��d�A)X�P��b�m6<E��d������F�N�����R�5��QQ�qט�Q]�KGmQ4��i�`3?��z2x��(�C����1	� Q PI�ef�lS:z��\�J.|GL�M�`b���S@q�z&#&dx!�Q~�M�\�D��Z�c糊Y˄ӣ����2���D�G_J�N-��� ��+�cf�T�2&������].�+4�:nsic�]��gO�R-ݭ]�,���,ץ"� �X�A�.k�h�*�o��E��o_����|&Ŏ��a�n|]�m��<���:e��֔��>Mzq���o���v�A������y�9ⳃ�ŭ�K�\>��m<I�Q�楓�������$Qv��w���&��:l�P�S�̰�HI�ތ��,���Σ��.�'�Zry�p� ?��E�U�ʌt�-��rV��zP���G�ܾ���G�Ӧ��_���F|�:�V��S9�/�<�́j�^�77z$ƴ<Fk����A��F
τ�G�4��g��l@���h�+��4*��Xz��,ǰW�%�!�o ���O�x���3�?/Eg^T c��R�ˁm� ���d��68�vH�M��6�W�ҷvt�ɓ���l7�"��/���Q=��N��8����YFb@�)&N��.��M���4��>Xp��U�bH�j���N�5�����8�OX����M���I�w�mF�dϮv� k��|�:D̀�ی�����b��;ҤO�=Z���J�� ,6&>o��&�
!s�>#
W$:b��91{G����r�����7cK�.YT��4q�+;�� z�KN�t;���f�5�M����Tl?�5�J����w��d/+�-��>���S �+�$;Q�Δ6}�pG��nը�Ab���gmzl��Ě�!�H��t6t����,ά�Jb�q4���G�E�����v%-@t������x$Ŧ��{3R���]�|ɋ[� ��a4~�uj�7y}y�z\׭����1��=�ݎ�2�l6���5lo}})��VV�j���H��@��iQ�ҕ$�m��?9��%����ws�;�G0�T��}[�ZF .�3M�Pƞ��.��	�C��5�[w��m�Q<���@��^���AM_"odT��;F�Bhx�\n��|Ҏ3,(�������4����2�}(�0���5�(̛���Jp�B�VF�c�3\*���	�.���V�ک�%���*\�G�$+`X���)�~�����Ge�bg��ջQ��Iq]qІ��Э�#v���^fX���i���N��*y@5���R8<9�E�4�O�{D��n�;3y�W4;�߷@�˔ᝩ+��Ȩq��̸�+����.��>��i�.�vx��ikqH��}!x�Dҍ���U���	����g�����T��n�2�!�p�ܧ��A| ����ʪ�6�晦�`�EI��g�vRL'��﫿h}$"�ʚ�~��V�+��}��hq[@�h@v�#@H�m<.�T��܇|&cP���)���Ƌ]"앸�&^$�B4��m;�Y�\��\�Nl~�V�*��'����Į"\:
� � ?Ӛ�f�i�n�oKVHU�n
�q�g�m�#���@J5a�5�׾�-9p�� +��BjN��e]�O�r�mm�.t��� kh�Y9r� X*���H�̰�%���T��sM!?�5ҭ�c��N�9�V��9�9F/Ti�,��ʕ/8]����ݺc���BsB��G,>�L�;\�[o�iEt��`��;�w)@
��n���T,!�I�N�������T�`/[�$�.T�-$�TTOIf�B�t�[��&��t����ck��!z�*���f�.�����/�<��f�M������[�����x�F�~�$ 3k� -]@�����rC%zp�O��Υ�}X�	��m�9i������V��aT_-K���ko�9��	Ms��q|}��[Jʨ�<�e=l��ޜ�{�l�]�A�7Lz�̀U-�N���@��M�:���@/9$��>瓏[��>��E�$v_#��Ρc�A�c2Ń����S�?%����g5[��3�,���+Ђ+C�3?��1�����Y�l-I:���G�8�k�0�~!*t)�G)����%vw���ԕ�Dr}�7
Ԅr�$F�E�E=�Ή,���U�D��s�ɸ�)�/{3��� +�p �͹I�%E�����/�i�kI����1�i��a���:�Q$�����F��=h-}u�%`��U������UR���~h�*v�� Sa
��}k�Sp��9� aM�!Nee�㪾������e����2�<�����骰�c�(��A�9�FA׹��]�f"�;hu yG�c�q��{�P��c&H2�d-ܡ,dy-<"��������w��~Z��B'!����F%ʄ��Ua�(rQD�Aq�.:���
Rt��A�t+i	�H�E�q$��Ωq-}�;��-��t�ɚ��B�c���>&K9����g4�V�(�[!�XG�����1%���7��FU7�1��.���h[���J7(B~�f`q3��4W�`�"(Y�U�>�<�^�]�tzy[�XVE�)(*M��NR�;����*B��cu�7-��Cl1�ہq1��U!��D׃
��8��j�BEl<]���S@Eo�:cR�+Nm�k�P/f���q^�L��C�~_���tv¾�mk
��R`[��QծZ��C�	��]�+�����TG��E�#3��!��A�E�E��jFw�v8�i�w�=<�~�>q;�L��[�gudcVh��ߢ|K�
�����V���|[(�}��{�� &z}^��������bw�5��7.��c���^��_c�$~i�2VBG�4D<����(�}���Ӝ�w =�����<�n"�QN�̤����t�{D�>���A�\9�@gI�N��AWM�i&�����MޟӋ�J�&%�1V�,��rD&(vE�r�c����Yf`��>Čx��w!N���	��I�0@�Y����RZ��5�����*)��&�I/~G�H��1[f��+"+ZJ�Ő��q�і[�W�2@��1��l�� Q\����nΥ�r5�HW��p�f�R�J�Ur��z@1��fi��d_������Z���u�d�����H����kaZA�̘[�w�,@�QN�4�O� �#�G7J�d����i�{U��D!������{��2$W@7�h�fD
�H�x���&�_�1�z�!S�1~X)s�ae����������\p)=UL���U4��B��w;Vk�i�m�Fy��j��P�� 4��9����tM��?ϧ���4�-���� ޭ��h�JYZ��yg|��eex�1�u��д}�|��E��e�*9��1�R2��'�'�A��Mn��$�H�?�˄�k��@� 'էh@�y'pa�����.�y��C�j�֪�\c�%h�����X��2��Wm��dY+-�3� W�"r_֜+��a� j���<�:���9bR!�ߤ�~��H�Qq��r�0�i�xϫH�9n����v�dКk#��>�.I~l�p��m��p1�k.��F)���$�������}�