��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��s������\�Ἡl-�y�f�����f� �ѕ:�nA�kb-q��_���ѹ(4�dê*���7��N2�ɐ��+ٞ�4Y6Mx�ejǴ�y9�����=���D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6��\\�l�����r9s��@'�k~�{�<���y�#���i6`#Ɉh:^[����*`��Z��|���z���N?`q_���ר�Z���FLe���Et *�mkd��^�\D�{�Ѫ����+*����+�Z����� ��ԓ*n��an�7�?��!\�ݠͿ�L=,���a���Nk��_=���}�7�C�#T��<T���w�w��ƕ�_�m�����դ��*���	�4+��Ch�S� �-�6�똒��Om��9ד�0�XZ\,��zF?|���﬌62����&��)��*�GXW�f�72�!%��F�c�R[���f�s#U��"� ��b��*>zT�9D�'���l*j<�$Hm~��ˣV�=	ʥ�>�/%��¸"x2�hW��t��mK�M��-W��f��8������f��U"p['���]��Q����ќ���W#�U�5�5�S�
P��܁NNɅǶ�9���#�S�V���1U걒'zl�c���+���os�S���Er�����\:�'B7t&���ǌ�u��Fz�A>�J�rL��p�F�	*�s�C_�BM�僐b�Ĳ7x��P���QEd��d�Z���ou낕Z�i(��[keY�^��1}�".�������'5��+Ï�,�.�*It6�-��{�⵿��8?�C�FZ�fh+���oj������6����W���>��ك�L�"0�M[<���<��g��?/+��o �E�>��XY�ד�N框/k�y��((�N/%�o_�,��!���D1Č�����f�p�䔺�
���`#p��$�P)ש$�˿`��?k{u��/DP��_��X���0�&-qDǱ�(i_S9(M9��>dU+��&_gY�6������$H�)55��QK\�LD�$���cl����b}2�v@*��+r�����`�<�yz�����n!�9���;潠V�}v��7]3'�g�W��8�}��0�9,,$�$���s8L"r��qYj�sU�S�D^؀��d�;Kp���kUW��e�w3��b�q�o�h(��1���r�HP%1�%P�y �)�7.2��Yw|m�-+�(x�7/����"́�I��4�����}�>��k��15lu�&�1�,ͯ�-�OA�=]��"I��D��JK6pQ}��Ϟ���8��;�#�-��?���?]�����*�����L M&"�_���W��)c�����}~���!�eJ)=kN�����I�t�8Op�+>H��88ɂu(�����T�w�h+9Ah_�Cpm�M��˯�<� +�z��Y)hdNq�~�ΦO�j�z&9�C�`��+�0*����M�X-�������)+�� �@��M�$�CJ����OwIw4e$�3���o�#7ա5R��g�һG��C5�Tu��AIBޫ���;�4T����9Ӳ�
{��H�ڨ�;�>Q��A�Ҥ/D@"�����*�\Uɪ�|�<$��
y`��o��ִ ��w�
�����X4|U�
�^�p2�>n�6. Q'j���_7��ÑQ���=TC�·�zI�5\C�R@��b�N�h�������P)��$]$��TL*+E�]g
S�q�K6{2#\`5�ݷ�����̘]�9��L ����q�W�v�����_<$oo�"���H��/6Ѱ-/��O�u�0C`��M�ƅQ^���F�		�۳�t�*��\M���T�SA^I �T?ό�Y��"�z,�
t%��t�>�{��,�Ws9c�}�؀��Pj~����K��ⵯH��"��v9!Ek�A�$9�4���w�2A4��:o
�4P�Ōp}�{ID�)&ڶ�x�DX}Fտ`u�k��p�V�z�""��7��k��>q���PF$M��|S��lI�?jb�)O�Τ�A��j����Y��~�y2Q�+������.�(��n���U(���K~����c@� a��vYq'�Z�����`B��K���T�%o/�M��2w�f�IX9�\�ڎ�1��V�
g@�ɵ�E!�����Om�]�E����^������f�~d�ͲA/�\�����X<�RDus��(:���DQ���-��_���' �/A� �K�y]����ߝ-E�[��ٍ��L���7�MYuk6;�+G���tT��G�?�O�K��rY��yk�^106M�B�m��e�ǜ�.�Ȩ�·�_;KW7'���k���}.�Lv�Y���W�����E��S����Ї��/�̳�&3l�b�Z�lx=y���LԿ�Np�2	sr��:�C�)��)��qA����W�@��.ٺ�����G�	�цX`6l���"q�G��5���`m1U�}�����Yc�j!<�q�ck�D�x�����Jj�ᴥ��	�b�o�@����:ڟ;�M�I�c��hsy������  `F��@yd��:F��Nf2�?j#RP3�HYg�GR�k [A���P�^IN쭤��9�+(t*���H�����Or��LG��^��|�QiR?�<�iE��d�F�U�F ��W���zZD5SL�4�o���"� yXE��G�ye[�[�V��THy�k̲���N�[�I��!tt3�P,Zok!�g�"B!kn(q͔|2�B�*��M�������	M�4���!]uR�_>�-���6����@?��� ��2���z���A���Ȑ��.��N�.��u�/������F.�����K��q�.�Ԗ��K���LX*	=�
8��x�AB���p��L���;RA*@گQ�]�,�牭�N�]C0��=����6��]����v�}�Կ�]����)+uz=u� ���
-��#�,*s�y���e�pO|���|0^��<��m�X��B(�R�� �Te�K�45j�������6ea��T�v�h�p��sI��r+d���E�ǣ�lk@2*� �rF�7Y�g$�X�jI(?6��U��e-ǚ(9�K `l�;Es�9V����&ՐM�$&zk$�a�=�s�fW���J���$�%��p	�0=���-��`?|��3�}�;ok&��B#���<�-8��?_B#�JV���c��j<N�n��������C��J&��Yyuot�"�?�}nVe��jq�-��p�2y�\��i��|z[�U�˒jC�w��ܞ���ex���`=:����-��#�tHܭ,=�y����l\�1$a��{�/�AD-"H� ��Ψ����iܠ+��L�EE�1n��C�E�#������hq���Z|�2s�"�����R#�G�֘�C+�o:�B =+����$�� u	�
� B���`K����1V7��Ն�ݵF��������2��#����� :�7ر����C�#�|#�s!����(到�~�^��0ƞ�0�h4u������0�]����˩~W#��B(;��ג��$]�j!�"!q�TC��Af�-w��="FG�(�~�LSQ.7xs@\��:��$����w@�w�"�u��%�r(.㽡�ެoC̡]�,%���UUef!P�y�3m�,��1�u#�!��DˠI�D*䉖+�%<���"a�YH��R��4C��l�8�s���Q?�*�2Wſ�mWFQz��;-��uC?��%Ҁ�Q$-�uo�A�Ê�y����K�w�:�����D�'�]�p�B{��"j�iEE������Pj�a/ʘ����h\?E �"�RD�UQ?�-�Х�6,�4!oጰW�WW�}F�e@ �_V�}p��<�I�����c���R"��j:!��%z�7��l(�n�a+ߊ߫م?�F���(��݆?��)]uzVl-2R��a�n�B"L-���,CF�`]t�2 YY�1��_R�mE�+��IuJ؆}�ɻ��?T��Gw���c�?p5k���1�ה��XV��F sH�)���4�߇%Z���Ѣ��7�Cmw,S���r˛��s�R��*�7���^��ڨv�/�yW�^{cY�����%[ۂ���D�Y�������x�c����h���[����0�H�2�uFx'ؖ���UL�c�&x�lJ.� �<Jfy�s�d���S��$x���o�F�'�>ZO\ij�hs��[_~/K��g��lÖ�0f���v��N���o�:P��ĩӢ��>\�[�~#1¹��O�}H����tg,"���2|,w'�i�D���!�����AU���s&X�#�ky&����մ�fn"�I#�}+#h��$�̘��qz@�A�%�gTnX�𷄙���[?�g�wխ�{�Bȶ#M��
z
�B1΋ұn$��S�����LJI�,JˤY`�G_�ur�<�e�����}��	U����9��C����f�̆ud����)���W��L�s���UC����a�D"�K�X/��o��Z���!pml�)0��r�D���x�r��g�
�Q�i��((���C��h�EP��"v�WQ���wHp��?�u��n�@��u8+Mp�B�
ӥ
u�����~ �uP}�K}}�;�e��/�]��c��=�(�#�t$=Qr�S��R�G�ʣ��%PtR#bP����.�o�̙��V!әѰ��8��En��t4W"�~�Ղ��}}ܙ�A�0�g#���%3�ZZ�fz���t,C�ޖ ̯����X�$z���G�b�-I����q�����ǌ�F�|�<9y`�RSAp�E�����ǫ�]J�n^��Zs���
)Q����H�Q��F�2�h(��� s�p�u��$2oڤ��煮�v��B:CX�u%JAe�;�@�3�����1x��Q�����^�ա�/�����������.�_��Z�a���j0ۨ`�[�;��nZ��S&�	�����IO���7N���y�w!�9ꂥ�0u;Uϡ�,pj������Ő��G`�F�,B,ToW�4�?��0ض����U��S�sE��{|x^H����墩��� DmcK^v���"u��|d���wt&J����̫�cS���F�����y*�)�b�(�hǘą�M��lxI]�Wu~(lP�}мU�W��䯎�� ;׼�nj: �L��7t�Y,�-��d~M1��;ej��8 Yt��
q���Fg�Gԧ7����v�ps����p�(TfbC�Ƃ�~����/9؅(�� T��u�&5f��Z����욳J !PN	�K0���O2@�@�\��hP_������D;BMa��j6�����?!�,�oW�\�V{1��x�cjbv03�ƒ�,��
c����o�$�~�?&d�������_���桧����-�V�e_��ޝ��y�'4R��E����V����Lt��W�k�#�&������ժ���eI�t�SL��7tԬ�džˇ��Ţ�N3��Wp
_Z�M�
7{�^QTj��m@�y��
c�]W���!��Ʀ��ҭ�����}sȡDp��j�	H��=����X26�����L5�QyX	�Wo����r�w�����ߠ�7��6�O3?f>�yc�٬��l�����<�ޭ���
�I�MC���H��t'�Pro�Z���������r���8��^'�����^՘�p{���*��1SZb���P>��wJ����T�V���	�����E!�7�%��	ݯ�D�D�Y�[���E�/�y����V�&������%��
�p�4o�rã�O֗��ֲ�3r�-�v<v��8$���y��g)G9��
�U݉	��
�%Đ�l��9����A���EF��i��b�Vt<3���]��+�Mٓ�����\쑢Fz�M�e�>�O+�Ϟ.}�)C������̇�?N!�cd!�Jm���2�J���&��4�F$F��1���H�a����ON���j��i6�hP75(wt�7��=��-��
S(H,�"�~�d�Ӓ�,i�p�V��V��:2C��]񎴆�Mx��s�i���ysW�M`�g��(��irך�	40M���}G^���Q�u��ެ�Y�4���i���S����S��T��?kN�������X��AV�����Jb�Ϟ3΃�B_ew�����H%S�ww�t�hm��u�N��ؑ��/L����J{KĪCȇ�8��
��6�"�� E��Gx��|>�U��T,��G��1�+�y��ZwƗ�=��@��wQs�(��V�p*��3ɫn���d�W���A�s<���Ĺk�5�R"��N���^œc�����>M3q��M��uu�m�Rm�T7��i��+��s'�^h�ʻ1�O˭OI?���~Ch���lu���*���IOr��j�)�؋�sx'q9V׭9!b �j�y�IE&���W>��(psL 9���b=/�m�
Xyʔ�6��ؽ-9i�w�޺;�gc}T=q���V�9��k�Q���b�A�)�`�w[/�i�ە�XP��}�"zh1�R�L���7i���Z#������E�]Y�S���\�'lp^�zJ����9z▨n`W#�R6 ;Q�yO!�3��ze�
7��?��}$ݳQ�� tZP�aʆ�R�}������oPٖ.���_���C��n�F����M�{��=����s O��o'�����k�����aC.�#3�4�]7����t5�b)�{roped���=��/���Vc� ��={,�p��7Z��~/��&[?��,N�p�RF�����g��W.�U��WVԘ�^l� /���	�yo@<�&�@��O��F��˩υ������`e7�?���$=�
n���\��p�
��l��#N�_+j�rELt�6tN*-�!$s��ܔk�tbb��+�-���B�����	�T��E��H��]�r���̑/�K�Ǉ�������f��+$t�����f��Y�)q4��� ��R��
$�h��Ե�IWM�0���ޓ���X��/��5w�!�I��\Q�-��y��k����;�i=�9[�\).I�(2�s�m|���qSGV�Yd��sbږ���o-R��RQ�BE���

_� �V�d�U�R���{�J%�������Sl�( �B�у����1b%]�_:v{v��KF=䞞����.@�Ai��r��D�����ٗ�ׂ��2H�ǿu�3 ~1������N�2[���֍&=4����x���>�%όJ�iO���+���"��EM���'L��0?��
���$�(���������#\lY��� ���8U}$xj� �GL�a��Z��U���Z�-��f|�uz�M�F���DjR�k��J��[�u�1���k��M@f����s(���L��������GJ��:�x2O�ܟ�4�r�|��V����:�W�{�d1�ë}-*h�ӭ��E���Y�ƃ�)��.��cjN�8��h�H܏H��D�b;��;y�t��@�8mgϱ�qY6�:�+Ү��1��Yo��M�?�N�o���b��@5�Pd��I����<R��T�|����A���&���K���G��le'�o(q4�5+������qW��%d�]^<�g�]�tG݄��C���f�f�b�TaC�o�^��{F�ˮ�����l�;s����Z7֑Ӻq�lR>�����G_�Zx�[cy)�}�t����)Wl��HrG���:��W	h���������7[�U�oĬ=RP�hU���y�4�h�;I���u3��8�3��;��i�6�K�^e���F��]E�Q��p[�����3#�����-_�x�a�y��i0u[kK�t�[L�z&�B5�����-�,�[IV>N�I���1�X���.N^��H�o��`6M��E �	m�Nn�M������h��k�ۻ���x��5ᗑV�	룠-�҅�j�qHl%�'�^a���L%��9�yˣ��*λ��.�xOw���qC��h�A.��"^��v��e�
4Qtf����0�3���%���0B�3�_*zs(Z�t��}��c��y��
�ז�dP# �����F�B�!?i�r�Eu�����J����0�^񎾢_V $/l���ƍ� ��s)�63̠����,P�E�����gv�݈?7õ$}��[S��}0��8Z_z�@����Goq���e:1�fQ*Y���'ۋ�vIN~(����mnU�7`4�*^�6�$N:��83��r��(5Z�2�o��D�2y�|�v��_V;�����V��!�)���ۅnK'EIN=�Q�Q�ЁG2�hZ��S�dw$����*0e���_?Ь_2����M�	אy����һG֮�vK�r;���*��ַV¿�m#T�h�f���ҙ�hX�&:���n�Dj*��L���c��
dzq����j2�/��\���e��PM��5CA�"�!��J�M�:����Z!=-]�_9`��T�瑭�����r�������\�aB��j�E�#Ε�:�N=s/H\-)@2�q��d�ϭ�IwW��qdG\3�	�b~�x�30�rf���z_���i�I|�``�{���aQmPs���Sa��Bp�c��d�{{9R"Ȋ.�_����qm���N<q��,�in�:���	]+�+O��`S��ɸ�9c�4�m�k;.�Rx^Y%G���&e�r
�J9���F	9�H�kp����"O���O#������ު����a:񾟊$GAC$I�*�:F�'@�6� <�q"�C�|ٵo4/��{�<��<�����|��/���>�c{N*�	�C@~"S# ��<���./�{u�� vZ��!(�����Q/��ݘ��Fk:2ұ��d�s2��%��4p��#|�w�P?OZ>I���u��Z�
�)Z��j�_Z�^b#ØU�c���}xH�E�Z�_�����++��d9*��KR>�� ao�� ��%@�&IT�Z]ȿ����bQ�E_��d
	6�>�w/N�=|շӋC8ku|<7�,���=�'�GC�N٦.`!�tɯ�<��r>�r���=����N�+h��^�^�٢\��փ���b8�"�2u�B���_r���^B��f�0$�9e�����T�d�<�h�E��X:/��vi�
�q����hhk
�4-L�{��`�bl��y����(�׼�^�/I����'*y:��y����'0ۗ1�#����;(�;[R�3�}��*7��3; 62�.!��ww�CY>Θ#.��LWϽ"_3�:/M�����.M�Ө́Ah����8���s?��1�r�Ԍ"�G����{	'�ae���X֩x�BU���R�E��G��7��i/��)'9�����7�v��T�����J�H��b�t<e�Ͳ����1,�^^�4d��Q��I���� �H��i��xګ�82FwZ>��{��	
p'���nL;iA��8��QZi-ٗ������%�=�.���Ҩ1-7zm�>3��j�w\6��y�&���h�$t�Al�1����Ų���uA�)�OW���ZD������4��8�(�!���wk���-x��k��Ꭼ��kZn`�"~yI��`�:�lIy	��)=�8��{���gq�"�K��lP�쏀q/I��h<��uk���w;;Qm?
cb�
�,���#�A5l'���4��T���B��H��R�]E��/XT�-�^؊`y�y���hQ�cC�%5���)�8��E^;vYi��i�24���U@}i��g���".�kh�A����vS��E(���<"эB�� �h��V!I�f�}I�%�fu��Î!���*/�_�/س�\�Gx�ITs�N|b x�#p�������ﴈXR)e�F���@97�o�0 ���k�#*���2Y��G�U��!�����Mr��?��2�vו{�������Gݢ$4����S$�x�p|���
P1ɜŞ�`J�N��˥?wBH$�dn�2��6f��{�ɽ@�%�[���~L�O��p��/�(���;\�9|�5����S
=�]5��t��L��9��1��?'��
���!��+��5�%Dfe.�<��ϖ�N?��y5�FDuAUE*��;�R��2Z�T��8�X�z��������ӏ�(2.|RP�[5�Yo��4�4\�)�N�1�_�?mߦ�p��0����,�	���j_a�<��7.������g*��#2���U����իV�C���d9x����H�+'��{/��"M�ZR f?@\R�t�_�<�J�B@��l�����9;��	���-L)�2�H�QE��i��������<�k��
$���'�����NI�⦼��z=G��;�V��[����$l���>�yc-�L��������Í�+���gLO����,�{�o�;w��.��"�/<E�_?�~-��qa�[%z��@Z��Ҳի��8�ov�D*bAϠ_�;�Q�T���[-����zu��>{`�\��OVkHiD�V����?�dD�-�*8.�W���f����!�ݔJJ��<�-�5���}𵡢��9�ZR> ��o�Rg��^q��6/�@�r��`��qޢ��D�Ě�[�,g*�x>2�W�ņ�G<��½�}��xU��G��y:�::��T��vc{�I��N�O�l}���5
;��&���^����{�F%�����M�=��k\ zmQv9�+}�9��v�L�4'�VR���Ke���s��`����L��[�y���UL����b���f*�B��蠺�;7����Y,�-H��A8}#�ѱUߖyBX�sDw�Ym�s�[8F��z��P�l���'<�fq�c��g�
/���S3��F��~$��͎�<��}
�fi�G@��\a��F\���P�Eiu�q�˚3��*L��<� ��};}�oC�(��$��%�`,w=Ϧ�՛��� h�9%�@9ľH�E�b�WH��j)O!�G�SW�Z����	�Mf,Q����r��Y���x�h����&�oKp���|�"�WE�``p��Rz�y�,�ƞ*ȭ�uc�ZNi�vXxj�y�9�̽,ݐ���?�z�+B�B���j�D*���t�h����:�Z��Ќ�䝽 ���A�E`F(���A;Y��ڃ��P �!�p�p���d.�]�yO��!7��1�H�w ��={�<��6���p�XT�eV �{�ff�0�P}5��=�H:δ֔�2�:��f��ؼ�U)ݨ_� �'O��_����4�����	s��FN�U%�W䓞B�>��H�7����XJ'��N6|���MB�?Fp�_G%�J"Oj`x��5$@�ܧzf �������h��,����3係Gq�׶d�+(�7x���@h��|Jq����dA����
�k*���.g?����q5씨�\��E���us[D�CY�m^�gy�
*���@JB��(k(ӪFm��.	 4س�-��G�f��߆����j��F'��i��[8�T��P|�"}ס�'���I:��#��)y5S�I��F��0�ds��(�ٽ�ԹL���)��� �J�_I���m5g!2KCF���\�������W��A󯭜zJ�j�C���\"��[~�ϑJw���U��ه5��>���B�B�z�pѭ��&�,p����4>��q�t$"�o�M(K�j&$��)���p4чZ�Y̙�A��Oh2W^�0u���ٻ���p�Aڥ�Z*N�riG
��e��\�Z�����Dnl�G�YD�qN��7|ɷ�r\1�S�eܚW���w+|�L~���+	�h��)�x�B0�)P���#Vj�ŉ橰!/�O��ؤ��Fx��b��Eι|N���1��-�8m(&ݥ�E�&$��Λ9���jB���FT�1	ԣL���F�~v��	��O-�/*�?�|�v���>1"�nP�c�x�eq�غ��* ��RV��~x���|2��8�T��K���g�+>��c��ȷ�=�G�$d��fu��G`�Q�'�d��������ԅa����_<�~�zn��@�:�8�K ��a�D̡�N()���dw��ګ�9G��Ĝ�"����C�pX��s^��v��9����	���D�v��L�QJ����6
�_��$9��ܸ��j�ʜ���u/��e��'{u�P�x�����Pf�9����p�e,>�k��ni�F�Û��[G�&H8��Ҁ�%�q^��F���3@4J����W5��K/:KM,��,3��/%�$YZ��
���}sbC������^�)o�4.�b�zkx�Y>��s���BZ���Aݚ��wJ̸&UJҼ|��B����{8A!�������R��06��h����A�����e��e\�r�3��ȑo@���NCEF,�Y����UHl��Q`$�"�8�����u��XO�m���%��:��=��r��}�̨�����W#E'9Ya�W�ԑ�'7�ң4�'D�_C��h���bx���>1���/�Dbw�o�B�]��^&�N��!�zy�wf�<i-֍"���r��7��Y\E.�_�`,P]������� gl��G<2=�-w��b��nmG��~A��NX�ɛ�w�C���z�2���f�#�#�@���?�n��/=|e �=�>�@[�\���=L<���r�?J�Y��.|����#	�6ѫ��/������]����Ħқ�~�,9�k�[�<��ԸuH��:h��8��=�4��g�;�OQ�;㯇��@򬉤b��Ʈu�ꕥ;aq�3�	jvnV+��W�� Io�^*����C�^j�nf�̃k�zǂ����yy��(�@h��z�'�%w\i7�T�uu�����Y�~�j�
�EmH�K|e�"��&�f��Ót�w��X:�$A���)��&����"fd�U��AÊאV���+(��_	�`~L$�8Фp�� ��~3]�jHM� Apa��H�nFt�����|��xe ʣz���(N~pp�E��,<!)A�V��Z�b���5؍Y���HPل�`z�B^���l��q�=��������q��n����%<MT��R���X�=���ϡo�L��l�	%(��N2 \9M�zR���}u��޵bsN�d2�4��S��>[��B��2��v@�؏�g
-�d��K3��,N��]?�����̾�� ���Mگ�FdX��\H���|�b��9TP��FN�D���J�}ʞ}{g��i�Wf+Tѓ�? �O����T۹�����U%���T����+p�v����΂�v��Keԅ��r1kXB7��x�j�7Yݱ�g�ֽ\���S¾ݒ#A>+F+�ޢ%F*@�n%{C8��$>�A5��`ҾN
�f6��]�n_���+z�KR�<j�n�Hm���	յ����˿�T�� ��F!�R�7�x���@�khl&'\�#���%����;��p�tX���<_Q2����U
r�X>���F��F5��ήD�5�ҙZci���%s'5I�����ն�5�_-�4�e����%���?��0)d.3���ں5����g����pS��{H��h����x@�r����;<�F�;�b�ds+*$�����'=��b�RIx�q���{6Y��8�iǞ%�V���1o��s�Z��樬<�j!���T�f�$���tU����_E�x!���-4?�R*�R�]�9�%���������@�Cy �W�Ԑ���R �T3d�2�H��^�(Rʴ�>��ⓕa����UZA�8���3sIe����*�ifM�4ßp*�+�T��u�5��s�g�mm��}v��!�z�p|�y�Jax,�%�M��G��xzUL(?R��T&���Wȅ�K�MM��R#�UyY�Z(����յG�߾ޮ"�0�+D�����	�˗�[ߕ[dd��ܪ�$Jt?����Y`���Q#���:}T�$��1�|��D�!O�{�p��TFO`p<4����f��U�S7�	�|�F ��l1ZH�m��~#/�B��/F�q�\{'($R�60�K�G�+�U���"���ʇu� �tV���	�e�yIk�d��L$g�C��s��a���nY�Â^9���ӏ��p�XZN�L�mE����Z��w����"�K�߭
vw��OF����j �L^b��n���#�>Ky+n����H�q���\2�2ܘ.kd?k�=�h��p����Bv�q�N��ّ0m>�DlU�v��4��F��4��f� ?#�{͌#�W���;9�:$��j���0�0ϊ�?-�D�w\��Z
+��bTG�����\��ǎUc��z�ߒ�#�v��X��\*��b\�p��ځ&L�`���'�W5��]f�i+&�}���B��L[c�0=��B�9��Tz)��ۉ��k�ܴC@OT�9�}�������on!�\����7t�����p��n0u�c"�l4';�c9�^5Vf�b[#(^P�ѧ/��Y�-yme�9g�1Ȍ�/ke���Ca;�0��`��`�BB֕��X�6���L�
�M�}�,������fd)�ٱN�7�S�ŉ�2��H4���-�%��'�,��j/��]`��;�$�V�����Y^e=�i �x�s�1*��T�Z^�rZ�r��봑�������E��a�i.�ϭ�ME���kx�އ���2IAJ����t���Uc���۹�U^��i	�x=�z�$�^��n�rZ�<���Zk��ǂI�K<ƻp>�Na,�����0h~���ց�(�=�(�;��1�S��I��]�@����ovM 2
�� �����d��o�Oxnv�|<�Xk;Y�*a�g� ��\I�b�j�\R�-�n]�I��K����o�����g}ޱ:�ֱ	D_���>�%3'SaE:�m63(產G��1�e���T ?�:�N7�[� p$«*ځ���l3 ��:�_��p!�g�Å<%��p��y�̫	��	v
rOV: �So�0K��e�]�-�,"G-�+�������ƘqQ>+��e�GN65R�\!C�u��P"c�&��21Uϙ��Y�O]B�"ޡ��R�0��������('�(@�`1��^�s�:H⠆\oJ����s�JP�KGxf�2�bY�=��?'����	��Z�S�v�`���tKVP�k�#ʄi��~�!��>|B˼�:M��������zaw��W%ɒϴ( ��옃B��Uϡ�l�) ��1��T�_��}2���=�ln^"7�f6��t��\����+X�y��@-�I�a�T��F1�WO�����R�W�n�|�t=k��v�����u����a��`|��D�T-�a(���s�[785���P�����U��dڢ# �LD���/ޫ�çM����_���%�=4��/A~(��xn�3�����zoV�|it�����k/�� �T�����R�Ӂh���-'��<��ぶil����.<�h1�Z̙��c�m��{���`!x
$��YZlN�"��dh� �*3��t�]Ҡ{�g�F�M��9���iZX����Z.p�ߘ%H�fS����jı�"���&�CJ�o�o�O�"粉�!�E_����d����`L$+�ނ��2!��$қ�|��%���[�����x֍�{ZN~>	{C�9����Z�����23���76b�e:�8�+U�G�kaOi�1�ZßtXx3a����'�!�B�dd�ʜ��LU��Vo ��j?�ݶ$4�W^�����j0�	��'��n�V�9�.�T֖����K�{��%�x���~s$�jd��~�Bٱ�4�׋�V��(��0�����������T�ꛩ�z�+������
�p��>��:©J"\8X�9:c�4s�
cs�f��-���fa\�88>��ݵ����)b�>�q��D
?5��o6���{I�N���:��@6������ V�yHv=ҝj&�3i��k�Qɋ=�V��P[%��#�!u��B�4h��z�T��L�Oo�����ߵ~�ޓV�N�E���~ŊN��q�Y]� �ɗÇO�۵m�<�[�г�=�K����x��.�Yv�g���jjC���OA�KѢY��N�VAz��gڔs:wS�F�>��K�
+����Sj����zp�׻���0�'�
�B�ݨ��W�W�P����K�,�;��J�%.+>Rm3b�[���;�i����;�-�R�q��~���#aZ�i�����p�w~����˦N;sg#��kpԘ���,�����}�J�vʽ�ď������G���Y���7�Ϛz��\9��M��4��m0� �J&�h�����R@�V�ͯ��%��}�S+d7�M��k�u�L4s�,X�it��I�'s6��ӟ�;��lK�;u{t���J?Pf/w}R{�6�m쮶���~a�h��}��5V�.����7�f�#��%�8�u6�z�$ȧ�+}�զ.�(�t�w��Z��zKTȳ����u���f�c��n�k3�l�^��I���}�	��'�I���/=!��s�0Đ��f��Ø�J��+L�Y���=ϗn:":��̀�����9��4ȓ�G�񼺡WRn�<;�Nl������(�D�AIk}O�Q�D+M�����k��"��s�U6��!4rM�~T�����[�ǧ��X��^�G�G?�
�!��Q��'V�?��[��i$E2��澵��.�?��E�J0`rFmI��E���-���T����GK�$ہj뙳�pC;���^8}
I�����MH���OJHhO.Pc���ڵ�@tb��Hz��J���2����_�3�lTͰW��L�Rsn(��ߢ	�O�0#��)�4�.epL�B�ET���@�Me_��
̳9��Sljz��|n1�)�w������̋�-����b� w�i�%����NXo2<Gi��z��a�K�H>$s/j��%r��3���ek���B�$ʕPf��o�	d�ǉ��H�4��,Ϭ�cA��L�Xf��Mo��C�%��q�?�P�!���r ��]�(�0������@����������m�_�
�,^3� '��#�`�/�d����#.UQ~�������!�؝"y��O�ò�Д�gǿ֗6q��\�=�U�V����b�¢�zdv��G�|�[��b��s����j4�������V���)N`E3X1P�q�ac"R\}�еT������p�v\��c�J0�7=��Y]!sv�*�r�hK��3���A��i�؋�N���N\%E"/��%h���OP�p����0vh�%�6U�̞������b��xX�u������HBb_�A���PQ��R+��w�vQ�#��J�L�Z��.��!b������=|��-���i�4$�c�Xrw�%3x����8�%��#��v7쳽�5 f=(D��m?Iג�-pN��E�rk���(s�{4��#���ٯ�1$�2�0۷�����3�y�C�FD�A���%�m0�ѹi�XX	�n��nB��̩�Q�f�5ZN�	'dr��&�ӥ��ݻ��z޸�iDd��p�_�>��sQ�y(e���GR-�K��m��ӽH���C�Z"it�4�(��Z)�ƣ�	p�7�"ƙ)�Q
�/�k���!�����S*�4�U�w�N2�r'�CGm��i��L�6��BL5g#��j۴p���(�z�r[iӱAE�&h���������xR3��v��$eѥ	h�)���nq��߲\�p�&Ub/5�{:��׆s*@����<Bu��0!@F���$�Q���%�[C*�I1����r��Y>�]�҂:�=\ ^�|��yR��r�A6��L)����*;"w4\~aq�Ǵ3���#Y���r��B��Øߪ�L����0�|�����ĕrp�)�b���7ɰ�:F�,7S]�̢o�����O�[�6���&�����z�荙QŸO`0=��@���: _�fs��7� ��s"�	�S#*�Rݚ�dVu�����b-s���$-��fra�J�O�JENoL8�͗O.��qr�*;��&	�����������2e��{X'���.� +%ʴ��� ���U���ޱl_
�
�������$Ei����t��Ϯ@���4�����L{�EΙ�:�;�:q�vPAq5;ܬQ0��^Y�G8@���J�h%�4aJ:"�e�R������f_tk��Ë�˫�3	�8��v?E��4�!2)}�36|�n��ڴ�'?J���z	�����V7�S��R���Na}�@F{1��H�4`ۋ��)ƺ���!|AG�q����{��O��N?]���L(%�+��m�D�g�EٷT0E�wO��$�����,�;�t�t�F��8�r������(,����?U��z����:��p>8!`������zR��r�xъ���C	�u2��]S��{ty��/�0>��K�Cd���a�Q����[L.ۺ8��[�Ccu�����z�}� �N�*�6����#����`fs����������Nܽ��R���%M4x����/óY̭�ݼ��o�8�(4�"m��Nl5�.TXǹ�/~����)�@q
��Y�X�
�©��j��S�v*խ!f�tP�K��	;�<K)
�{bF�Ej�K��WvG�� �th��D F���r��]�K,��x��sF�P��%\Z��W!<F�0%��O�xyq�Ջ�8���ṍ��s��ƈviiVy@}�7��`K/�F��7�zm1���wG����� 5��s>�n�|��ydM;IP�F�6$k�tq��я90�?��i_ӓ���v�Z��@�h���!�S��S���(P�|�z�d��㰋��Q[����վ)u'MJqQ�pp��m����J7+i�y����2N��3|�3L�䘄��������A��l���7E�@P�zH{�lqX�W���^���.���]�|�A�le~�X�JS��$�Z�좪�&�p�A�%2�H�H��Ac���`2�<V ���ע��17��Z<>A_k2�B/�W,��j}��_���޼�Ǐ��K׋���V�	�`�G�&0?d����a2��C$)0��S��JD(�
*.�����Ԯ�6�޸I�滫C����>�fO�,�LX��*�=z�)� ���Ts���l)��ͭ�3F��Os�M��/��}P���.���='�B�&�+�4��2��8jz�%��[�e��J�^%���|2�̃I��EPf6$��P�'�W�2u91�o����Uc��^��;Llb�!:����k� c��w}��爠Z��t���]�^��g���N���#�0��>`;l�n�;��r�>*��.��^	w@�����>�B/vD���(5q����Xp%�U��&+QEʏ;��oJ���	��t���H��avp����I22��W���9�֦--��nɔ��ůiWܓ	�M�Z~psf0���^���H��v�F�ϙJQ#�5a<M����:*��
Ы�>��Su5u�]=�`�Bz���`t�'��7<͇<ۦ"q�O�+n������W��+p-�c<#�a���>�8����:���h�L#ǁ�4Ƹ����W�n`�����=[$���J/�T�B�Lؾw��`c��.��v[�1�K@J�������Vq�)au����w!A$:�DHT��.A���7G�,���i^��mT)�p�n�6�Dâ��?o+j����DLB:j�FВ��"�"�l�U�)���ζ�-��SVxH
M5��G��)֝�����H\U^�pܫ �?�.�O蛹~[���-��d�Z3��-�}9�;P��c���.jw�z�O.���
խf L�OO��g�xzӗ).��u���K:���ױDi3�������B���a���eS>���G�E��n��̚|�,��)��Q�L�w2
z#,+��6�����,~Qu���74O���>�4�����b���H�@m��B>�pE���>�˄�-�7(5@��`8�b�f�L���թ7��`�����h��y�S/�v}�j�G C"7�ŵτAڡi�������������A��SOe%sy]�����*y�h�+�$�(TU]�b�PlV�v� {�/'�����8��!�-��{ :��k��R{�p�n�i�l~��:�q���eN�ox���S-6Yk)��!n���^)�7B>�&[@�6�x�Q�BB����ko�Y�d��ow|�D� d�����O�?��/nJM����N,�� �&��/v90�K�Y�S'�{�q�fW��LW�'��C�XK�bsؙ7$[���D�f���X��	0�fz��������f~��}�8��Ϝ��j��G��m@������CF
��n��U��(��w���R3��\���g��C�8�ٵ�TD���V���������\'�����~jF�f��>�O>K�^���lA\��Kբ�քh��$W�,ڻC�Θˎa�^[�l���S�m�'�*��l*iC�%.�r�:"���S�/�AD9q�䏖��:�R��lK¦D�|���E�0(�,*�Յ�K�`4�4���J�>OvC����t���8�A~�&�C!񯽺����-��s�9t���Sǟ��>�>�m��?�mYSr6l�!L[�VO���v�>��kK�]:��^���E��6;+�?�h�������tJ��QbQI�?- �44�Q�����F�'~�D��R6ފ0�ྼf��U��Q�X�eX�W�mESQ$v	�r�wG������b��#�}��cB�C�{y��zL�섚��/�4��t6��!9i��A�� ^Rg�#�-�� ���TB�quF�����!p*��q3��t[�s�wI ����Ӑ����~����I���;e�h��a_u(���q%@�Ey�_�݅T5�
��>�ܛ��� �������� ����^[낶�L0�LO��1*�8��?�<=2�i/U:�E�3�%{�|	���%��9-7	j��31�/5�#RG=��cC^7<ȕ��=�Њ�q�I	t1��_�<���k��$���z�8� m�$Y����Q�P���u2PxI�=u�Ů��S_�7�M�~�³k,}6�\���� ���kײn�F%�Z�)�E�>��P���:ƥMp���*K=p @dQt���CF��M�����]�Ǿ��{E�$d�Tk�7�
�<�\����k��ԉwsHb6~��ո��
PQ?���h��G���!��*D!iy�12 }�b��Ϳ�Z�铥��	
͇���A�24x���;�|v갦�E��!��,�Vҫ�M�����O����5��5�MM�Ϲ
;Lz8�:}����*U;��=�`���r� 6�SH��'�9�Ww4�/��?S&�^��1=)�ju�/�jO��Iz���z!��o��J�Uv���t�����]]@�+2=\J8���1�D k��%�J{Ѵ����[��_�Q ^�A,��E�5k�gȚ�L%�z2ss�u�P�[_���]�^q��[��������P5���;�T�lG���?��n�l��<q�ݻ����g�M^�LO�>z?G�U��h� "#|/����x�)�)�B~A>3�hr�&��y�j�� ks��A&���L��i�Ƞ&f��v&�n��s��0��͋��?�`�¯��Vޠ5�A���M"N����B]�6l3"�F�W���r��)�A��vi��2i������ȗD��+�+t���]i��n9����`i�JN������3�C������B����	����o#00=�0ˠ�[��O+�Z<�ŗ�����(!�cfgٿ�Ƞ�_�� �G�`LP��^�m�񁪣����qڊ,��0SF��@ek@����UO��K��QM-�tÄ֨ʛ1C<�mf@Ⰻ43�f-�j��Y��wb�w�̗��|?uQX5H���t[i�p�8�8��'1�պ�%\$v�-�
��~H[U`���W 2�[v�M�>��M���M��S��q0l��ȕ^w��1�v]�� @��u	<{�Z�5A�}�wx����0�8i�������~X(|�("�>����$۩��%��N�Qςgm8�d۠����$�.��C��g��pE?�������{�HB�%F���~]9%ּ��׹[�2�KpL��cj� �֜�d0y�4534��4E%ɕ.>�)�d�R�%2I^��k��ӂ
�`�ZNlm�;U��+�*/12݄�֣UrT�x�M�L��9��Y0�"��aR�,y�Ȍa�)��O0��͙C~���_O'���Ef��u姣Ã#?H6+���"T�,=��b�&�SS��޸w?̵�T��>ǧ�\<!�Rk<�6�ߗEM�<eaI��������ޣƾ&���ǥ#B��Q;Y�_}1-���g�X݄-7�%Zb�\��g��M_v��n���w]�Ce:x����n��h:�x�6v���Z�
�?!����[�p~r���r�_n6	+��eQai^���z�K7����`E��{���s]�֋r��s�!
mn���\e����M�s�s_��z�
��n��L���y0��m�\#�n����v[u;p��E�KV�Sؔq���>�`uI����i��|�U��lyt���}�P|��Wb�f4n��8��ڜ2J��|��ߨ��Y�ǘP7��)�$����y#�cx3x�8M����J&-���V�E�1���r|���Q�O�7���8O�Ys��"�ۙ���i�f��1�F�>lA��ɉ)Mߕ��t�8H��+m�=V���$����(
��~zTN���������<s��"�x>�6�^�=bam�oß)�R�ek���̮�T��E*�����*�����y����k���`PB>SB�~�����`S�:��d�8t���x�`<<�k�aWH����D]�Z=���g^]*�xռ&؋��u��4���U��9TB�mrK�bw��N��)e�RYZ~*�L��J֝��:�׶�n�����ze*��}�n�ȃ�kp�\;��?|�v?�fzF�G�lu����B"�4�		�j#�����B�Ҽ��OK�SZxB�a�3w�B���v ��ElG�H�V�&�)��E%ǅ�E^Kd��v^'�M��k�j����,E&��ȸFib6��Z:G�x]dPa9�Bが,^��d7K��&m#}��圼������6�f�d�ɹA��@U���#�N�|;V�g�S�-�F�V�@���i8�V�jWc-K���04t9��?�������c
���lc��C)D��/ӧ&���n��O��1!̏��	�B�R�<��d�s�ዽ&����[�Y��?7���&�Ƽ��"%�#��,���8�k� il@~�n,m�ю�*^m{x��Y�?���y���1�9��u�~k{���w�ĨۻWYa@�G������\�(�c�pf���� H�ċ�>Fg>����i�d"]�p����Dv�fM�aPr�SԂ%��x1�=|r����Ksq�x,^�>D������C���	��U�Us)�:R!���&ZJWјh���]�h�bN�y�KT�/���#Z�����)B���D���c�ۜ:r^?�9��]˚/(��El�c��	�6B?�5[F�^W}j;��Y�ͩU��p��hB��;1�ĝ�;�"⚉'G�)�Xq��4A�$+xy��c(���}E�岉g#��=f|���vRf��)�����Ð]b���!L��b]6�ȄI��3�	�?*�_��|tzdA���oҲ3[s����(�n$�q^����"9�-����f��J&�j��7T�X��p��9Yʲ<�D��`��B�_L\W.��P�S�'��;$�D�����x��eP��K��E7���C���v��M,U,�D)��7I�GC�0��RGY�O��kun
�xuj��້�;c��7=��W�`�r���~��P�W;�&2�2��N�[���*HyL|n��V�8�@�A߉f;��T���������0([����j�~�sۿt��YI����|
5�`��7X���c��n��[Oz@\���#7B@E9CƄr^x�g�0��Un��8�^���I�����w}ǜ;Æ�D%�z4�\�s����p����
Y�HT?��t��y�R:�LMD�u�F��We�#'���*b�u�ÔT[�����]%��a�O�!kV���Ǣ�Y��&����㿭�`z*\E� u�~36M\�q57�G�_]�Ï@�6��~$���Pݜ�ap��"2uF	�Q���y=$6SM�{��=�ԅ��w�I�Id~�{�!�;�'���l��D@K�8�=:h �./ʹY
���ŪX�gK�����?l#dk�FW�0�J�8�mk���d�h>ρ�隃<��C�l�Fd$�Of<���sQ�|2�QF���8Đ�IiP�C��v��Sd�?�]�,��843��x?��g��S���̀�J�Փ�"�H�\ҫqH߷�v���U�U&è�����Kw���*6e�O+N�M��T_�77��{� �Hg�
���&�X��,�)��N������C6��E�����(o�� dw�.Bq�\H8��AQd��a��*��	]m&�yE0�U��U��ɤ��#�n�fG��5(���UEDg�D'Ę>����Ȼ0��uP~N��Kr�Gs̉k\/�������2�����j{��	�|�fvxVq3��%���6$��#a��ſK��o@�V�㏠��׆��Ε^Ħ�W�P+^#m�"�Eߣ�d�'�_����4/	�����Պj"R��̋���G�-ߩmN���p�Z�D��E)�ָ�1B
?h�s�8�dќ ZX������('�C�|�Y6x=zް{�J����		�t�{�z���M�iu��1�j�%���T��g?���d�|�;7E4�2�J7@P
�+��G�f���s���f?����;�8D����ܬ��"wd�����K���r�Z������Z��(B͙�'�����Q>�t�Uy�kkt~򿖍���ڦ�;�t1�����O�@�5�5�ƪ>�ȇ��ۂ���a�v�=���N��(;�!401{�Fj�ę�E�����&��s%���.s=�f3� 5B���W�.݂�'�=�E�����=Ý�|��F���[��׍�Lzg�����#%
}�����Xg��ԨTI�9߶uue�-$~oQ�f'�B�0t~kQٯ�Zk�Q��^�6Vk/�9���EB�Gchm�+��5��'w$�u���Bv��.ZlZ���l)i�`��	C����⺵�>���-�ط3���D�����ޒ���|E5[hk��3c�~�؇��T�����`ߪl����=u��V{}��0`�1�ƧGO��H����;^Z'D)ωj������c�Q't �����e�E]�B�+|�̯�!/�Xi �i6py�.&���&�e"A��-^i�US�X'f��߆S�`7�� ���'E����� �f���(�CQ���f>k��G����>�Uc��5$��صؤ."�%?V욹I��/|������­���	s�b̕r϶�r�:�Azi�� �z�g�`|Ѥ*kS�CZ1���d"�jK�gH𸈍Hu�4����o��һ7���%��[%�%�fxgڀ���S�DW�%ُГa�0�/�|p �U����}hV�Ӂ~K)�����o��]4E�����z뙛]�������;�	������w�Z��C��|�Y�U�7��d�=�+�d�+�rN�G��8?�)���_ۺ��o�݆��(yD��(���N�)�i�0D��z娩�,eu"�G��������]b�r��mc�ZVV��_�H�2�Z�e�o��ҿaJf�l���h�i��&#4����бF:\M�0�̙	��JϢ��VD��}�^2'14VE�����N�;�;�h:\������<R�a�W�}��h��*i�����o�lxP�Ɏ�>�88)�j����߯+�#��Q�3ϨW���D�	�qD��Zv���3�
�T��-s�p�t��/�FG@�	p+F��Y� �ZW����Ae?��et���)a�:MH�V��/�`7��@k"FÃ�J��ۼgwA�{�.�3�ԏ�/���Z�]���I��ڮ+�KkI2t�b��05r@�7�1m�2���S6[1~���ߎ�6�s��j��?�j^�&�����'��?#���&U�α+T�0�k*���x�+Z���m$x�2��&(�&Dc�v�bv��m�t x>6,��
C�@�/��p����;_��P1Am>H����*S�%����a���H�\�M�f#=v��s.�����_�^����xX�_u-qY��}��ѽ����@��Q,��̏rg��	?�6/�A��	��f���۰ڿp��V����9ъ������m@]`ކVݢ&;?�����3��[���0��&A%v�ar���Y�h����o��˜�@�5�YoP��Z^�!h��:����N�s2���n��8m�_@�l�A�+�Y^�+�{;�&;�d�����#�N�������^��x;��Z�b��쨇2���c�T�֔,d�Ѽ9� ���s�ɦ�|]5��Q7<4#d�4���;-,{k��Փ�u�o����I�08Z�J�GQW~7���i��|����ޣ�#��>��e��KU0��Bd��,i�;?�~Ap��u�|�o%@����|��"g̎�i�:���^���[����<��SY�<����	i;i~i?���o�b'�g����D-]���1��f���ڕ˓�'�+��43�F�ĺu-�9��\�ԝ����)_�S����%K�I/�&��:�M/r|�qم�ʘ*�{nu�:1�n��|�R��;����XKPt��g����1�=e�i�Q����d|l���ќe�RX���ǣ@.`�@	�n�C0��3�YƳb�O&�a���[��ܑA�\������������DkӤz�Y�|n�9%�MN�k�r��[\��q
T2��_>���?�a�ެ�6nb��Ʊ�8�{��ţC��0��}Yۮ��[���=�)�M�n��©�5���W������ܶ?���	��Kȓ�$�(��+�e$8��C����`���/��q6P��qn�B7#�� ��>B�l��g��U�\�{._'�d�'UI�]qs��!������@� 
���o��*(�N#"�7!�\���1���ub����Ͽ��gМ���B��8_]Y��o��z~K����g11�O��
����ph��G�r��O�T9bb��4�2`�V�����K��H��[���`o����g�*���054��?TG�!�v�V���1�d�wrn�o��)cJ�Uz�g��f��q�w��i%V�1��w�U\�H�v�H����X6g�L��.`G�W��*��8#�ʉ4���EH���f�6�T�n;R�U_(������t`��\��8�z�q�-)J�~9�P�K�ka?��ٔomD>�5�X��3%*D�C�)��ϔ�r��R��o���e)�d�� ԡi����(�i��A�D�D4y���������{�c���V:<�&(���9�dW_���vШwG��h��Q��#&ד��t�gįR�~���C�?�@���e$���럙��s�he�훠'�K*�3���^3�����qEYk�n��v,1����f��%�A�P�ok�';T�5��,"�uߤ
Z��杌ۏ��������C9�T�b�m�e��"U�-t��x�细���"�Q	J��,]�����Fk|m��20�&���.��2=: �ԕ�7�S�r���t{aVy������?�+T4\�����T��6��b��8�������f�%O�I$�B0�󲪃9==��B*(BT'�I��̳�� �(@(��lw��� ��Ԟ��\��z�f[3��������2񩮅�y�7Sد*+�ָpXV6W/W��gȁ������M�/�w�3��p��Af� 7LU�Ѫ�u�Co�:c���.`������� _�P�O�X���M��'7{1H_����pį�����)��E��f�k�x3a���ܝ��}�{��	/�I���������ؠ�N~���׀P~��Ջ���;�,�[�bǶy����Hr�+�X�dt~��iwm�/."��F�aI���y��&�<��w�z�I��˟+�i� 𦏶�XMU��-|mdh��5�{�ܸd��%:��i��n�R��"絖Bc0����/3�o�'8����	P<z��.Y-��s�̲�_�8�d��Pe)r�l��JM����'���|�H����f뱲p�[sn�(��Mڍ�ǔ5����{M�q�8s�-0�"ݙ@�(��Q[kۇx��	hs���%�2c�f�� ��-q��r�Ӑ�>><3�P������T�����/J��3��I�:H۾�1���i���]�[v��k>,�}*b\~����#R@�ꌠ�]�p]�	���D�!g�a����{LS݁԰��mܐ�,w��ʺ���'Yw'���:8k<�3�X+-���3	<U(�(ɺ�P��Ҧ�pe����	<�o����t&�.�٦�t���\[bD�b��
!������Θ?�^Q�<d�ѕ��}J�y"~М�Z*�r�մ���0��&�	��PSP��u��j��B�h�G-,�̆X��Y��3�S��\�G�t�ܦ�!�e;�ՓL�j�e둋;����_(de�!Qy��rEB�*�A�Bĺ���UW�fⷘ
��	>ȪU>+�����h��x��TQا����m�	*����zf����2�D��(-"¼�i�����d�����<R�@e;����ҽ*���}�m�T�Q
�S*��0̪�˔�����)y�"UD�A����8t���ר!�B��Q;��2�%��şv�^M�t���o>�J_�ãH��Z��*�ǿD��q�7;\qJL�qs{}I�����N7��/�dWK���u��O�׶��r,��.��K���	�v;)���GЙv��ҬvoEb�A@M�6G�f&i�nձ?~����<�c����)��ڂ�)ү�f��mJ��C�Z[?��URހ��+a�f�UU4��V�T4����x���?�Lg2�\Q�ͤ���H���s��Z�ָ��Z=���x�X��u*�v�b�^�W�x���G��$ߣ4�5[r�D�TM�`�zK��{�7d�=N��̍�Q+l'�g�zB�ᶓ�uz�v|�\��G ?e�*_|Oڟi���ѳxq��o낷���-I �b�E¯6���=3d�ot�a�c����������U�윊de���
�-�N�l�s��?���;.���[	Kd[F�>Ȭ�/b�Z��]r�MRuǳr���d�g��G<��¯�@C'T�q�
O��]�+�����k�ˣ8s�!7^�O����3m���'K U(b��/z�s�@�n��mnA�Ygr�	<Es�vP�̂��Z�VZB��竉p߫z v^M=�빼U?�Tgȕ�cZaS�)��H�~^��c�z�����XSj�b�b�<N��?h�%@���S`���g�m�"΄	�6X��"��~�;�=�u�$�X���GyĎ�<��w���a�&ri}�ʩ�r�$�#�Ȍv`��%ބ>�r��B�,״���+�y���a�e:�OJB��P�`��q�wZMj�ZU�*_?�g�!��I���v�I�W�a��VF%�{��	�~_�`n��1������}������
�}?��>�����@�hl�*$�p���R���sSz�k�%���^�_�K����+=���� �AKn�a�ޜ�<Of���n��ˢ�[�R���}��H;���; �#0��˖��@��F#��zP{O.͵'^��VةX�� =Σ���,L�ˣZv���si<6�	��eU���xe7FTc$t3�Wt)϶rT�>�ƚ$�G�V1�t��=��-͌/.��>���9Z^���+���'��O�J���IS��Yz��H��%�EƯ�`�a¥���y������P'!�
#��JV��:s%l1䁨v�Z�#�;\AY�W]'@Ӕ��С���'�:i����l�_�\x���y���T\�]�:�Lc*���uWx_����jBukP��P�ȍ4_1��R�SA
��+J	�_�T/p�F�m;��teg�8�*���$�@�=
� k���|���j%b�+QuUM�y��o�^<�]Q�[��-^b��,�n��4��a���{��r���=#�8���&\ݯVH`�������I�u񭈎E�R�.o,��US�hv6�|��B�NI>�N_��nnw?�!�Z�ߣ�l�K���1����*��� �J8�x��6�o	1�ko2�Է����mQu<��^ aH�>���G������������m#_u��H�U�H�l6i�S}@���w��w���`��/J����qv$]Ok��ڨ���!b��40�L����s^�{~������[ϕmʦl���r���c�k��������4
�~��;�LI��EK�<V���­��f��Y--`R���$�t3S�	u�(2�	�a�W6�S8�d1;�ύ� �C�k�B[��wfi��irm�
��(�>�f�U�8U�rHbm�?Bi'��^�?�������L�k�%*���z��+��ϼ�C����'i�uS�m�H�� :�Z��a�g���� �X��2Ø������I��} �n]�/�K�\�)�\�����Vx%�I@�H�`�z�U�t/���{�1*�#��	�Z����2z�>�~���|7��qD�¥��v?�Q"�=&Px�����%(���Y7yն�->X?���Ӫ�ވ��d[�g��;,��,�6��
��-��>S�1!�m�_f.��.��˩{�`�Z��j�����L�ؠ�P��"�ud��^q����	�sR���_�,�I?+�t�F;�G�������o�_�0��N�Y��Ew����la��� ZnH��1L� ����~)�9���۵S�A��AH�㝼��lw��H���C!ւ�Բz��Ֆ�3�;1f[\��aҰ�]�ۼZ�2�N����)'�����oPj��]������Y�J_jЪ:éfQ$?�C�U��{l�\�ԇ��i�Qޙ�?h.?)�PMT�)ictf^��y���W_���쩄)�B�_Y*��,,��+ߓg�ưu`�{h}���U�*�';�U@j{}�]�\Fid!��X��mWOb�;}|>
_�7��oCrM�W����U�t�3�����U�G)��ɸ� q�79������3�=��%��H
!h��T~����h��_���/�Ȇƣ@X©W�S�X���r���(�ѓ]	2�t���	�>��H��;H;�8�y@���Of����?��xO�IL�(���ĩ�@�������r15��V#�k/,�5�N�<~~{�))�sX���������\�3V=`��"+����&eI��u�'Z_@��ب�����q?Y�ֳ���.�_Z:n��~C�ym؏���uĕ�6�?v=�l��{���Y�]�����?�������uZ+��Uc-����F`aȒ��n�q�$K�2�8͢�۟����}�(��k�RIê~Z��N�Q,�>!((d���uC*��'���e�����u��"��l�4I��nf��яؚ���;r[r߫G�ߖ{e��_(�ud�m&��$���t6��l����
q���~sbh�{�6��o��|lV�\�V�N��$C��5[Q<`_�8�CK\�|�v��A9��%���ޣ�xM�p�@�&�$��X�x�6��@|	�w!�}���~�t;��j���2���ٜa'o��FD�?�Ԋ"��(,������̇�i.^��@�2�KJ0�e]�
���0�B�$�j�!�c�����۹�[$H]���f��hk�S�܏��/)��)�4	��7�m����#.�4�_"�t�A�#��� ai_�^!�3$���ԅu�Jq!�H����QY��ж[_��}+�,��/�x�ב�~�Rhi��2��Ɋ��e���(T���%��q��ɍ�s/��L�.U�D��@�=��S�fHEu:�*�����t+d.WKQ�z_0�mA\��r�-|v��͗By��0��B��&C([y���sR�:�UR�dI-)��v
9䭪��6�B�`؎�^濉�b13�0�*w�<h��4qҊn�+�ҬMu�u)zl���A��&���� �1�u��6{�����:���� �\
48�]��dh�M(���I����D���9��2���v�ר���O�WBܨGNVˋӅ$0��|S<��ƴb�x��������6]с�(I�� 3
�ur`ƛ���y!�D�uYhS�4a�D�>�](��
t&���aS��Э�P�xW�H��0n;`�aǌ�oS�m��k8Z)��%� �J���w��K��h+ݺ��?�:*�P	Gv��l	�Ǵ�^���zW�.X}"e�惉<��T{h�G,�����)�pFg�.�K}����}tפ���~�2l�c�NVN�46��*��� ���0[��XM#_�,�[��k�R������u4���������9w �n�Ki�ޖ5{ʤ!�������T�E(�\:� �cK.T��"��c��_p Lt�� :tM1�w��Ϣ�v���WM��fLWÙ��zI��ܤ���G�a�%��xg=�z�,��
ж�ìƊ�㉢=OT�V�B����4#�H(!q��zR�'���\�|�D�pQ$Al�'FDZ����<m�(z�Ġ2(\��0O*5@�HAp�mb�|�=Hl�`��!����C�>�=K�vOR6W��tc{t#_E��ӏ�5��ΤMk�K"��y';�n}����%2�n֙��S���q@���J�#c�C@ �����p#���R+wUS^7x"�KiN�j�?�[��V�%���]����� ���B�	 P�)��y$��=X��*}L�;��=�"1�_V����3����>��e�CȒQ?ݵ��n�����1�%�5�-	��U�>�c���<��g
���������e��!\����{�� )� ��Lխ��q�K�֮�|�r��?����L��O-,,R��km�y\�I�
�T���F4}�q�]Rc`�A�ϬmL�c'��;i�iI_^��!�BWsIx��[T��"Gqo���eX ����QR
��=�PT�FD%a��`
D����o>&�@1Q@t_�8���B������HF�J�yzX�ld��
·��.��϶��g)�$J��2/�ɇ7�j\��.������D�ޔ,ڐ�؄'�2�`� ~�[Fbw !G~_?��\��6F��;6��v�������MC�ȋc���>�G��Y���K�f.=���C:|hy�Iy6a�nB����=�>�%ÅH�q��O0ء�v޼+:�P#8�:�b ����խ��ױdd�$�v�^Ќ�nxt��u��~�p  ��ƚ�b٭�Mx�[ϭU�\! ��c�YlY�\��͚�R#[@�^���YY�����b*��:�z��>�Q��>�*hpl��oRV"����*�<����3&F��H�^Ӏ��K���yD�B]�ܸJMy���X�fO�۟��6��~C�o�^�b<���L_?�	��6�� 7x�׸��������d���w|]ep�]<���
)���q	a�82	����r�ϡ�`�p�k�����i��֬�#�#Im"p��X�(���f2��g��� ʠ�x}�^�S�~�#�Kj
S���*�H��k�%��[�X*��BAe���g,U4	����dɮ���p���{�##¿c�4�L���m蒒���0!�M�+fܫ���o�T��^qi���d��'y�L>ڧW8
�p���)���F� 9n�O��Ф�{1#�_OQ^��;���@:�ֆE)�	5�Nc���i��7��������j�����ψM.}�N��+r�:�Qk"|�E �GE��7^w�x>��u�j�)��w8�`���򶜪f�jU銰f��_���.v�s�S��Zފ�뺈�bO"�_A��b�2'<`@w/�E1�:I�-`�W�Bdt�1�?��Hh�k��lk��S2�	�(p�����f,�+h���;.E;�E�6j%4�li���_҆�fh{_�K57R����8�ՠ�3&]�0\�&
gN0�(̻�w���gD���Z��-�U��@т6���Q�U���m���N�~���0k�]�M�!֯f2�AC	��m��u-��v>W�Q��iO �k�	Y�4��� ��{�<T u@J�yp�^o�T�8�t�՝Z���W�}�s�+��스���ʻ�ރ���sM���+�`�'�%���j'�ͦ��M�!θ@~U�%Yz�^ozq땯�]W{����m���)�4�;����,<��8WX�PKR��j�Z%�#���1��K����~>omm�I�n@�?�BaM���`��T�.�3������s�k:�k����.��v���6S�s�ilT�C�.�(/Y��- y�<��u_&�����*�} 0Aj��R�����{�FP��<�_�p�g��!����k�G<ߘ���c�L}��4g�F�G<ѐS�#;�9�ve�I+&������H�D���^r�IQ@� ���J�մi�ط�:W��N��O`�T�Ǉ4~'��d�X�넔�yz���fE��`�9�5p����|h�����yþ�m�>4�NSX]Q2�޶!�&���,�����Ԑ�ύ#�#�WE�˖��X0�Ac8�:;�\�k�!�a�d!4�\�S����_hX�\,�&@�2%-1�by�����f�R��Ɂ�K�T�H�7���
�/��Hyc�����G�.�l�ӋYS�["=J��pz��g��]�E)�M?L��h>�@����t�a��O�JLN^�Щ��d�{�^,/�+D���G��;��F��ڄ��<�5�F��̠����#�����M�~YL�,L�p���i��_���%7�5tA�����ﳦ��A%H=���}����[�\�JŬ��*g��ɣ$��цï��B�cd�g#���
�#lX_RД}�cke=47d�v��J��;�'U`Ze��7��ʏ^I���ؘ�Q���� å�cͪU4����7���� �I�1���Mu�7��xrO:��)])�q���,^4����lt^E
�l��GEY$ �1�����+�9��nPiG�!GM@�� `!���颺�؟�2�J��fG�ɐ��!��n��J���XsQ~EHRs�ʥ����m���'ah8�����}�zi�(��4 ��ݍ��/���0���ƯV��l�#�F�}�m-	�f��Ylh��������}��h+�M��9cz3��	��� ��&,�s��B�7�iR��xm�;��s��o��[����#��j�R�p�-lX#FC&f����o�SO$�;7��_G��z�lg�|���A���m�X���4�-N�Ή��f\�ְ�\���'�{�T�M�$�W��X��ɍ�3������֓�Ӂ[:J�4Vp����
���p�栞���ʧ"�}�q�s�����C5S�Ü%�o����ljJ�R�YNC�'�2�V��n�����s�j`��z������ơ�
0\3���Q;�<޵I�/���1G�����Cf�[��:���q�)x��z�\(T�V��@�hF��1\�n��Y���O'�I���0
{�u��̿����I�?�8����
��*�`àU�� ���0i��ǁ5z�_f�X<ܿ�]��@�u�?����z0�`u��$���ʒg&ۢ��37�q2�Ľ-9��-^ E�+D:�̎��F+6s���� t_&���s�jcPc������\��.�+� ��|_�����E�r�d��G"�Eb\ı<ݷ9J=�#�2���mJ�~E�L��^��ַ�1ݥ4t�/��#O�!�_1��Cu�`(E$%{E�� �����]�r�|�P<|]G��@"��+)��UF���e���������=(����O�Y0�������@0��/��ڋ�����~��1��-M���q���7xK[2�6[$�R��ϼ\|�-��h���C�p��1�/(��@1���_Q����-���~�(�\�Ⴛ_���ݚ�TL�U KY���M�T�	O�Zl���:��`BD$snnv7�,!Z��!}�2[冓��϶����whxo���&/�E�;�J"��S�l�O���`"��/kMN��`>ӹD�=e�2I�;5�
��.{�'^��5W��ñ����6.�t�?HEA�m������2�g�b5�����v��������+Q���ҍ����f2��v��uI�Bf?M�VV\ }1H	���o�r`2�)�m=��Ւ��*q@��U��?P��a��4^�f�`��d��ރ1Y����V�� �������O��D%$;����sb��~�mxWn�}NA�E�z��a����3=�RTm�5BA�L����"�Zr���1�J�iJ���F��ٿ儥飢�n�����Gד���F��4w���@�g�}n�8�MZ�<͂�Q���r��1�dt�(�ˌ&�~k&.���^��"��ki�Wg�૮=���Ͻ�[�P�^F�x�Z�$O��
��t�Ws�)���I��W�~Pt�p�t�:�����V&��kt�"/��0��1��/�^����Ҁv�e�����Ζ��
#��2(����w��99JGμAu�.��8�r�z����´�jz�X�[�O��9�s?��>a������_Ղ5~�#G����.�`Gt`}�ێ�E�#L�ẜi�:�����-���A�Q���HH���2��@����=�r�
l>ⷸF?Q�"���	-�<� �{$/��ad��'�����pd�4o��%&"��US��'�b�
L��Jiq\F�]o�:�1���K��]����:	MJ��B�y�+[fQ0$��XY,��r�!��ҁk>3���f=ĝrFd
6_��Jw^��9yhE�?��,j�!��@o���l�:g�5��� N2��z��0��
}�HIЍ ��T���y�l���.��B��)�x�q�2'J�h��'KGIh5(��h%��NR�� {����`9U]�Ʌ�7H_ _�[�E�c;��ԓ�\B�I���n_|�q���j�?��c�~����%^J��H��'ʼ]f���3W�!Ye'-�ߟ���K�
����RP�������z���e�xNҰTd���>��4[������q��J��A�ſ�%A�^�>F�u]>��>%wi��M��gyn�@24�%�f��w���#�g�d�k�Zz�lV�>��SO��{<��#$�!d�J#`$�~����ppvwZ�/�-��>�,�3vQ��NU�4>�_ը��FSB���\f���>	�~�]�*�m�\.�Q�O) �����xY���f�mK$�l�wN)⫰O����������ȸ�O�\�uFtXY�)�3O0�<�7d�~�r�����~���)F�b��m�U  A��C�ԕ���q._W�k�#�F�t|���x��T$�b�8_ĕ�a؂C�C�k���x>�k�a�"e�[�*�w��es���DO�K|>
yC(�ܳ��i	$��	���ת牀�X�~%+VO����L��qX��1C<*��^�]�������D�i�9D,.�PA��m �r�k�1p������w���_��؁΅q��DмvP���ڙ�,���n ��A#\��ݨ���y���י]�Ⱥ���`��ϡ 8�v����,j�X�#Ȼ)����4�V���R�}PMT�s�-���1;��A-q@��,E�i��*��nID[+���S,p�<C�Y����j$�3\V��o�M��������R�3��W�0\/^�qء��6�΂R�p�e�S���4=Å�'�w������ bG��w��#���[<4�"�]9�	ܥ�n�[!�^���M��1hHg���+ğ�Bp�����F{�l�?z�5PN�>�@w�	!41�43��ܤ�Lx���9x<��]��K��Z�uE ��=3F��M�Vl�����p��w�١'R�{?�T�<�"���l�Z�0}5��)����#5�M�J��o��Q�P+�6,-��̩t`���Q����*P��}�Y)u��<v��A=�o]�ES���@V�y����t/V]�R\�o���|��P���p㨬��7�`ؔ�+w}��`�&�o.�z-��"�R&��"2��uB�e��9��P�VP�8�^
 �г�X?6v:�hA�c���\ K�Rp���`�I.x;88�'[��9O��]P?i7���d���8����ч���0�X#�D�� < ���QVL���	�Иa<1]���y��BH�yb�I%�Y u��	wK�a4�n���}Y��Ǻ��-v/c ZW0��4�F��g�L9�*+��{�
���$8���������*������R�x���@�!]�]�^n�Y8������;K-���?e>Y�hl�#�8�z/Jڗ<m����w�]�Ԩ�uH��0/_�8��x-Q����J���Px�,��Nn��P.���`�b��C����Y˵�"Nŉ1� Cu���a7d�_)? ��|ߟ�t�7��ʝ�/+*1�bڞ�����#!%���t��%�s˃c�p����zť�)�#�*��&h�0��vG��y�����uR.��(TC�P@RԃףcR\����=5B� **{/p�TB%}���}g�p��tL�L���k��\ ��������l3�w%����ح ;utG��A�,��BXIM	����]�-Q�T��\��b_7�G;Y~�",��)l����\�k]��1p���촯JZ�3Q\�	�^�`�h��]Z�C�{&����]!�{��� 5�E*Íp�~�_�G1:5��A�:Rt���:��~��/9��Ȁ���nH�C��S��AZd0���i��䮇No�&�E�����zݷ��~���S�����Zn�d�z>p�g�1��W�v�U���L�U���h�"{Q�������)_U�A��,�F4|����$��{ˀ��!����K�Xl����i��7!	���0G�BQ2��	�髙Z讟6�I��7�q4��d���_��e��~V��1��P�9�ٲ����VM��_�j;�)r9��[���H2y���Qb��ςL�.y�D�n���-�VJ_&�Y�N����1h1�Q�Y�Ӆ��%������^��I���0�u"}}vJ�l�д�_7
�_�&ؿ���?�i���sEr��_��y ��I�M�I^}���j�c�����GeG��t|�;1ѿZ4O_�.�U1Q4�DKӰ��6�,B��K�x���n܊���>�2c�A�x1��q�g�_n[
.���.G@��*j�]l����\4����Xc7�k��@�;E�D<�ިf�]��Ѽ������<�*��6��?��t�K�����R �H�(7T&䓋w#��]�=J��ɱ�mex�N�y�����s ܤ����xc��m)z��P�v�����Y�'�
�f����V�'����3�M�<5:e���󿚵�&'�Ωz��������V��T�@!�Q�kc���T�A�CKq�� w�|��.�n�g��x,�
�H�MӁ9F
���L,f�q�k{x��2:��O)n���"�+��$"�9��z�!��5�.P�����:���\��X��d����ΉC�YTx#%k{]���Id�k�P*x&Iՙ����	2��:��#	�a7nq��oؤ�q�0��1��b�O G�T�#���^�X�֪C�2_d��7����
�i��og2���jy��!
Šה�=�Ѳ�N{3�W>h��]i�#��h3�H&��+Yd�~�`�^�G~7����?��'lm��r�xXKZu��}��D�$�XE\Ϙ���M@��A���V6�T^c�\S%g�F/�utD����c3�;��E���zt.d:j2�.��D��}v�(��yA)����wg��to��fFA�c@Ј�$�̜V[�(�-���'�jZ~4.�|.>��F�R��_m\� �6V�x.�v.(܊�YT�Bn$���|A�LT����xg	|��c{�>�5���ؔ��|u:,X���z��4�R�����˵���4�(c�4��v#b��y=��7�	��������եW��8�}����I�'�#r"c"�8�3��u{���0D���)M(Ш��E;?8-��oOf�JW1��N��b�߲	�ũ�|,�d��];�i��=�;[K�*�u��P2����-Σ���=e��Uyၖ�+؀a��N��ȞQ��>��צ�.��f��x ��ns-1����о��(��\���&�7���T-��ʆ�6N�pF��;�$S0Y�kq:車��lJ�h�#
�!T�f��\��G�E�c�IM��Q�����"w�3�A�lTa���D�����g"5�~�&L����[^���d-װG|7�2IQQ��H��'h��Dμ��&�PH�l�zJ~����af6=k�T_�E��vl��Ʃ���N��6��fk4�#�3������#�_�Yz_�0���E5Jڌ�C����(��#2Om]�t��^4;� �2��ȭL5����vV�j�[��`��l���<���5C��n�b��C2ďg#&a~�q�d��Q��u�?=��y����9Nr���v�_�@��E*�,�~޼ �ڠ/�;�B��j�S��Q��n9���ò����=Ş�ʱ��%����M.���:��8�1޶U��h7l�=�OQh�U�I�@�=z���lń�ks-�!h@�'x� k�\sr�E�¶����I��Y�J+L����ze�S|��Y�-N�}D�mW�׶�<��K+�(;* ��q�j>bx�,<k*���fsvr2�aN�Q�W}#A�.�L7F�Y�d�f�}b�Y�"��b�$tw?ڀh�q�}E�-V��ޔ.M�T��s|��V�$a&�v�oD8���4���i�����J,�=7�vB���ƚ�C�X_��^$q�W�mM�:b� �v�V֛6{nȉ�o�WŴ(�C����MWm�N.��E�	I�`�������IGZJRW�n���%ެ���iPŀ�c?�ڈ%�/Q��.��HY�x*��{�����z�(��dv�W��i�Qv�{�z�6t���҄|[�F� UYb3[�-5���`��4 E��jA��	aB��u�˫.9�����Xu� �����:�BF!����`�n��J�}��.4�=� {�R�O���@���F�A��
�I�5����2Z* ���w�i(6�Mc�򚦫���\�Rl{U�2N����,�J��K�8�4$]M~��U�R5�%AQ�8ko��'���!]�w�}+0��}K��� � �J/u=�:�R��w��uq�k2�<�ދ�\N�a��Y\4�Y��J��_<�������Λy��&�ll�1�j뽃�H�NJ(6]D�k�V��v�N��L`��M/L#OOx~|�T�( �i25�U�6�$��T����*�R�z���ĕ\��L7��سP	��DW=ADL��[���fΘ���!�F��yú�u��Z��^o|��-��`�נs�G�z�C��ת�K�z���q\Lx8��f�:ux�$�.�Icr��t�6�ݥ嵫*O����ZmmL��;�&�LFs�杫o2؝����9Fޅ&Xٰ=<���5��z��N�n��y�KI���7>����{�`��r�W�A���
��U�����g���k���J�4�?W@֓�A2}��(L�w-��IM~ڧĺ[��&��;=x��K��"G����M��-Ï!�7�P|�e�*�ƃK�1��hGxsx���D	-�M���`�e��(�9��x��6���|�(�s�6�5⌣nf�@QK�3������-%�e��#��>�w.=a���܅x �.�Zv�ط��G�:/�ț]E�?��?`y܀|P�iNFv� 1�� ���X�̷�Aً�g�=���Ĥ�E��#UT�H��4nv�[C�x�7!i���PX�Y��v~2��A���G�3ݔ�(�<:y��b����x!�4�&˻;T�A�0��
��R���@�b�r���aSZ �v�5d�i�L��<^.��g���#פS�6��\4�ܛ(r�W%���EѻoT��ǮԞW���9�l3&�����SI�C��^攛V��$ȣѾ�G$��J#嘷�r��a���`a��V���A�S���4���}4Oq��/�,M�1(ޱ��&~J�;)���,}�{҂4�0�	l�oKuL��y�v��b�-�+�D�C�O��W�x������I�v��f��M�r�/�+�M̅�3+-���%�m�iC�Uf�P��j�d�+H {�&j��%���'5��%L��]��48�e��B���^�y ��폛�i<�;|�c��O��ux�vpʞ�[�	��$.��y�������� ���P������" ��]�5h�ܲ�x�~�3���~��Z��������EMI?0� �r�p�����5�H\j�<�=��W�����)����j��ҚN��v��壐m>�\�����B�j%�� �!���1�_le��itg~ދ��a��9Y�^ϝ�
<���^V��Gv\]ߙ���Y�̳m�U��ѯ�#w���%�h���[�F��T��3��>��(c��[ʆn��;�j�z����E�p���Bsa��S�j��2��-�N-<<.K��n�kЗ?/}:�-�;���&a�A&SQ�S0����c�'"�8:�ާ^�� %�R��T��vD�����д%����Þ��d�����ti-?�mȞ���u���C�aߠ�֏�S�R!Z6c�8�%�B��<e��CK]`����?!�gW~a6�.��o����(���IBnx�O�P�A-1E�Su�U��= 9洽rwL�C �eðC�wX^O�\6asM~�0'�2������0?]��z���p����\1P�Qj4��_���A |�$�vFOS޻��v)��1F}����u�P��x��f�˨��eJ/Q;d9�����8k�����0��e�dHx~%D푠��b��/��I�{�y�x��Sq�)F��(̞���u�K�.4��@#�{vF����"z�U��<�o�>e=c�x���peR(^k\�6�E�g!Sy��̽Uc"��%Qo���^��q�Ӷ�Ů�p���W��FD<��c/g��7�~9��V�S|�����2P���j�M;��[~�:]��u\@��YXtّf�W�ar�"=%?^������X�m����w��_�P	�1���L�"ʄ#<�����Q|��/�,��uZYa5a�hR���:��j0�\���K�铄�b}��8/�,I؊`>%�`��S�WkЈ�6�'�ڂK�8�u�����ߓ>B��;�n��/a1���7�&.ň`�.\��&p�~.����i]{e#�pN����G$:���ĉ�\����k�
FP����S�j-j�A����^��z����M5�7���1�HO���V:r
❥�l�|�bJ&���V�p'/����h�X�JPJ��F����ޚO�yctN���`���`u�ܖ�E�)�A�x���P'O�U��Άum�i�/�-s����{8I���p�N8���uId��vz:�B���A��xK�J��19�n��{l����(n7r+N�	��"|8%�њ����"q-�I���X�s;�d���9���@���,��r�V�
a���C��W�����M�q��x��QQ�c�q��?�9���1������S�=�S����
�pt�Yz��ۦ��Æc��E�@Q��SR��U�|���l�����T�V^=Ү&�(�ۆV�jZ
���U$�K�Z�w����Cl�:Q'^�t�\��8�߅_}�p_�}\�#��go-g��$���l;A�V�B%��R��@Ξ�wt�� ����@m���#m]�Ej�	1�v�B�h
^![��#�+d�ԑS���C�����va�
S�Z0���]��E��N���\��J7]�s}|~H�"��:ź�c���%�1B*O�ŌnU�8�w��v�Vu|=רX哾�}t���Ǩ�/�8�GkE	bW&&�R���C.BK���8�s��P�������w3T87�j�gV���H��Ye�K)�R��͎�%����>q�C��Gޖ
1����p_5++/V�a<7����4g&����D`*��{���Q�d�������������O�YB26R�=*ޫʠ" ^��ȃ�1<����`��T�cY�/���!r^�@�_M���$}�z����X��N +��(C$\�%�Wn�ղ��ӞN�hN�NV>��A��4�v��/��g�(�G�`���u9c?������"��j����5Z���`C~��(z��zR�M�$!�� a���;쾬6{��,�B��FJQ_�`�\�<��%s)�_��quծ��ik�?ۡ�A���p�!�Ǻ��2@.�t%(�S��}e�SJ�>����Vy`���m�ΰz�*���'?-���F���z��82Q����b�M~�w0b]���s廦�^Du��9�#5�x�d��\E[����ESiEIk��vX.C��ЬKuŁ��3����=`�}�ɖ���	���z��3�*A�'<�&��5SZ��uYoOa !;�Ԟ02��R�GL�O��`U��o���W{�6��=�!~���߮���.z��%�߽h��ѹ��/(Aۏ֐*�g�>���h=f����dl�)���C M�l��R�K<9
��v����q3Yߊ(/w�1��@�p����A�@�[V'�pa��Ɇ���
��RQ�3Å�LP�k���VC�e�J�u�@�Y��v�FNs>)<�Q��`CSl������4}?��G�N�V3�k
m�#"����@��Ȉկ�B��Y��-n�*���4
w{�LVgj��Dn�ɠz74V��4���
|g�s�D��ɝ�l��~�M�����6��5)6�Lz�k�'��fk�S_�Q\ND���j7�q�g��!��R���R��-��ș.E,S���Q�[?{��;�\�5[P6A�xtDY�|R������^4͎ 0�{
\��֫Iė�~gz�g�!C=�y��x�Ⱦ���h�H��愁5bv���7 o\�`��ZsB)Q����~�jL��Ɍ!�7����h�5(>=]�BJny�+5RWq�ktxZ�ZY����c�Rz��~n�]��F�<y �UZrkZ��dȓ�IGȣ/7�nT�w�T��t-Ls��e�����a�MF���AhΏ�d�h��O�����x ��G:׹BhW������?�������8G���F{�'z�koī�&�|�7?Z��r!z0_y�2�Z�xq2ccT)66��A��]�3�S(l@�Z��/��䖦�Nw"���sR8�E2�{7b83ѩ�Ce���=�Ƈ�������t�xx�Q�{��nY���2REP3b��P�i�~�h���2�oxqòsRjPK� ����Q���q
��ا����$�
��9Q���qE���+^��w�_����W.�^�H��s�����;p�Ώ�L�!>e$]��n�#dWq��?�����6 rT=|�K�+6�ס�i�G$��'Y/1R���8�p��nuHs�Mݟ�08_}W��qn˙]F�#,ŏ�Ъ�h�bb�O�%�Ι�����l�x;Z	������$>�=�o���!)lH�����e�=a�����}��5�"F!�Ä�D���(����3�{���|xI�ݱ7
dc�cQ�@3�����I�@�����0�M�|��,����؆���sN�&+���:��� ������(�rޚ(쑭;�Hs�U5�,���2��Bu��:eolffVg�>����>h�,wF�ICgO��_O��W�\��jP�a�.h����L$���h�\	�U��[}�+P�r3�)LI����>`��D�R.kOwl]�n�h(K(��&��aʶ���4����G�5E����S[���kPo���r%c���z�pc�&6	�hD��=E�s��g�zķ��^>4\9w�!j,���.ts�x9��[[�N�j)�97�w=�e�Q�jK�Π� ���Vҩ3*�!B��$k��[�����H�o����Z��WPo{�� �ߕ�z!������;��f.���jqش�ʞ��t`��� �԰�B�f:N��#�t�Ic<���ZJ�h������ U�U�ΦIb����=]�@�G��J��7��}J%���k��c?�����C�1�8��/�ʞ�$n�t-<�{���5���wn�VἷB�)��RҊ�WX�	�2� 5}�OT�IT�`�zX�p>]���H3��;�,�d��fVٟ�Z-��ʜL$����ǔ%m���~��6��j��V�� :�e����u=涚�,B� �e<\J��*���5�����ָ���\d^�-�j2��H��G�"��~��y��S[e`�v�B�^��Lx�az)�����`��������:5��nq��a�� �͙�*��`�@�!�J9ψ;��7��3d)��cw1��������*�M[f,5�3�:&�y�s���*����m(`<�s6翂���R8�ޝg��t�����T��<"��P�S>��ٓ��b�S\�'� �;G$� �H�~v�Vk���"��α��1>At?����C��1_@I-��']��ja����ۻ@���C>'U��9O�p�&]�_*\xJg���
9���M:.|*��G �^�����-�����L2zF�[:�}�Y-!}�qq��x�?�u�(�fP�5�?v�D��M4/<hq�~"�Zq���� 	�,J���_O��Y�>�����P� A������G0B�����r�x�7�A�j��QJ]��2̤J�k���#y��q\T#���g��{�i@_�y�#H�YZ!Ĺf�/Fs�"�(9�D��VQΈ�����݋^ҩ(F�۳�^���[?N��_����Bk#ic��� �x���k�\������ݘ����+��^A}�z���3��خ]��i��ʚ5�Ol-�_�9{%<~&��'���<�$ETv���j��A�O���{�DP}��S4bm��AeW<�%V�O�Uc�3vS{��?н�	fwH�:�T0����xo�����2a�����z�Z��y:g$�s�Q�����h��BI�r#~�WJ2D�Pl�]�l�����
���Z2\�wM9Z�ԤԒ^��#�瓿����U�y��ӻ�_X��Gs]#:���*L��`dbd����.�"A��R��#�6'��;e���y��ck�F��uW�``�;��	U5-��h��\qMGs�V�:jy79�jAՐ�C2<�%4�֠*����L1y5�XJϻ9�k��6/7��\��n����P�i��	*�b����H�4@G�;<` ��?+&ÑZ�s�d�`^�'��z�7�9�Sw�îG�n��!�+���U�`R�G�jI	��,D��~�Xa�#�}�*�:��`�z�vzGR����a�[��s �I��ݪ�BhV�v8L�| �}0]E'548*d旁�M�E����i����q �7�`(���:޹�QyXO"l�8FS���"F̜�X2�'����Y.�	 �����0�c }�n�gg�a���{[�{黑�Qe�w��ی	k�H,l�&�H@�AD�"{q�`l�
����~��f̂K_@���`�,��K}����p�aa��Ӌ�[Ls���)�Rvh�B4����aʀ�q#�#��4d;E`-N�DU�MTc���tCU��r �������oY�b�{WEN�����H��y��1�g�����Ֆ��.8�҃ �b�`��ʭ
xit���&O����6N�1�;����o��ij��C"�W	�!�{p��������M\H�h{�Q
KRD��w2��eoq���!�N���ǁ77�N�7��dNx?0��(V���/��o���c�V'��#N�_���a��a�d ��N��fx��_c�{���+GM�M)��	��	���%p)��/:�
l��m�S����$��1�7�M�^�IY�eaJ��9�7���%�`���7��c�迯'��(�BĒgO���:�)�k�D`^7��%r`��I��q�m�0k.���}�K�Lb7l��g�k�ۃ��X����5'q�=:P��)�<��}s�>F�4oŢ����<���֎ZL���S�J��Ù�#�f�GA�U{k���;��+�XE���@���	�F�DP�J����*�����e ;a�Iԟ/'\��jc��F�x�tʄ���z)#D�l�a�9���1Yq��d�2�d���X�K�K�@���%����KG��)��	������Ѧb9K7��pLw�<���maܖ��H��{d��K� �!�A�O�p���4n�E8|���ߘ/�
��K�ڑ�["Y�|��Z�˓e�<@T���]��~8ǫ��]��^M�A8��ZyG��8�<v��Awv�y[y�x��.��= �4EB�@����/k^x�4E��2������భ~3��[�؏��"Ki�ES��շ�^�̽ �>��p�h��-*ۍT9G�gz uFY}�i0�T�5u�Y��0��0�%���
�P���.Sy0�v��G1g��Ir��Y���.��b"�D���A�a"Xi��0��z�L�3x�QTr��	H9���R.���*�cƫ/t���]�ǽ}O���)O7ef���\���M�HS�!��h�j'��P�S�%�����~-h�	�j �!�X����K�9Ÿ��W�(����uy�����T�y��^�_&�в&�-�z���XN��~�N"3������|*�r��~+7��sa�#���&ؐ�)i\r�O3�a�#f��Dk;�h� ���E�c:�-U4�kp�����FK�V� ��|�����6��,@�_,�Ƹس v���	j,���HJ�|�$���P��|tӇ���i�h�x�l&`8O�Ii�v#i���L��ߚ$S�h���Rg:!z�9�|�V��gd��÷���Y��U�W*]�&�ɏv#��-�Q�"|&��|���R�{�4�,�3�R�xc{�O6,^��J�h��>��bd�ʕ���R�ݜ�Ry.c%�c���킟Ֆ�\L����y��>F��2���T�bأj�o8�}i-v9r���	,��G��#���=��7h�d��.���I�a���x��aE!W(�Dj]�K7����@
䁾ư�?��&u��;$M��1N��Y�%%�d,;F��*�׃Vw�ve�l���8�ol&���u���1�im��c�q�Z!���,�E���^�%\J�trtB�,ʱ饧��J�I�� �#�h. Bj@}<,4[����h��&�eF�$�E�I|�;�q�5N���@0-ux4�G8���Xs
{j�,��>~w-3�ɡ����W5��!�b���Ib]����˒ ��7�P�yTF�Hr���.�ؚG�Y�37�w�HJP��}@��9MZ��w�ycS\�FC�V+�l�E6����B�H~��N]�iaLp��<9��ax�}�鈐�ʁ,�}�0_��
6�A�(�zWK��?t��A{4z���y�S�,J��x3��\�?G2A�A�.D�w�m�Q���+=�>k��.$*B�lS��4Ol����!�VeW=����?�=�0i�'��ʊ����G��>RU���q����)y�M���SY��w��dl����Wl���ނ�T���v�Pj����T�C�~���V��W�#��N5�+Q�)���{ �
M�Q����������'�-�gnM�h㈷1ש�^��(�6=��hWt����,������n�;?ZSW1i	�e�
a��c.$��Ļ�"�&L3��2_fϴF �:#����:1A}�$��/�+pB�Ǖ�|�7@ф�!N���e�0Lp�npTd�џo���+Ӳc|#@��7�r/�떰Lz
#�D-e-�����T&ن�f��s�)*�C撍��o��7Z�;��i�Ѿ"'�m1"�fo��k�@M��}�t�t|�r��y����$����Y�t�\b�~�����%�0�k��HRb$E)�d�~-.��Q�>�mP3�S���3āe��QԽ(�M��H�J����vg�},����T���4�d�f���y�:�Q���jU��r�~�R���M�]pSC��~�f��h��E9Ҹ��I6Jk$7�?+W]�3�K�a^]���%C8.WH�R���Y�SI��z�2�O'\�'u�w��R�;�jT�,@�z�-�U@�[Dƅ2�.���/_*��ꠟsn0nM*�VJb�)�m�'�
uY�N�b���4�}���e	Aha'0�#��!��a�SŘ&O�|+�aH�	�L��:m;CkI����O���:�>͹�����/ʋ����9�j�T�#gXD�o�@��͘��-,��H�j�J�۶f�_�g:��o�s����O�u���n6������b ��ّ��c1�~���������.>%k�	��t�.f���½�d�Y+zzI����pX�+�b��CiI�s�	��D�������e�\�QB��YI#jM�� ��zo����<��\@l�Qmq?cM@oe�5�UP�����ۄ�H1(�؝!����*ސ���N�܇����R�ŉ���z^&�Z��
�R�o}��/��r\�����t�"���X��u�is�����i����8�g����Z�Y�gM�@?Y���b�O���Y-�_^��";i�E�Znh�T���X7qSb��.�CW�6�3�t�k0B���|c̵^$�P4����Sl���_-JP�a�@J����`��~[RR�@M�-BX��m�o�a�L\U��C���"<����k��}�����E��Vgj�2}E����dT�}�T7^�|9?�گ �י�����������|��w���������U4�q�*b����&w\�e6b^�� �k�̌'٬ �,�Fi��ꌢ�j摩V���0]#]Z�����;�^�>��!`�(bg�)�U�2�i��U�x��ч����Ԇ�/ �-��1�$u�f󺜟�;p)�%=wi�^��gJ�R,Y��y�d��h�'�m��fG�Ô���R�ğʴ�$yJ�p�Vl����Ec]迖� �SȱH2��0n�͞��E�٘K~U�8wYaԑ�x�_Fy�0�"j�cr�6��髌<'��{ܾ5���)Sk��~e8-?�%YP%��m��]�,	Ds�trh�,�pPw�eCs*�A[T\!tO����I��H���ME6���,��ڕ�Eu��Y �GM��m����`��҃|bӧL]���#�ɤ�OFm��@�_�G����R�A9d��}��+M�a_RUx�_H�a��ȏ$P�t�������8��_�{_��K�e[��.Ҟ�R��hآ�9�6���g����1_�"G�����	��3/X�
oX�GHgUc�O�6i �vn�I��	�C��YU�1�\��Gc#��O��I�ԩ� |Wy�ri�ø�U��Q��T�/������8c7��lh�	��GQ�nCx����֝�4��Um�v����D~N{[/�5�ua�L6�&8��xHA���1�R���a6��3ܰs���I��7!�M\��;	N��"/´��/�9�.̴�+u�`��N�*�ˡM���H'n��e�����y�5
��c�����=�{��=��9��
Z��>y�Ϸmz�Ŝ��-O� N;� H��烝c�)M�=k���;4Xƭ|�F���G���/ ���3P�T�O1��Ҩ�+=�ߙ�f� �7��ho<���Ћ���)�p��3 �^D��vIN�v4l��k�r�����<�\F�RG 5%B�|ܿɻ����b~u�HR�< �L���q�: 7�^ճ�<���4d�_��FR�N�):�-%��r�敯 �(�bx�P;>���LM�i��3$a���������1�����ݕ'�Jn�ql���y`���8��Q���a�k(<8޾� �J��x�� q1��%.�k�;F�`�����Ù�&k�#s�	���/]�������<�����w��$2��|�wa3�sLBp2����ɐ�W�g��n��h��9x	6'Ɲ��!�����a&�M��	�=�`@�:�|�Vs�I9TPvN)�� ���k�[�E�mr������<��`�n!g�`:����1PF�ّ(��G�Z��DX�;@�K�\( x#��%�.˜�ԙBl���+L���i5_�� ��C>�c���ɵ�@�1��ݓ�T @(7��߫G�aB��@;��M6�y�Nk�jn�?�+�	D�Mn3�O�=`Reګ�f�#�����S��?�>���z	������$2���Zc�ϻ��jGG
�G�}2<�{v�͙��#�G�Kǭ���<6v�AX\��)�SFJ�*֤à��4Ɍ�w]~�q���V���3�2�EL�b�g�V�ϯN�e*���Q�Sk�Mk)��h,��0O��L��~���m)!��w;�^"ͬX?�����A�w��������zP8GbVj�D�VS�1Sq�O��٤01dIr��h�͌B�u�8�D���4�� �ݺ5W9;��Q�5�_ħ��]NL��̙
0�JI����]��g�<��%d����j�'O��N4A]2-����i��)y��M�{���}�!S��p���)r� �0�ZYy9r��s�����R�����C�!te,7+m�������N~ ��Z�Ǹ㔕J�Ѿ�ޘ��$��J{g���Ds����ƓO҇]j]0�?8Yv�r+�6;0��$�O>5g���L����w �DF��8��1v�Pv���������8L��7k�ͣz.������z1(�l��f����n���g�t��SE-�b�17^!@W����L�����Lj�������cy�.���6��6s<�;�m�{���O̮4�)��x����Υ�X������pC
W\ݝ�!�=�[�D�ѹe�b�c���[n}������		3�yK�L]C-�'Zv}��������e��� �_g���l�ePV���K�5�Ғk�mxW�gtw(�%LַEԕV廥���J3�+�\�Ӝ��<�G��̮����֏z󶖍�@����;��=o�i�����l��#��2Ui�=dڹO��NX#��`&K���̈u��[6��R��}����%�CC�Ʈ��&���]���s��A�������)�b�l��j��"�g�O��?�b�^{�p��M�q�2:C�s�������{r6�U�O9�'-;м�k����*LD��_�:�7h�Ok�fn�L����X�_w�nb]���j�ӏ`0�����<4��)xD�g�M�^����W��6��}���g[�|+����3�0[�o�HM�<Ju�Vs�`��xW$�yM�D=�Q8���*P]~x��##]	F���~d^i����gd���%p�O�Zɪ�SK�qn���2��'ww9 ".�g��rZo�5�����1�үǊ��!�e��(�E�t�q�\���U�����D
I@���?;���^i.�$a��U�ce�p;_7i�W2������f��>z���#*ĵ_ߥ{D����m�Ze��kvo��@�*��v:u-�2��='�KG���7f��*��d�Q� ��D@�C?�].����q�|&��$��+�ʂOM5��:�����y��P�H���r���2~��S�'�K� `��:����%��z���i�u�b:��V��G@>�����
������LFq��F�	�V�;oH(���g�V�m�{;=�cG�����#M;�oˣ��&��� 3?�L�H��~ԢgV�w��_�f��%Kv�]Qs1�;Y�g����fò��ݷOx7m�+���a�k�Ou�|V��|
A@�aC�T�
U8���n���(Ý�S�"�44|���	�bg�@�U�B���ź�=MҿL����#sv뎽��J�3��E;3�6�,�������[�Î^�H �����x��A�g]<�p
�@��|��X#�\)aZɽG�[�^)�&6@�~^3]M5�B!_l�2~���
�췃>�<(�xH4�������� :�t�l�\A�DN ��|o+�:p"�~��:z��bU�r�j�7k�:n?m9��k�ƞ��א�N�YH��ITv�{�OR5ow�)�D��}R
]͏�_��4;�qk�V��S��VT�v�`��/1:��*_�b�e��?a��-�[���YŇs�[E�'m��3�D�ZUt�3�=���n~��Ѕ����N�D��3������׋00.޿˖ڱ����y7MM퉣/w���'0�v�t��F ��D
fkh),K9F���7n#�6����C���j�@8'mB6Iq��#��v0�l��g�^ۈ�ޑj��D>g�`²L��]�O��W��i��GKwjLz}�	�r*�y��5(�E��s4��gr���G�3�H]1jǵ��~8���m�Ʉ�q7�������8�AubL?�'�/���9S����W���$��^S��Z��,_�q4��|ic���.�]��[�	�~���U�����_h�DnO��/N��i�kkϓ�Ƞ7&�u�ҡ��k�j�����8��r�QsVv�4���.����	������$@��oޒ.���1e�˥��A�Z��\%��s��|���HV���X�a��s�f�L:���U��;��0;�` ��4�Kr*���[�����t�U@�<7�?��v`\Z��n%WX:�@�u.��J��6a������p?b �%%w$�b�w��jfU+�d�*�b�������`���+]�j�PJ��G�Mc}���(�����>ν���jͫ���V��W�푘�1[�Zǭ�bv�%U&_d��J�0. �-�C��`�h���<Ye����'�+�V���fl�ݖ�:�#G�F�}/Y���!n�A�b��7M��o���c�cܓ�qC�P�\���tFS�d0����R��f�K����J���{%��Τp�9wF[��{;z괱���*��.��Jq�{^:s�u�l��T����t�V M�2�FYqC�t��c˯봑
���5��Q�Wq��tÄ:����@����r����b���CL�z�B��k��,�G����Y��N��z@�y�c)�Th,8��R�����0U����:�{x����Ex��~�5�/|P~��S܎<�ܦ�DZWq�VfCTȫ�6Ur`u�QؽB�O�����/Z��K��*��%��Y�K^�5���!�a+�eC�_c��u߹�W��d_�sF���L��U%���$�0{˱ZVmU'�}���<m#��ډȗ�aG�d�+ˢ�<)U^a�1����@�76a�:�+��S��5a�J2"d��V�*G*�]��X�0��A��O>�չ �5xQ$�4�k��E��/37�,4��6����S�|��U�q��� �]!B*7s+��&vϏ?�z7��#aeM��G)�p"Sw���tf�)�޹��n�����Q� �a�jd���!�/�Q�t4�(�
%�R=�-ĩ��@�О�-�k�hw@T�����Ҝ����r�e*!>[��8���=��/��)j6���z�_�C�&�!Z�:�6x��lGD���Il�D({	�/�
RȲ�>FS-�d���m�ι�' �(1>{.t!5��,�aI�ƈѪ��mu)�G��n]o��zb�ڄZ�J��=�z61���nn-���7�N��] ��U_�-zK����Q��<e�U�|��v�i��})"�-ݬ��"l,�*�m5E|��^�����q�T��G�6��d�Q�E�PE�����f����,��S��u�G�Fx�8��jX�A"��֌��W�8�0�-\��+��W�����g������O�w��qi͇�����Ҏ-���&��;�7�O|��L����*4л`�������#�x��}l;�8|A����*�.�m� �#��>��EB�Wݿ���}N�rAL���QM�A���V��S� G�*���!y�Ⱦ3q�уĵ���;a˃���ݱV����ϋ�8�� "���R'`���7�K�ȓ�=�2s#��8#H�?�����pW�%7����o�)x9�FcCD*�pc}4-��7����-?����G��;'�B���/Ƚ%��������<���})6|���)F3N����j�p0��ӛ�	s�1|G!��%��@��c~R(�b�zj��v6�1W�|��0��U��&���g���7���wK�]�~Re_4,���Ί����5I�_�� ��G��蠋��B��H���_�U�M���J�R�|U���������w����N��|��m��Z�\[1�E?��N� PC���7�pGd�*=����P�XJR����ɭ������@���� >�b��9�G7+ѰZLͷЉ�7������r(S�.���\��%������>�����h �<����Cș]
?��F�&1s\@��-R�.��&�e���Gp	J�Iȿ8C�K�?�/)���KĆ3��w���l9K�y��d�'oW����)�yg� �E�{���b�3q%I��i~��6��~�EX���Т��{�
EK�����,�A���5��zZdlр��%Q<�k%`S;�6��j��`}�*�Gn��z�ƈ�ݪ����2�mA�,�GJ7�!�5�ڦ`���ک�AP�ثϔ��-���&����.��)	��5�->� �m�A�H�.q
G<ۑ��z@���(��ee�oN�Aðܞ��ά��]��"���H�=2��ꓚ|�g�-���T�@��<���t0�#n�O���_ğ*X��Bf���]o���)�6�yU��
�э.��F����(���P<�����SC9I�y�`�F�`���eAF�XsFV��{��Q*� &+v[C��廩�����г3��X��$	٘k�f��q�S�Nh(������C9B w��E�m*�%�+�;����Mp�)��_�&Pz���3��8���f�'V>�!rw=�V\ G�b"YY��C�����Xi�!�G{�þ�u�� �NF���e��r⹖Η�:�rIN�"*�2��F���j�}K�v��DY�/��k]����U�8wO���g�W����X��6�R��i���$�!=~�,��]후�ʹo�>��apw��\�b�b�)ԃ"qt7ӼQ�Lc-�s�g,���+��H�3���Y�9�����%���8dp���Q=6�M*�iǟ�?�X����˷	�F��q}ӲS�G����%�$=rD@�ȏ�;�
$&�9�5��ͷ6��	2�߉}�%d�[G�����;��| ������Oˡ�;�i�������ZZ�~4c��NQ �HQ�Lx��Ź0����b�%�����l�°�O1`�}���L�H�Ų�*�C���P�z,��˒�6儊�I0�̶����'�q�"��Ȫj�Ě��]z�#�k"�ƃ��׏���� z�"�L%��ә�Pu�l6��(�h�h�xLr�6�)B�>J�S���_�ȊA��`��]�s8�y�[|����|@Un٢x$hο`�uqy�}�|u�i[W4���J��-�W)($h�`�½����?{��E|j4�a�z �]a�G3H���^�M]"��6��-�:�)|f���{�3�P+tE8�}�<K��dyq�����������o"D�*��`�r�	����M�o��c3�\^��.i�=Q���#��̓?�i�I-��?iznV�����w�	8l�K������a��L�|Ъ��ɨ����(߽��Mh�?�7�heu�G@>� ���CeQަċ^ �ֻ�Z��V������Fu�� m�sI�$�3����n�u�in�Y=���dбjS��ǟ�O�0�a��)�c�(������_.�<k�0z�~z�~���};�7�	�x;2h�N�s�1:�N9�Fb�a�ƉpJS2�z�X=ņ�-�Qמ�x���6v�\�L�(��{�?I׿_@��=E����p�f�vM�#I��H~�Q��RxqC�7�7��4'؆؇�ﰗ@��� ~9�G5�]�i�H_z�;h�h���XL��O�s�h�\�o�<˩�|������CzM��˔Ǜ����)���~g�kx��6(��dCz?�j�g~��^���v��^b�;��>��#��F�Y�-/h	��3����23$� H�{u�@�m���'x��.ņ���a�5R1h���d�<V(�^Q��-qʉ�����ܼV���I\x����iF@8��zƂ�a�\�V)���-�?����ow�q��֢����� �����|m"v���d�&zk��<7�!�Q���+-����2�*��� A�� ��3��j��j�j!�yMU�l�v@N�� xݝѢ�h/'�v�G6�k�M��������ջ�jʏ��4%�x1�A �
1���R7��G4�.A������{��K�	^�n_r�JL)������i�xB�0 ��VF�x���)O*��!%�D	G�8�稁r5�t�S�tʝ��|/��5�3:��/��s��d'�n8(���P/�YҨE6c��(�'�C��Zm�y������2E/�9\�6V�.#E�7�[LF�A|ʻ5O��R*�U���{_�$]Q��=�RlT�P�y鷾�yn���'������2n
��ԗ�TU�Y�iv���S?<��[6���aAt����?6?�Z�7I�)O���f�!���P�Ԗ׿M��I>��*�ps�� Ι�[��G#���(�MB���_r(������2��	�qe�d�r�$����3��(=Q1�i���OU	�ܑ��E����7Idr��^/Cj��|��>�Rd�"��"ƚ���5�3�{O�M��۲�5������e��6 �����k�a�!��5X\��Z�b��,�?k"��+�������m���*��f�/ �⑋C�{."���׶><�ߕCC�<�DJ5�en�%S��f� �7�OP�	P��fIZ=�}s����]by�N�z��T��q����4A1G��N��^!%C��V�w���'4*�ZIS�O�k˞TT�/��<�	ǿ���;s0�o76��
�\8��թ��=.�-\B`摊L�ӎ�f����-����۟5�#�O" \s��?<��%�vE=6)7D�[a�_������l�b8�aȇ�p`&��/	;q�<}�M�7=�vh��LP���x&�@�}����q��$$uc]91	����g郬����Ț<���bQ��F����iԄ�h�9xL��)[neC1w�䢼^x��T�~K�c� �NyTU K��O�E� �Hx��y
v[Q�O/�`]�+��d�C��	*�]�S�i�v�t�3>��~YJ�1J	0��X���"�F��ڑ�L|�gT�Ѣy�I��&mU�	�"a����0��G���w��=��"�M����E�/+��Z�"�W���A�E�6tz�?[�5�������T=܄Fb�0K3|�����0��<kIW7tI����<�[;���J^��+�✨���)���gE`5K_L�]�w������ֿ��z<���	������We�I�LF�h��T2�-6I7o�������E�h�ǻ�o�j�m��|��
���G�/"���eg� �3��g8�ƥ�J�5L�o2tm�ۥ�Ȋ��u4߷������H��SP[#�9gR`�3�	~�4�O��-�l�*.����\qJGYbjt��[�rhW�����T����⾩{20�v�k���a�O49�a�h�=��-�	xak��wT�h�` �Bk?�Q?é]�6�^���(	X������ڒA�Yz�_% ���Y� �WH%lZ`�~��ץ�Ӕ4��l���U����}�Y�}��c`�|����a���6S����O4�w�G!d#�M�|"��Ff#l�\8��R�,��W��~��D��/�`Νе�6or��4��k�;�]ѥ��ND;q�ڭ#�������� ���}�JāQ��RqO�ߊ��(�'1�%U�7_�-��0�#�}���o��i<�M�B�TfEqg�Jq��e�
�=���>�tW輟�btf�M{I J
kLb����c���H7�m�å�ý����,�V���f�"�<S��e窬|Q�1(\��W���fZW	'�B�$of�}W�S�g�����lm�8~�4�q�k��z{Pݐ�8 ������"��3�9Y��t8��h5+K��2���@����GyN'֋�V��Ǭ1��]j��V@�������+c��)��5oՊ5���@ˀ3Dm�:h ű0ի7�Γ�i/i5�D,.1!.K>�A=s-Un�b��@������� <7����ET\P|Omy*�֍9��?&Y���YG:jh���5�(�}n�a�DM�S��EB�{�K�SWbKW��	Lcq���>��>ѷ�۪ؗ��0��������,l�nB�`�>p��pbX�p��?m��s=��5�e�I9������VsuZ��!`B�D��u�U�T�����D�Rto�`�UV����̚�T:� �(����^�W�4�O��{��c�0�D��7#y��2�Q�T����V:jR;&�$�|jY�sx˱�/���8�e��� xpY�4'3�͓��.G��*�-'���FYج0F9"yb7d���^Kc<�'�v�d4Q�۶ ��d�"=@W��O�6�(�'Ae�G�e���[�Gm���.E��Ml�\i=yFh9R�����6��b�d�!k1TL ��j�u)�݉��0bOM�ȧ���6?��g���qiV�x�T9"*m]]�U^�=�L�s�=R��h�@$CK�ѓ҈1��~���'<=��y����Ca,�S_TK �E�
�������+�ͫˑH�<��l�6�KH0�����?b�,jn;u�ǎ��s��#��h�e!b�Q�sie���W��E�.�S���;��B�^tza-�{�,�}���5�!B���g�3��8�B{���G�5!>U���n�de��\�6E��M�V�� Y>�I�{39F�5Ʉ8�٢��L�Q���<��bG������/�m0�S?��f�@Y��?�R��Ctm��[>0�/d���-�>����i���%�T���J1��=�+����~���̢���P�y�3���'��4pa敳��T�"�\�mRnqC^�p�/g.A��k#�"�V�j4³�����_�d&��@a��L�����M��,;��f���jNN������
��������Xܜ��C���C���xe:��|���ugx��`�%W�>)h��-ϥx߳����a3�!كL\c�G��\���v|�=�)�bI\o��_y�:���wȠ�_)f�,{P�d��x��), /~�0�0{�H����{�y�
�13���v���s�́q�{��j�� 텙E�k�ۍ�[/�t1���NMK�-io�1n��Ѐ�R�}��"������!��⋺��'�m���&����K�P�g��؝���h95�	j����E�d5�P>0!S��+�-iD�$��#G�O�n1��$�nG_�s�g��i�6�1�ԡ~���!.w|���d����(&�j<��+ټ��I��"��Ŭ��Һ���~Hhm T�`[��t� a:8�rb�M��w]B<���E/�ܭ������h߱�"�-r��?�ӡٰdd2wa_�mA��j�e�]��<Ȉ2�C<��Z��!i�����~��[q��@�diqM'��t��%5����*��9?h�k�4&*����H�9�	Y���סD��f_�/w�6$(]]��%L�����V��2��U�n�s�Rv��~H�L�T�~�o�C����{ �g�����a�Y|�9���&<�3O�:�V5��$�kn��j��O�jke[�`���SQ`	(��A�s�4���7S��0o�������`.6�ѷp��Q@��Y�VӤE���=���Z�(�7$^��͝0vg�u��+e�1b����R?<��,��?z(XfH�p�x ��tƔ_���	y۞I ��t�ҍ�H)��۞&i�?���9_;��y	_F[�G���ڲN�#Ps�'ӭ�b����hP�Ks;6���Y�|�L$�m-�f��Ս��R����eWC�۷�D(у��@�PA�
Ş玶��z��S7���2��7(0t�����L��j{|)k��+5��6%<���F�]�	@��^?tz�`�֎����5{�?��~�q�}���WMj�Ռ���m��c4&"��C�� �C���1!��J5�~o��T?.Ԛs��R�ON�8��ӈ�L���h�ۀj���^� �\Gڔ���9����s���{�������
�o���^��@ge����e��2:���uO��e��22����,)�8�VD��A��#�{ޖ¤&��+�B.'��!:QD�� �y���*���6/���
:@�P��p��J�𡅾 >���K2�ɣ�-�R�s����)�����[鳖%	���
`*��q��<�Q� �ia�KA�,��Z�D��N�I�`:�;����αX�K�����}�c(�P�ؠ��]r����xxOAc�ѢT�\<ѕ�H�T6������D٭���0
�`5����]�|��9��5$�p���R&3��>���$3�=�t_� |(0����1H):��U}]g@�/)˔�擲X��~8/�m�Vq`r��/08�'"Jw��6�S[тQӬ���Ż�������q���/U��kt��s������5n�d�K��_/��9��l=���ܣ����	�����������4l��iJ���Z�?�!@�h��Ct���ڙ�iX���9I��m^#Q�m���$��$�V���qN\�_w�߰�Hn{i�0O����&2Wz���`��
yBPn���t"N0eʼ w�X����q��|A?>�x�%�"��d�h���r<+w��$�5�7t>3$��*\�)����r�l�#�jC�T���7a�g�)qe��S�'�}�Fȓh�U�tu���\�����|�,M�c}�O�����H�� o��<w��v59g0������lԖ�P_$�S�_E���&���4��y��Kǫ�"G�-2$B���
�ɔ�L����S�6�ۺ덊&"�=�ՈĨE�5
�A��m�L�>�D�+(;��v�n�R�+���H_qІh��W����.%��A}�u�� O�Z�#��l�K�y�-C���A�Ќ6�7/�����&s�zhU.�k@+�俵`\&Ȁ���pz�s�L9�C��E��9u{D��
}��+��.�%e���m��ljZ	��G3�������R�>I�c&2*�]��`q&��{qe1����"���!F�K`q�0/(Sа%+�Skw��*�~*JL�+� �������$�@��@V-�h2l�+�F^�坦rT7i9,~�=��p�u
�&豀i��jM�xb-yY{Y҃f�b��>�7��d��a=�=�&�,����=�5��Pm�)�U�u����Nz�5�	����h�3f��|l�f��o���P��xo����: X��5!30$�e�L{���N���u�8 2X��[��1A<���� �c���LX�c�/�Οߐ��|:�
<(�pvrMB�-\�K��DO�sy<�����h�YV�7=�p���!��5���_�
$�eƣ�cK��aK���EY���r���:5�P.�k�B�7hˈ��u��SF3\�1�Z��oѤ��!~�q���`�����]1	 ǨG�qӽ}�����w�ݙj�'�}D^�9�9S��,�u5"��U%�|�I�b��j���V}�ۓY�O@�ƽ-F��GI����_�V8�Ź��m�A�`o��z����^b*���6?$�����bdc�����g��0د�#�T&��C1_����:�����[x륚j��gn9��:hOXf�ټ:�1��&v[#�綉E�r>�?�k��+'�?7r�Ί��s���4�h�����5X?�ܧ\p@�#.�,,k&�E�H����Sa���e��5�D�9����$�}Iw�8R�aR_4$��I:���7�Jste�C;��2EP��D�!�x�al���DT���!`����-��+�p�/뿔�]�Eݖ��P�[k��$y���+*M)��P�D�V�g�XA�"��pcS;�B��wF��j\|��-G�d��`��ȗ�A�%(��j��QW�*X��<\�l3���U��]z�4���ŧ�$����l;3��X8�$�J岝���O��.�9�4���H �mX�?�z0��ʟF�|�Os�5��o@d�a݉�t_�ޖ��,5�ϣ$��S?@�N�FD*���p ���Y���@�'�4��ӳ᳆n�s+�#r�ՇЕC2��%�n��]�� ���f��*�+:�@��� J�.�B�޻�&��jr�Sf�*��P�fXQG����쵟ß
�{>���D�OŮ+mlY�bP8������:���� �� ��*�uWÕT�*���mk,���.v'���t�ޔvA�Vѯ�hC�d/�䵬?�k��1�k�=E��W�RJ�#�Q<����gZ�>�u�eڒ�K�%[�.4(�	�v�R%�Ȯ>�^_�N�RZ�����y�1s��i�~�=�]åȘ�fx���~�.�����q��Bڡ��'���W��W��h�d0`�~�q���VN�U�L+�D�a�$#���i���n���r�/�R�,݅=��.{~��K{!�s�r�����>�t��͉�F�	/��\�׻�i��(�N����u�Qg!���J�ZK��sV�Ƶٻ�E`�x�!?�w��b$b0�;��z�y3�4GmX�+vP��ẉ8����#�|��}n���`/}����p�</���<Dcv"��{�O�����y�,C���b^��c�b�$隉�K��q�Tpȷ���.��k��Sp�@�ֵ�Y���,)�t�ܕv�$��DzEg1|p��u���~3����!qO�)����
�.���Z��N���V_��&-��sEU8!e�@�&17��w3���E�4�H�ú�$�E�vT�R���\��lW���*|f���,�k%���^��L�S�n�I���_M�bނ��ފ��	��9iR<�TQg(����f����P@Eu��F�Ȟ��A�,�=<����ծ�it�WC3�%��]�#��(�#G���ƌ���� anM�� |�@��A�)�:�h��ˍ�Y>�r�#�t[I�K�`5���'��Uq����@d3�:�
"~����]�®���2v��<��C��G/�4��ҀTi�-E�Җ;�����2'��kh��hB2����9k�+/bm���*��2�	`C�'HA�9�0nm곕&���n���_׎h4&%�A��MYs���˴)L��Do
"�����ս�?�\&\~f%QK]��_�x�Z�`��;V�k�b"�����&�xK˽�=��T��
�*��m�Zm�"G5����Ō:��0'�'�;}ع�a�S(?c@�zI��܏9�[L[	N >���/`�e���������r;m�:5���A	نa�ʑo�3��v|��M�?Ԍ&$���7�V�ຘ��l[��u�K�G+qX���'�(����m����2*Ͽ�h#���8l��s�f]��H���2�I%����}%�ٗ�����'0��,Bß\n�/g+��ƀ/yq&}��� ��LO"��x,$������U��?�BɤL�͙�~�@[h(�.�b^V+��v1�s���Py`a>f$������`HXJ����~��6���8���,��D�bF�'b�P�4�$��#�թE�v�X�B� ���#è6��\g5��C<#�Ѱrb�w��x�����U�O(�
2zw&QS'E��8("���L?e^��Y�e��	�(2>���@Ea��o/�gk3��ƈctF�<)���gU&B�k^@/8+�OJ�+#�m`�oe���7q���-ԂA0{D���Ys��)/��*��C�^u�'�	$k�8
R��(L���,t��7����6�KU�)�+�s���X�/��u�7�����cm4,�^	&�6?8�C�M�;�@�l:*��S�+��i�lS��lb��ժ��0���zɫ���L�1L���o#B'��[��P�^f?h�.�C����<%e�nhB:��]�� ���M6�UpV������k�R�Z�[~�L�q�퀸�X�Ae* ��Ǟ�K�ņZ�2Z�V�oBDI�f\X�	�'��{�W� r+c��X����_ 	�������Lq�������Ͽd4F��ߠ>��j^2������)�ǒbm?)Hp��#ʽH�A��W�g:eOs�OF�_2>w?��^��f�Z�@�Y�4��"2dB��d�@�ue�t���"�  �%s$���]q�8�\�E[�c+��u��h�О����`mes�+pA�����K�`y�"~��p-]_[��,m�����^p�ڴ�5(T�^��P���� 2���K����E�S��X�M4�3�ӚN@^&(3߶�{�/�@ɒ�'0g�5�.���H��Rl�Clq���*�o���F����{�I�o��j���,���?�{7
E�����^SϴKYqr&���+־D.IV#!������n>�����Kڏ�D �W��6�.D��k� 3kTL�@���=��͊?�f��U�K=��V5�ɱ˷Xp�f8�`�yX9��&�&~�st�0rsudM��|��H|z�O����\��6z���&-T�{��q�}��(�eGV�/>>?��o��r�۵�Q�fS`"_~,�y:H�$7c�i����$��L"Ić�_�JVI�-�����F�eE��i7�����2k��,Ӟ����:�����o~ �MMR�1� )aw�O�8Pr�{��d�jmO��9�C���HlB*3ދۡҡY�=>��k��dF��bl��)2�X�#��\�b�|���X`�|\Զ�~��=~NԻą|�O'����I��������~�`�<ע4���a`'���	(Cr�gP�v��l��9�`�7X����v;��hq�8��cK[�>W�6�I�@�5�;!Xc!ᘔ4�U��MS��x��"�,EǊXΉ�r ��CL�d%@ZH�����,[�J~e��;���KlL��k�j
"�U�O+R&^�Ƃ�No���D:�������i���&O�+��E4fsD�C��4�����ӏ�A��Sn�����:����q!��@=�G��#G�17��W�w�U��^[H��|��bzsjh� ���i�l Űݧ7�?����������֑9�BȆ��ꋴK�G�t�s�DQJ3�lsx�yc���y�8�m-�\������J^ǛWoK������W������4Ϊ�R�J?�/��7&�����g�B'djtu��AI7�i֛�C=ʝ���G�)��.~���Ս�/`��9�F%H;�f�\P%�"wH�aoS��dMk�'�TY̋-�Y7�*��d����Lq�bG`e9�#?���}8<UEG���6���?�Z�e��B��.���z��0_��q��aL�S�T�����ʉoتe�� >�� �^��[�������GE�F3�d?ѭ��hZ���N��Z��N�q	�p[��e���n�ؕ\�G2�8b�+�$$�B�'�,?��9�/�����P�伊	P�iY:p	�VZ� ��R����b:��)&^`���j�j�i:~��!kk��W��r.j�|��S�ň�,�~���*�3�WfY5�0��79��UC��ո*E��1���FQ��ʓN�P���(�S�.��~�����:"Ś�jBE}��0�H$�rz�u�xε�-1[TI5:#G�^�y]C�b��W9m�Q�!a��f�>n]��p�{�$��xA�T�9P���%K�KGB-�'$�0���ӟΩ���Ͽ�SX`�U?q+2�6���ى�3�
�=���PhV{�ˆ��ڔ�Q��x�@���J�6 �8�KrP�h����!�p����,��;|`�߸�}^ܻ�aFiB4��)MNatȚ;�:`����K4;?J��Z�C�\�:�9�@:�	�(d�S�9s]�Zھ�
�͗I��g�������M�y�(^=y�b�,)�K�Dmք���S�8o}:�&������w�Ag��n�Ա5$9�}��dΚ�q9�����Q�P<�#�Qv�mha�)cr�4��Lwi����8�K���x��6`�	�P���'�w�.��m��2u�C��^��߅�s�ݗ��/�2�w�+���yf��MB�r�KU�y��©�G�$�X�\XGҖ�@
�#*Lr}j=׷��dTV��c�P �AO�D��t˘b.�Eo�T�riZ��8I�j_!���Y�}�}Ȝr����p3��<��3��_�E��!���]�����:�L���%Y��p������&>��Q"v��o�Lgu����,�e����9ct�y�Dm��% @�ݻo�'SnRK�Qh�s '4�傰�-�� ���>�q^���������G���6��3a��9o֡	�)d��E+��P��t\���n��[��F~�3.G8��]�O]���P	��l@~�Z��-��Ņy�䃜$�=�0�~�n; f}���0_���G�3�h	�J�m�%�c"�Ĉ�~���n2&f.2�Z���w�)�Z(OVJ	���9��/�6���epw���KQq$FM��}NzT��^ň��D���4TFa��|������E(.���a��C��X�G�Z�H��B�ܢ�� ^ǐ���K����FB�\i�<
_F�t�0Ԫ�R�1�?�t���٩8	��!�dE��n��ʆK?s�x��u���fJYç4W�P�SN�H�_�94J��k�kC�R(`P0�Bd�`���X7��3�^��'��g|%,Y���=��܀+2�&��<6G�{�'� q�N&�B�3�8�����9���;�%"�e/�K�Wl.]-��l��T�b�����'�t6!�y=����n���^�+V�2��^%�-�O8 6e	7��6hoW���֢A$��=Ԉ���~���S�9q}�5	���o$�H�-u@Ce�斫	�j�\��~�W�Un���������u��33�ޫر�9v������#�%�T�>�˻�M~����(���7+�`�Cxz�fo�c����Y�HD%����af�i�4--?E~u���ZE�S�+2��x���#��9�C��^s�����c�5�o�xhO�oZ�.�����{X���y-����#��׾
�v�Wx�#����d�� #�1O2x�;��	�ˑ�O��:f?���<h(׶�?_Z]�^���U�L��X`�<I��wg'Pܶ!wO���g������@�-"��{O	�^J�K=D]���x.oY,�����?hs��~P7�Ym=%�f���0).�#�T�KPE��DM�|�6s)��s����R�/r]�s�����a�IJ7�|a�ֽV�ޕ�+p$V�����l~ ��*{�n^p@�<<��#�;D���?O�����^�5�T��)$I|(�C��V��~�K[����xY\�//�%�(��40�dM3����c_��ۍcyP}itU�-#p7�OԞH���#lA�N���j0ՠ(��	�k��� �׻�hR���*�I�{_�f��1��K il�Ω1o��p�A�ae�zúv�w�LB�~$M9T5�}#΢����?�����J��Ôs	�uG���s����6Յɣ�O�ݰnc��`zQb����kӏ�B�^v�zV�B�;q�6ֽǝ��'WnoI�*\�wA�_B"��.a��T<kxmz���+B��'�?���M����+�+�x`�a��Hc'�=�A�����_)7y����11B_57����b_�)��p�U��nB3ڌ\S쑦��h�����H����)��-�ε
v,PWX�E)sd�@��NP̓���5X� ��/OWQZ��d�7�LIƇ����!���n���PGʐ	12��<�ε�,sن��`��F�~;@4�D~J�V<q�!_(r�x�X�S�7Ro��s�pw�k��n�ū�t�I�����}[?9!T5'�LnhO�l�}ם��w�2��J�v�ݤs��Q��&|��Td��B�|�� m~S+�	�U*F<��B���^��ʛ�􆚧���]�UgBXq��-@���q����/����&�R(�~���$O�W<_+F�`Ro+��H�U_⭧(�P�=|�ۓg�	D�e~_����/����B�|7�-�<B��Mh3���yg{��j�ٰI�DB�0�w��ē�(���#&��֍�Ob!9ha���VwP<�P~4���̋z��"��Z��f��p'�U����	*f�Vy�X�0!<vҊh��i>s���T7���b��w%�Z՜�^��/���=}�,a*�%T`���Mԋ��)�r�r�S-�j�^XX��:�r_s^&����|�y�g�
h���6���0�=cR��%���#��C��<��x�z�}X����\��TW�T���킰nls�N���)Y Wz��c�pF���� ��f"���ϴ���&��I��ga�V.��f0�)Ԋ8\��6�����靸���<�|�N��M����f�����)��KQGz��s�y�d	�=DK�N�@�����!�D���q�}x ���1�T�5��n_Uٔr��J� �j�ͮ)e��lx}�x�﷯����R&�!w~��AUL��K���bU�+��(��Gz�2�S^�b��of.���H1�=є�,��ݼt�����a&����#�*�ơ��Nㇼ�^��닢�~*��MM�\\,1O�~����IJ�C�E�b��d����sY9Ҙ`�y���J.7M|>��f����q&�5������a	lTޖ	6JD�V~�AA�
$�ag^�ɑ;R��웤��L��T���4�W!���g�nx~DvI+ֹ&?�E`1�a��&Ey�.��cc%	L��bo6���|�<WL��B�&��U����է� �l����>�~��R�9��M�s�"�����&]GtX~��7n����4�Ƀ�YI�~Uu44;���1��y��	�7��A����(�խ|�]���e%Y*��K�ڽ�}�k3G�޴�����
�.��*'���VAA���.HB6*�d+�r����l;�*�bZ�'�x��D�4tyr�	b���}E��@���q�j�OM��s����lEC�ˬXkf��xt+�{p�dω%#e,N���'�3�_S.�����g�V�"
�Ż���R�����J��'��EOtv�3��򈵫C�u���#�Ac+�ʽN�����5뫈V��,O�����Qc!T�O�H6�uYW2Q����I��`c޽a�\�_L�(g@���6�g�E�x�����
�ė��Wfބ�ln�mN��M�q�e��m��{Ը��^��wwn�6oL1VL>w����%�M�B=�F��ȇ�ǯ�Nפ�9,PL�H�z����+'d/��t�X�v�d�
��<V�30��6��Ɋ\��g�j�'/X�D��ϰ���=��Q�_��;��fg�oрC�L�_�����(�rq��|mK~B�[�_�PT5ёQa��M�+�K*g��Ҩ.��Z+��j�oXѤx����l�����l!�
�B���4t9�x4���84�1�5H��G��^F����V^݋��:���<[�BW���8�F����
b��r81�f�~.��~	���}���i�FF!��.`W;��<9��{�3װ�����N����檗��@�m��K� ��k�m�h�V�`?Opg��ŷ	]"�ϗ��o�.���\b��؂0S����:4%R^s�5�t;�T��0�I�r�7.%\%QM �,��%	���,��Z�7Ej�z'_��a�_�P]��u4^X�� ��lꏧ�㞢sֿU[â����F�5�r���o�3U����R"�E�ޯ�z�F�(��E�rFr��B�h8��y���j�M�6�d����a�(�c��wO��~
�z5~���q��'u�=�	I�V�����9�?HėN8L	˳
���\GAtl����Tmq��1�ʠF��\w�)�ZeF���P{֨�#˕� e�� �~n�/V@�w�q���O��Q��3˺���d|�,���v��n_fː	$r2	n]���l��Y`����6�1x0��3��� [�u<�������D���Á�aŮ�k��(X���8{��?@ۏ�ӓ�y��&�T��R�%#%���],;�8*0HW�aVUž���[A���Xh���xɷW����0��Y���^�����<���]�F�:oC�Ǧ$�T�}��y<�Q1{��&1h�����1a���fZ.�v>�q�e>��Ǖ�>���㼈���sp�&��>��K�p�}2���ӌ��)P�:7G(��z�H"�K1>4b����eQd�D�����[8Q�|�]��#�2Y�ح3�L]L���q@�@n�n=`I���a�q2+9(1�`_��^��~Ҵ��FfR���GJ
�;��e�⏶�KN�����8!� �������&�+�Od��8�=�\�yEIr�E�h��3��N��%@�β��o㳑��`����hEF����|D��������>C}#�(z�ˬ�K���+2Uߊx��'tk���G\����(�/�o�(�)��4�u�<�s?;z��}.M
N��A� <mɶ��Ĭ� C�dt�_�]��6�JNݎ)��VU=l�@��2�;?i&���*���d��&f^�d��T�<��=ܿr��q���ç�'HTĶ���LI�q{B�u~����w�Ã��4�!i��#�[[܏)���PO��Ɛ6��W
B3���>/��!�F)fl�[�XM�z�lZy�BcJ���Z��@u"8��IKk�����:f%[r�(097кJ6~3�-�M��O&y(���i�ٞeƲ�Ü��9'�M�)�2`V���I�e/I��bI}��Ĺ���΂��I.�����#�$Ky�
��삓���Mme=6ضf_�S�H�/*�e�rɨ!5Z]��r�ͤ�J�l0)��-?>F���<��L�>b̌�h��x����f7q�B���o����1>�{�z÷���Q a���:]p$�@B�(��Ů1䇭�.
�Ul�J��q�$J�����}��_E븯����c?Gc��(}�ڇhX%�5� �,�L����K`�zW�o;�4�nЪ�ǀyZd��L<��M��׿���`���8��b�@-�ܘp{JΘⰵP!]�Q.���V��7������D)~�󴛙�h<��\ݮsN�P][Xl{�������饜�j(����C�7��\3��%�6HR{D�%����$�/� ��-&@�ƕ�lnm'��*�)�n�u?J�}RCx��E=,����nÊ�&��SYmT�kf�*