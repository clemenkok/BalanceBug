��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�!��
��%Y l�׾�m�F��������2�pD�R]8z��~lIհ��Ԉ'��T)��"�֝�|c_-⛃Xe�T�8A����phK��ڜ�5�z/��,��M.�?"��{"�RZi

�<�I!P�F ʙ��b�P�Dq���}Д&Mv��"�j���ʦ������Xb�+c\�I
Q��i�� �~��D�>�y�ɖ����1���|P�94Dg-���g��!�� v/����&:<8����<�#˭,;����)�f�w�8���I�	���`���.�W�8U�&�~.~��=j3pW�.I~�-���|R�T�6�%�{ZzA���g5��ᓇ����,� ����r�����ߤ�{y#v�Z($Vn�jg�o�=X9�&�񑬉.0 �K[D����Æ��V��]��Ƚ�'Wi��`Z`�ա���;�f��`7W��� ��6�j���h;]GG&fEޯ_�|S98j�����5Z	�gHR>�;Sw�ܹ��U1U�y${��U��:�6|S�Wn�P�9�|�I�]����`5���袛�3��C�0S����D����\~�.�������I*������R��(�;�gхg �D��Ć�[�	�(F�84�1�?�ힳ.m�0�L�y7�о��V�1}�lP����k�j��<]{¬=?�x���r�=���e��F�{�c	y�Kxn�7��'�· ����@���MG��=FU�)l�[Fp�c�NfJ�l�(���p�K�\��i�o��GG
٩��*��G���<h�צ�eq�L�鑧1H<?*Că?�@y1��O�w��Rm�W@{׿&O�ϣX���`�`��п��]�����3��a�Y�,d	y@�u�& ��^��ҏ�`��T/�<��i�,\&��$�=��;ܚՔ�Ʊǡa����� ���K��������e�,�S�K���?��w6նo�U�h����$�H�oM�S"�4����s�'�J�~��X�C�9(��{���\�4�0��]�����7����|���!*��PRqhG��{FkЄ���/��EZ�E�d��pW-��4Vp��;3�����~��˸��y�RYUw�����)R�;R+�l��l���C9j�3J����Q���U�
���V��hڤ����&�.*����#%��Y��␜����:��`\�u�8��gO�x��*pA4��ݴ`{��}П�q��,!Ve&K�N�i����v�@G�c8e���E"�P��Q/��Y�%]�E��M��L��A%a�^�O��-L�:Ƅ����tÄF ����	8&>wv���^��ޯe���0�G� |W�l`�ݎ��'I��@�I� ��ߓ\��\̖p_�3�h���ޙNa��
V�����+�"�נ
��(��'�"k�G���n�d���&��'(���<dԔ��[��ک�G&^h�`��YV�f���:V�p�X(�b�9�:��J�$�K�'O��[%"!~����ݲ/�1���t������h�'����vU��P|Y����^Nu��{��݁�̙���o��S-�H8�P̡Ԁ`$_�+�-~f�[�o��n`���D�̑��wm��VH7�i��g*g����m��/�E*>b�1��E��1r���B���i��\� ���yK�#k) �Յݍ�LF��>T@��م�d���ׂk��� ��֬�dd�{bm�<������h8�B"��GbH.}=k?~��J{�}�;t,|oP� ?��F�S��4i.!f�f]fN�m�)���	��Ш'��ǣ��~�5�@H���/`Vd��f�GI"��0b���*O�֊�����dPmx���χ�aEǺ���
�u�B���y��F��
������@��K)6�t�r �50���1��[��ݼmܭ#��5�L�
�	��5��Z��Ԯ��f�'���t�iN,�%�a3��
:in��:�p��=gx��[e㈠�X��Ҧd�tf�'�{e��"jzX�H>�.%8~4}��C�?���_A���˹x�J{oy�Z�����YO�Oh��ыf���9H�2Ϙ�>OX�6���ia�ò{9,o��|�c��WC��iGl����2WBC.�JR,|�y�����|\.��E���OD��hDo���ן�Rv}���!�l�|3Wx[�6S�����Vg/̏�u�:sٲY�{��Z]nQ����Mǲ��J�m���'��&C'3��*��`ٲ�����@������K����p����)���ԧ��m�cU�')��Y�/���>��	������ҹ�j"�	��9_XS`~�2�k�\�E=�����$��ún~I'r����2�����б�+�����8z@�)��gK�&���N��w��e7鹠����Z���e�;,�չ,��ՓZwv��6�P�g�9��,-"�6w�p&���o�NV�,0 O�ԙ��:	��������ͫO8���d�N����W2���������ID����>Bӫ]��dq�hzO�i�����2�M;v�peA?�L½��`�.�"��J��jy:\l�{q��Yt���JB�N_N���Z�ĩ�U���g�=-�M��^@'�b	~���iڭ~[<�U�����9}�@�W����NK�TyJC8��l����Y�6�>�ٛ��K����©u�Yol5�D@L.���}#yl��Ji�[��ܖA-��`����)�s�����`����s2�È�G9�p˓N4y{� t�\�bA�T+9�ֳ���#����a֯q cnz�5y�6���W!P�F��:��=��P}�>���|hQ+�^n��L��O4��q����|���.z�U�̵�gd����,����dS��I�i�ǻ{�mӃj���f����M�:á�Q�b��{�SX&� ^1�0�:�����``�G̊;s!0_[+j�@���kd�D�n�Y,��rSG�B�wv%�z��Q9�l��j��^%�c��+T��VJ��:��E�>�ً�'�2m"�2���]�7-�vi�HT���I��������J�l�a�nf̶5_�'f�w����鴉��m��Np����i��cC� ���������U',�&ŗO2�ᶋ$0�E!S�bQk+CH����X���[*S�7rۭ�)Ә.��'KK̊T���;��\�ӧ\�~�0�6ѽ���_�)�X,��*>W�40c$/�-���DM
�x�P}U���x�g$B��(R������)�$�S�D���u3�y���Ӱ\�E��ga�L	���Y.��G�k�b-�&�ZS~���}� ���Z��$�������v$���Bh��j/�6(��Tx���_K�:*oL�q.O�B�Z�*�?����dx��v�$�n�^z?38�ѵB��*�5v���	L<���'��ч��<	�f��� dSL�[�_La=(}�_vp�s�[�f�^�'I�׵ӂ���FD��JNN��͍����<*a��+c��q��4b���XX��L�� ��x��C�̔��Ơj㳠~��Id�E�/L�|���z��h��5��ᗎ0;��ռ�T��z�<��{�@#M��:K�Z@D`�m�|�@te!��g�c�λ��p;��hm��np<*U�g^/���7~�1�#��pS|�=�����ܭI~v��nw�5R�W��{�$vjC� ǆaPs��~����,����]z�������G�T~��>+�Pn�y�}̽)�;�US~M:	��"��j�����7�������ɑ�Ů_M�	<�U�L@�ٴ�1˂Sx6�q�M���oVzդGI#ڜ4�Ldg҇�{��E1� �TC�C q���l���!i�b%R[��X�A����=_͉O�Oʳ��F��N�}��n���敭v��{�%�A�l!G�H���1vZN�{!� ��Xw�;�HӪu'�o�sk@{��<�=HȈrGAvp�lGJ�>^��:�c��a���If5@G�d�r'�m��L�Kx8l�оzc��.%�;���5�.Oq��n/:(5< x[������V��b@���p"��H��;�U����ۣ��T�a�/�h��uXpX������C�ž��ۺ��셒[x�|8�ĸ��O�-�9�At�����}b�^X�o^�7���#�=?]�I�Ř�l�{�b5ru��44�_�����N��qo��}+G*.�rR/��f �K�O?;���h���7�Z �+0g�f��n�~K�@=Εd��;(���TPn�.4�������(��D ���sd�#�RpLEB��j}�Sr�Nqj>D����[2it����%���)klfꃮm�:�{<�_L�!Ҹ��z�G-���uMb8�E4s?U�!T.Sٌ����(M �j"���Ǉ:|�[3!&��f�Y�,��B=�2F� ���B�8�[�*��*t���.���LF����?�A!�Ή����J����.�+�Ѳ���GN��P�4&h�>��$;^��#
|No2}%25�&!� �E�\��З���хI.�!�;�/^�6�QߜD�G���A��e������"��R"5�����+�S��+�K4����g��θC�?B��z��"�S����:�A�-�!FǠ���J���,�5/�� @��)	g�ZD����ߦ��Y5ˁ�	%��썦R�o6��Z�-<�d q]�C�&���U�hB��pQz�+�4���)k��znU����.Uժv�s����
�5</ruF��p�V�G���.�&v��I���<���6Z �N���/�q߯�~����������O~=HI����H�T��)i*d��ĸ"�[�q��n>b1���yw�V.���d�����zqՄ^��o��	D�[fCD���y�3��Eq��O����=�` ~�J����ّ��(iYn0��Ĳ��c�<�m��t��%�$�b�G��L�[�U��:/�����IĈ����B��<��'�Y�-b5e*ߐ���>��'Q5lC܎�e�y�Ն_�������B����B2���.����_�Oh�Y'b�L��(�cY�Y�۞L�9���Q���2T�3>���l�g���Y&t���T8I���nl���M�Vx�n���2H��#L.W��pA�%gy*�7�T���_B���`J?EC6�3�(�[�4ǚȫ�����~x��ݚq�7f����^����,�#r[����7vS��K˂�,��&_��S絓.&uSl����V�G���z-�����@b^/��n��FTz���+��,j,%�w�-6����z�H@h�o��k�-*נ+����������4�B�X�^�CI���=q�p��Ҁ�!����Q�o*O?�a���?h� =MI����=G~	�<Y"��2��~���,��նQ���\!�<I���X��я��L� �����V\�F�Qֈ���I��;z[u��Z%�]���[�̯/�	�O�>1D�m�"�5c�$�\ňF��� z�ɸǈ��[O���&\D����?j�Ku}2+�6T,z!g���I��p�2�iiI1	�cU��|	�ek86������K�!���}�����e��S��v��s�0fٖ��y�d�A���$� ��m�����W��.(B�`Ƚ{�j��?��g\��:VBk��`�ܣǀ��ѣ&�f2V�"��tYo��[-�v- �D�0�	�_ 0?���A~іl�Y$u,�Gi���| ��u��T�5����.�+�o�������:�l�x~�?\����0'�dj�A��9�J�1�?�>��cS@0�i��F����
�_L俅����V�����]P�w�K�W��n``O��H��x��q�L��q���5+O��z�0�>Z^r>��K^����}�l�|B���Wp�9 ����0*�4ʽL��{~>1Otˣ?oWȈM1���������h��=	9R�D�-��l�M);�Ce��K����4ߔ̠s8�,����*`�9C67Z�z�E�[����uh5T�$'h��㏂�0yh��"͓�'�b���~�����ĵ�'��"�8���y�g���J��B��V���P���fJZlQ`�Q1��Sb8��B	*E/<��¢J���e�>���̎�..'�E��ٹ[����4�I�3����Z�����,���Ǡ},\Tf!J�'%�n<Q_c���s�c�&b|�$���sF�$#)�y��� [�%�v�b�1��5^����:ꀞ�!2�ԯkX6c�e��F6T�[�L^�d$X�{`RV缩���#�� �o�dO ��P�F�[��H�zlX(��<�3�U�_6<o�='{�������5�g�^�U�4\��%�a�^rj{wq2�$�*n���)�L-9v���>Y1t��|���:o���a�(`�T��԰6ű�hB 4��`�<%ap���Pn�a>��q+m'�}Qk��%���"�OD����G]���)��/q��O�ҙ��ڔu<�y�d����c��hU����'wH,��pĥ|e�s���ft�J'��r8�	��uG���5d��NV�Ұ�W��ǚ5Σ��Li-{����Q�����Ź]I�Vxl���u�|�2m';�d�j��%�H��:�}�N��<t����y�Co�����Ԃ{ꥵ:C\��M�ӎ��Q���XiF^�ߗ�^1 ?T�{�I�D�Ğ��e{�cm1�rbM�R���5v�8�xh��3pM*	(r�z8�7�b�Tatΐ)�������CY��|(b���
�s,���:�^ذ�<�b~7����2Ko~E�3��9b�b+C��s�C5E��AT�2&�i�^;�I���n�T�{��C�7��0��%�ב,�Q3��@��C�˵�(��W���[/Z#�
P]�H���<W.v�_�t+��n��w!$������6���,!v��,�� i���z�`Ҟ$��������D�,%A�O����߯�6��o̻�X�3�����Zt���c�����8ө�^��.WA?�F���ĳ��?\1��I�9 �.�M�(�ȃ?�����N�]�k�n�P6Έ��ƿ���W���h&��7f���N}��עޙ��X��mߟ�<�_��p����-�`�͓��}��_�;c[�Y� ֧�0�YZ��m�1��Ů0�E<�)�Uo�-�XP�H�5h`Yp��B��y^=[K�u�ä�x�t�Hж:qr:����`����H���R-� c�N`�>�;�{�\Ұ�/$�h�g*,����y퇪J�8I�M��^������ߎN�<��m+��u�)�+P���W�r߹T@�*�A
ss�q:�6+�$\���kX8�j5��O�ۑd�
�8ԉ����>���?��5�Yo�K�����Z~gK]�~�9{ꅶ�pgf�'ver1�"����gal�U붭^$�;��C��M1������<䋂�W�f2-����2�6�H��vm;���f��N�J���1O5)u�<.6}q���S&�7�@�t�B�>Mj[����z5�^��7!qW\�_;�^�ÆF�hbܑEnw�[(�=���e/���:��DӶQs�}xb�$E6��q�z�N�	�����1NCy�F�/��Pjg�p+�ί��F˞[�i\�}�l^��iz���)e�� ��/�i��+�#ҕ4R/AG��cz�>o�I~ܔ(J�J�����W�%M��n'GRz�*�i3x��?M�zA?��M$���X�����*Kż�O�ww�q��UJ���8f\�舒��x�p�E�ٮ�ڄ,D��-��M���%�\_�����
�s���[86��i>.^��WM{m�x�{DX�}�k��5�@���M
���j#�"�V})�����M�n���A��&�"����	9��p@>�C�^~��&�,����j�c��uˑo�_������.51P H��$�����U�b��b���0�fAEV��>ź!���0��7Ap��D�Ap��?{@~�����&u�'�8��5F+H敫�P�yp�\�s%h�����z�e��|��T�49���O����yЍ�S!q� a�0��~�C���\�^���<t�f�=���/<7-�~�uF4�i��
���O��[9��X��Whx�șL�Z�z���dއu�o��S�)���kJ�
pdB����Z!�~W�6�ؖ��k�&��Ty���"e���e���<K�gZJ1A6�O�ǡ�z&�ꚙ�q�����gp�#�.lo�i*�4��>qS	vu�4��YR�cʂ'��a�xo�2~I�Aw� BR�����NX+��􅌗�O����O����9ѵ�t�C�M�x�L�c�	i��1r�G��sf0�_���D��N��I�:�`���*mj���S:ƛ���A��q����i���ŭ�}�-�;�
��R1�����<�Si0Π\���i�=��c�x�5p�1H2��MJW�X����O�t�>�O�9Nr��m��@=kf�Bq�Wz����y@���|X����!���k���{U�A:����jU/��fe��x��p�K���H����)�֕F��kH0�~db����7��W��iH��V&4;j�<-�����Q�	��� ��]O�?�	:�7*Bx��ߨ9M_xLj��%���^�8��5K��t��iC�R3��M�8 �>S�F�O�:�6��N^g#im�-�;�/�]W������2��9J*��XI���UK�:B����s�����|�4��.�LM&�c��C#��'��Ռ����j��Ԛ����F�F�9u��1cPPߚ2��~��>;�u�|�E���'��_�F�I�6��s?>��"�-�'�'�6v��)E_�O��pa<�D�m��pҳM`�:�/��j�S� ��_N@Y��d{���LQ1X<c�C�gY�m�������E�S�Z���!�J;GLCFd.��6�ߌ��,�t�S��A����΂_�!���,�4�l�H`�0��
G�!�1���AQ���3�"��%�i�
�.Lzw�1@�hwb.�Af�.v.�i.�7���~�\�o��r�A�X�O�G�W�=��Pׅ�l�Pu�sic�madaC�$e���	R��Z�a�2rH;�=�˱@s����&��OmK+Z+*�\�]�4�\+N��,K�p:��Ӽ^����0+����3?�Q�Ю�#���=��ja���Yn��/5q���<�ڍiM�>nm���ׁ�����\F�G(w���*�����&($5��{��B*�O�6�.(�նK�u������c�7髤�BU@߳cL�k�V9�Ƭ]�u����
؁8��c�=!-���h�p��@w��
�����,��eQBp��i:W�lJ�+%-!��ӕ�ƨT�a�	+ï#:4�^s����^�d���h
˂�5D�sP����d�(�uH����y�7V~kv �z�?ޛ��=��TR�SA�'S7�')�2�Qh�+��D��-��?��o�Q��y]t_˶v�����{{YXp�����3t����k1o;�@M%����6@R�9��Eg<ż��Y���7�Xq�*�&��RG>*��U�.g1ʘ�����솤llk�낪wh[���@�k�GmN`ZM64n��ڿ:��If43%��r���I������Y�]OU��!��`�<����9��+AN2�e�gOA����v6��YE2�+E/�rs�M���h24���B`}{�J� [��Y�K
�H�_\��p�^+L1h�0:�P�}CЀ 2���}A��p�hD)yrT+�{�'�F����&zA�����BM	����`|���Ϣ�'U�Nʹ���*·��+�1��돺�w�9�rG����Ʋ����1�,�S�DZK�������fwH�b�h��_�pr�1��)��p)a�j��ڟ�:�<��.�y��_Aƫk	m-��(d��	cL&��h71W0���bά�Q�o��XqO�����~����ݟxgS��^�m��6�~�UaŊ��C�CS���ZZ�Y� ll�ˤu��e�]_xfk�1���NL�Cd��T Xx�2�K,�1#e���y<1^ ���ozš�������>9��J��Kp�0l��!'E�\�B�C(�j�*\��Q���'N�Ku���tV� \�M�&����qZQ� �j ��qZL��T;s�3c�2X���l��")rH���Э��+ɒ\��5�b������C�=s��P5�h�/O��S $��Q�&�"e��.(_�囹Ý{�^�q����KPH�:Q��A����%@	�2=�e�h+�^$�"�]oN5d���)?�����"�0z�s�,W3�(��i�J�Y�ܿ;�UGɫY������-x>���J�	H2��u�1@��P��>F�3*�Z Y��.�� �a��\>�n[�G��{�I�=ρ{���K����u.��cMژ��m�x�����t]�RN�ҴM8��ASN�XTs���A�!<է2Ǹ*�q�뫒�������)h��*�2;S�vVS�Ʋ!1�^�#�H'�3!Q�Amb�ٳ��%FT�z^��� X�{�3�0<Xt(�M��H�,h�w��}̓x�ĸvGm� �xb��P7*3��S���-|+܈:no��Ƚ vN=��v`9y�A���N���[p�.׈{v�ޭ�.�ã���$�����>�/L�/wQMh�z���j���IV�N�Du�%ʳ�X�N� ft ��>�bXVo�i-i�H��x���9�|2�1���v z?s>����r�2��d��̭�Q.㯇�虻�"����B�`�ܶgC�w�)M^�&�@ر�1qR���۱ņ5A�$�'U�}��^6E��N~ԆE���Xs�وx�^�*��A4�[^��?زs2(SN�g]����{��z��K��_���$8��s����tQp[F/:A
}����'���`�����+�^�`��:�#~�oMU���z-��y`�Ui���y�zl0q�4?�HhW�\���-�B *T�y�e&��8$�\(��e�o�#@���@a:��:�-��s>n/E
�ⱦ#3�= ����Y+�N�+=�uO�R�Ǘ������H����?�Kaf ���*�+�>������|��W	�B�F;+V#?�+����5O��~�s�(�܊3h);Ƶ\3�	ӵ������7��;��~W�n���G��s��9��
�p ���rQ���	p|?�'����p\uk����e�zR/F~�D~f�N.�8�=��Tj��֭B�C!��߲�/�i�hc��.�㘡���ը5;��1bMA�
4!eN�_�v�GG���Kc�l��Wpu�k>Yj�Vbz<�(��o�>��J�`��/q��])�#3l�pB'���-ë�o�	x�xo�}�9 �cGU^�"�fLR�uH�h5h@�_�RO���Sھ�����M��?�џ���)݆u:�D9���U~�%�_����M[XZOh�XV�`�dӝ҈��o�����R���m�f�w���pl��ʱ�2\:=�۔�L� '"��\'w��{N5x�jd�s-I�!��nn¼q�z�Vȁ z��X�:�]�(C5��Ǿ��<�������*;���u)���?�;�!V���9D�7T���nd�S��CY��'�}�)Y[�dR�ݯ����L~BN�S���GS���i�-,w����Zm�aVႢ���/���o��u�Z>:�ntw�����U�7ۅ]lQAZ�Ǆ��U��<��o���0W��|vr������Z!2���M��.<��p=sP�|A������A��*߈���l!Kfb��nq�f�y~�:ȕK�`����2�j-"�I���{�-V�u�~C���o��f���	8�4T�E���6R����j��	�yNs�/�,�U�-FZ�%��s�e�d[iN[9���5b!��h ��������T����w��a^O�q��.�FB��r���
[�������p7D_�VZ�����*|?��4��b�w:�l�����Ӥ�b��ϋ|�E-+�!�5�j�P��_��T̅v��?�qI�SD�>>
�3�M/�0P�#/8`Ňi'�rJ[����sJ'5�X�هj��F�?�tq�6c��d1�����S���G�*V5D��J=�)�Fq����҉����SzS���!E`"]۾��oPI94&�@7�m9q���1�Nl�֣��$;�c'����Mqz���5-EԨ�;O��;��:��ف��)�:�N���0�m�MXQZ�H�f���� T_���,��^	��BK�/(�>����5�np��`y�Ѥ���b�/���Q��hZߞ�֧7�����z��L�<�yy`F�+E��o�6��Uމ��?����A�B��cQw[���N1���,�ֿHY�.>yBˣlA�t�t�O*lG���H>���t�\B�+k��u��P��G`��x3��i�	�?�Ao�-O$?<�/l�=�o�b�̉���'vfW�ӡ㊥7����nJ�c��W�+
c{�!��ύ�,����[�Ǹ�t���L���r�O���i�c?r|��s�<�S]�G��n��&KSS�/�^_�T���K?؏B?�CL�l=���oR:���l��K���Z�� ���l��q���G�s�D@wr��J�R	{�#h)�"�����;��P������5��)�xM�s��Y��O���4����դ�8/ș���a�g�ʆ大�g�T�����tG���Kh�0al���˄>�s+&�����P���S���� t^r������"2����җe��K����EV18��R��[΂kJ�Ta�p��;�+e�������uS=ߵ�̻9x�8��Uq��Q���؆q"��7Pv���`�L[���s��=H��t�݂���A��� �;-TkA�(�o�����P3z�p{l@c����ُ6"��N��7A��aӾ���է�$�edP_g����'D��Z9���m6B��km�xr�D��a@fVsc@ �^&�3L���N�k�۫&~��uy�q���;���S^Lu���D�(�ڲ^3��ؔ���
�G�n��<S'c�f��=�Z ��=x����2��ܵZ��U������d[�
M�Ě�{���2��#�D͋<�9�\;D�/�޵7���������6*>�KI�,�>(�J�ƿ�b���EbM�4�ɔ]�;Ƹ����9@�-7|s^x��P6ZN��x�{�Ub��q|���w)��G�D�������&�昞F!<Oⳛ�ZP>�Bh�)����z�,lG^�l���1.6�.�Ǖ�.CO���U��05� ��It��W�U-��c�!�OXЉ����1�EߚB
�\?"A.&�Q�Nh<���h	Ty��/�G�����nS�%꽁P§�����]��j�Յ�M�� A��3N6�K'k�J�2j��_�1W�E�y] lQ^56�k���a����b܀6/��#f��}�M�cI x�-b��4��ǔW���=�!�@�Tۆ�2l�A�����kʦl��zA�wF5ZO��Va��iY&%��.�����Qa͚�;�"�����.-٪��-ذP��6�hi�,�����{W��>�],��m���}�����L枘�����s��O{$P�<�p�f�44���Nx0���>�O�Vfma�Bv��n.���r�"l��*0��-]̨�,���c*L���`��A� ���(泥؊�$aW9�~�%/'-��eK�O�cє���
0'����:�By�{��	���4b��PƝ�ʁQ^��r�ƴ�Y��7��\QG�}k���᧧�?��j���}�}���T�#^�7q�]��N�]`Zޘ4R]Ŷ�Di���Z�]���|���f	��9
�� � �Į�E/2��Ϥ7��OP8��`9ah����E�"v��s%^)��&�N��V�57Wӿ�hR2�%̿Zj�;"����s�����7a/�WU�/�_:�Fj�;��<&A���PR��cE졉ڽ[��.�����Y�9W��M�H��`��M�36��Br)@�[�,�m�aOd-�_R�4�bz�Sm=t��>�e��c�w%|V�^����D����h#��Ir��<DeI1FT�gh���y�?G��`� ���M8ꏨ���_5�C�~|W�J��Q*)o��dWY��%���L�Sm�s8�s��s��<A0��1�.EH�b�˚��
����	ZU�A����͖�$�fvq�=�n
�����c�C}�6X`'d�`����w��\��!�#oIIO��Gڙ���o9_�3�y�y�3���D�7^�J�t�5%A����3<%VE�$;�b�r�����Ħ�
�8��@� _'M�ݛ�w�4�{�<st0�
�Xl����-�T��x0�r�ּ�o��<v&iT)bj�1�0=��YKm�D$Ʃw��5�3��養������G����)��9�*�v�i�K+G�����e���@�>.i'�\_�(2��nt�^�!��S�+GM�����}������_*}�"�N����؈]��i��l�4���(�ƞU� +���?N��o®������)�T��}F���%f 7DJG'��g����ca� �K�D�<�}���5����H���[�jɥ��&¢Tz�L�a��m$C���R^���P���ņ�� ���'�X��H�쌵�*{�,Q�6��J�`�� �F`���ԽB�)Ξ�~��C�9d}>��bku�&`��R㈢��g�,l�w��h,ڃ���L8�q��`������J�,����nD�ߜ+b�_t�X:���
���'�B���܍�5ۑÁq�)H�@]��/��swT���`2)��k�F`�]���Wb>iz����q?$.���p'e���d���pQ�a�N�7��s{\d�;|ɡ�u���x��2d���6#X���U�X$�Ww	�7&��^9�)��Q���L�OV�sVi=9D� 4�.�{;�X��ң�GU������۰%�nM�]=��r����2B&�*t���!Sp��~�4�l�oG
���P�Rn�@� :�~Y�жLݳ����Au����A�o���T@��2��+M!�r��	yfqL�,��6��K�d�%n}���]p���&I��z��6}��
!TZ�@(���<��T���DF���3�5����2./���ob
�|xc�����Ӌ-����!=�kG	}y�������e����,~�^� PҎ�c3�J,&�/?Ϙ�A.�pq,�/��NrdZ�ٛ��U����i\�	�
K�
����'+�l՚D}�s����Ԁ;�0ab��	ٯ4���!b*�U�M�Q,���X�f�;b:D$*��'�9 ���cP�^�%m�%�q8걟�c�k1���y��퉲�� eX�2%ݔ�%����(��ywN�g3�ބY�eEm�)��ex�q�;d5�Ͼ4��C�Uɾ�)v^63%ϙN���� ���<U��9Nm�<*T,��E�}&�<�}��Ϻ�	�Kw��/̟�G��$u�,��jc�(Tq(��	���TIdr.��1�'��;t�oh��.�CӠ�U�ӎGY��(��>�o���"��d�@Q��vߑĥŉ7��7�C�u�3`�CR��~���Z�f���P�|˪!&�Tmd�����ٷH$[��x2
n���v�{e���D�w��-u�p��1��$�.��NxZ�7k�ü�A�bq��3K�Gox�Ѿ��n�k��=�2�RK�p�duL[�d�M��*�gX
4_�L�m";t}����q s�=��)���W�Z�N��9#����}���%�'\�FW�2�*�gi
��
M��NԨ
~���,�Kں�9��^��z@[p�X�K�:��LU�#Y�:�i��j��z������bM3�1g;��GI4O���ɥ*:)f��u�����qeZ��z��bm��1fJe���Pa�Yڢ���lL�e@�+���e�a��7�u�
l� ��g�*d������g�>�8Ʃ�=^n���["�>��c�ߩtc<F$-~ܵ����-5��90�������q�)�U��U��V�>����#�Jӡ��r93�����E�7D��z�&(��m�Sr�:^yD�y���ie~�?j*iY)�J>�ܾ�U�"yI�sl�z'��&6x	V���\58:�4�;~%!kw�ڨ�0�t�*��a^4�9�����*F��Z�x��Щ8�����l@�ǡ�����]Ic�F�|߽3��u2�)�Ƌe)�r��X$aqEX(9y�8�}5h�h�x���Y�4
hވy!}�r���n�D����u��i�3�V��q�*��b�o�U&�H��I��Jw��UP��}����4�7�U��Jy�j�xP�r�%��Sq))QG^���8R+m�%�<E�Jg����Js=���VH���S�0�7L�%����Z��$r��֌���]Ȼ�`:hYHȷ �yn�[��ZXa�E(l#�t�����xb�xy�G�	��Q���E�<��,QGR	d��v��e�����UB��m������)����w�o�V$��QUȐ�-u�j�=F�\��t�E�t	����7Ik.��}��=]�g��c6�,��o��&�Ht��n�Fs�C���U��A�l��)���]Xw	�5Y)e4�<��BL<��7���d����1{_�I���#ꬨ8�3{�WuO��ì��N�*�D��𞳝�"E����+-|JM/W�܉��r��3�`�?��%v�kGt�Vo��Å�8P�S���[*�/�^ňr0m&&�C��L�ꄃ��x��aח���D��wEt�v9q��z�\�̙�!,���L'k'S������
�8�#C�̑����@�{F		���R�[.��4����VH���灋�ƫ���o��&��SX�9���WXYK�3�����e�0 yM��ymmW��%�{�C���V���cɤ?������t��q�n	�O�QOG�Tŉ<n�։	HXM`��<u�7�*�HKG�;�u#U�q��^oH��2=X�Y�^<m����P��a��KMo��:�A�R4�"���Lo���T^�5%�1Fnb � ���Jd��M����Vx �s��ݔ�i��߂�a�C��Wv4*t?�
��N��� ?�ƿ	��w��5!�~��ݖo[Ë�� fo��+�r$�c
7����C?h�2��`������7��Ջ��L���!K׫�����kHό��4Y9xN_{E����~�Oq��᡽�,,@�D�-3�0��d��t8S"��S6�DN�j�Y $�d�i�R;���sxZ��M��np�&�Ġ��,}��h���F���jm�lԹ�o݈f/��Ƚ]�t���%�l�����.&��-���H=ѭN!�����{<o#F�$J�w�xo�O�ҕ������$�oԳ�� ͹��i2�u��} Պ�d�0�O�'Pk�h
LK�,出��v͌a��M�>�Cl�Ի�f`͂;N�h��|���Υ]I<�j�ŕ1�Z�X���	8���o���[%gu�s���6�cǿC�¶���;� |40V!���c��>�:5I77��=������r�8Ռ]/[���5J����%�V�޼���:��q��j��c@��֚F��>+�y����5˓Vԛ��lN��F\p����T<�a����y�T�S���^� &�Q->$d(���R\]���J.܂Ƽq�pT����bH�T��t�,Ⱥ	@��l�OΊ���|��xF���@��Ԟ���=�=��G������^
��weʳ4	�a#?���6�^oSF�U���6��.V94髲��o��Bp�=��vE�c�5 ]	���͌9'�\���J�#``eN�P^��^*k}ld�o*�����濠���9��j��H�e����o��\nl�4�O�7|�z��Ք�B�������A%,��Q���5/�T�������1m1X�u|dKx����f��S��}��69iW�%�ͷgb�u��/L;*j%���Afs�f�2���7����q�@���2�ōCwzZ�K���]e�vlrA(�o��Ta��5p2�h��v��_����j����M���v����>1P���w�]	��A�
D��p�P�.�U�V|^�^@j�V��D�^��K'�i�rO���2V��j�
�ZL;H,\/���Y3V#�}ߵ��K��G\^�;�s�tΝj=^��ʯ ~o>��x�G�/+�md^a�"��������p	�{#��uױ�+fBྒྷT6L�B `��s�B��(�5��-��4;����R��jٲ��(&�t�ߩ��^j��=��-O�"���I^ozgvR�@�8����CnT�oOɤ�=��4ɏ!�rLG)��B�y�*��ٔ�{bْ��cֻ�]���W���fE��]�&�)�D7�����YȞ�^ߗ�3ܣ�� Dy�5�:����H%	@�/�¾�F���;���
5����@���أ
�e6����W_:ڵ孾���*�X��%�L��M<;�	F�*�$UXD(q��/�k�;&3�����f_���ʛ��SGP��g����}VIz?��#���F��5�u�G9\��IZ���x?Н����:�3��fFނ���?=��M�G�Vx�C-3GI��L�oo�>�x&�^�7l��i��@Y�6��zxz����� ��+����T��D�E�{46�2����$�ջ����PP�,�_=�ң{R��}ux��� ��Bq'�`]b�؅jdȵŝ�3�/��ӭ襆���:��v���a� W8�����0����9�$�ҷ���<�wFߐc��13�TV����C�^�e��N/���N���,A>��4(����R�yM�{Q��D޴�>'��ٶ��VW�fM�a2�W�F��vhzf"��t�v��Dc4�uk�	�_��@��s���iX3r
�� ��B�tB�<p�p	�}Tk�Aq���3�B�(�l�z��Q�S���H-Ѿ�w�k��2�Ke~?f�k/;����&$^ܮ3y�9(cŌ��:WnM�D�c�7A}��7d=c��v�?d�)u�ٛ�3v�ߦ�!>����AQ�/�d�B�I�Z߯�W��� y{Y��q'��!QkI���<�j"K�#�
����g�F�ִ��SeĖ����M1��漲�#�c���dx2w�(�H��	� �h�U:D�E�-F$��R�0�[�b	��*�=�,����|�)X�Zы#7ؘ+�� �x_ּ���Q��"C�'_�.�q�'�*�6�ӑ�x�����������"u:���r������^�yخ���M?����3���R�}1�R���e�/`���R��{5ˌ9�C\�?�>(	�p�髕�:U��qO�Ü�oj�B{5R�9�iN��I�����'��̤��s?�:#�M{�G�tŁ�Ӛ�Z�ǻ�#3��R`E��F�<�ǅ�Y��+�s���,]/z00,-5�e�\����ǆ�׼��iq�G��G{"�!um'����Z7��/'(�lǧ����^��EdSg~�SE�o0Q�s�l��	�4��[�E��ժ�a��]�$��Mr{_�����۲�݃"^~F(]<���RY��8��]o	�. ���P��������Pp��-h[E��͝�Y��X�+���%�Z��))���P��+-�C�zj�7�n�b|Ҧ�B[:�d���aO�h��#rꏰh��
�2�tK��X_���/T�(�x-�^ڏ<��J�����o���X�QK=c�<=n"3���pY�CJ s��I��"�Z_-�lX�Wp�L����ක-�3\5��2�f��.M���ã�d}�kO�\'vV�i�?�C�wHn��Y�(+�q�h�Sr$q����M	lD����ol���ޤs�ה�z���B{�b�XI���b�jQF��R���rк���S�i��A�<f:����ʿ�")�x�O�[�vƥ��)i�x����#xT����g�[y����b�Ct�ȑs��y����6Aq��ȱr�v�@P3o[�I�=H�������:����"������zL������C�5��'���BjHM]�Pb[���?6����/wx�;T@D��k�Y,���m��l�����J/4��{xd��i"-C�nr�:��ƔJ�	L�ti�Oo�,*l�������'�ۢ⩕��e��j��qEcax5�`n�hG,+�Ho�����4CT`�݉n�.�BOYE��M���/]/*b��z�2��9(��h��/w�s�|~����$�/:�:{�_Ӆ%���D'� ��>�	3/&�e:T˅,ј�R�j�H�<+1����-�b`����~�� ��"�;xh%�<�=Y�+������J쑪�T��� ��#�lGeB��t�l�����A���l'b���� I$�C�jם-��%��I�I�%V#&C����3L�������9/�]~7���_Q�c!����)�&@�W�:����pG����P�� ��PQ*v�_(Y���%q�-����H"m�c��B������ v�\L�e�j�oi4�|{9�X��n+���]�@���iT�<�i��# ��u�XS�R��q13�'�>j6�>كC�W)��fm��S}���Z��-`S��b����$W��ێ�gA�vĳ���*���[_3��<��a5��&k��˴Ivw��l����G�/�>J� ���![w/��bmO��M���)��{�g7�?�w�63�Z��|H����2_��%Q��������rw��]��Z�^�݊D�C����~	ԯ��t@6�A���V(����"F<Ȩx�e�����Ŵ�����~F`����f�jZ�EYeJgU�M�)ȵ��䨁�ί�%9.�B�3�|]�+�g��{N[�(������+N�)mxk��7�~�3ҡɛ��b ��u�IOdO�%~��������K���3�
���-9�G'�w��Z�rW�9h���$�Fd+�g��AlO~����S'1i[�.~a?�M�@�`�k�(�N"�{f����Z�껿>�Đ)KE������&�57��B8_`{� (0ф5��,�@(�%lF����&_��4���=;��)�� ����"�_��I
���� [F�^����ȥcm����`K8� MgJ��?>%e��b3���o�>�Ķ*c]����*��l7q�4�mo&�9!\u{�������$b�4@���%#E1�33��QY>���v~Z�$���ز0'�|���e�!�Ky�۱�N31���E%gFA}����8o��+�<�!��Nzd�a�c�}�"c���(�=ā�
�U`��<���pq�a�_���M{R���GdOw��bƊ���;H���V��v\�@[��L�C����9���C��uJ[����(��Q���?���4{�D���b���e����Q��s˕��5/��n3kkI$ݺM��4�֌|J.Fm�|�k�T���Һl���Է��{gt�A[]"��BE�5��+k�7nNr�fb��Y�ɜ�2|��}��7�פBs��Gd���TP��kP�7=����%��v��'H���=�Z�����
����)9��+�ӭr#���M!Aނ���}��~q�QU<>�����6��3�k���eae�!vBk�d�9�w�G�c_Ps��{.�M_�)r!�$-�(HO��F�.R^LE�M�_M؋C�~F�m����w�R���LzmO꯳RD�W�.��V��buj��h���K�9�["�M�������S0��U܉��1?sta�B߃��4�)`��Hn�wt�s��[#�żHu��#���\��:�9��L�n��?���K��"�����l�"3���$I[��g���>�)�Ke��'���n9t�k���T\ƾg1k``�W�q���L��`�_�����i��5iŪ���xb�F��sL��$`�N'Wղ[��GΊ�{�5ח�h;p�z�(_K��_+O"�m}�/�T�Ƅ�~�� ��Tp�v�N(��.���f���b囦
��������:���?��핏S���
��D�O�|�щo@�K�?���bN/�׀� ����[y���y��-:_�I���bM���\��ɣ�]�� �����DsRy��C��)�/��A��%\���0_�:�,ДxeG�j'k��߄M�	1�`v�,Q��k���esP/�I83�4�
8��yC/ᑠ�|�U��C�D3:Sͱ��̔4���g5�(Mʚ����'�]�tM@o+�]���v���3â\7��I�HN�V3>�P,c�݀,��<�\pep�N�/�,�t��,ċ�^�ZU*w��IHg��3@���e���[�+ʦ-���N[5���8��@%5��`:�k\� ���w�V�ǰ��״j�'�P�[x6Ku'�D�0x6�텖�� (�����;p�� �����*\�u2�[�Ȏ:�݉�n�<8��_^d�RV:S���[膿��ڎ�$�����=ρ���[\�q��	{]/R�T)���J8D����'4�)_��"��DAyf(��0xF;�K��n�L��ʧ=|/�a�#1h|��3$3Ƚ�@s���!��I7Yb;_���&�f��Ḃ�pґ���E4jxq�� [����ԬaIhQ��#U��3��S�?��,RJ�C)�A2kt&�(�m�u���Ϻ?Sf��Yg2o��̸�x�㕵}��wa��;��C������1}��VMOQ:J:��9�Nj��d �&-�����x�f�%{���$�l���d+e�3]����M!�9�!U��zXz��mq09V/���G�s��W����2L�m޴��!#2��z.`�2I^�1X8�i~ƝC7�B��4���������\wh@�rz�wA�R�&Ф�p����za��`� �]�6s_mV?�:��O�h�V�p�(2hJ�׺�%�\�V�2��U�W��r� �Ř!��0�Vny�خ2�IT��.϶�k>��'�����9vq��e�g���c9p�(�� qim�6Ź}��o�k����P��~WU17��	�X;U1�_�&x��M_B���f��dP������7 �@�3���j��D J��z1k�:�Ɗ~��si
2�v