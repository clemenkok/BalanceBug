// Qsys_tb.v

// Generated using ACDS version 14.0 200 at 2015.12.29.11:38:54

`timescale 1 ps / 1 ps
module Qsys_tb (
	);

	wire         qsys_inst_clk_bfm_clk_clk;                                 // Qsys_inst_clk_bfm:clk -> [Qsys_inst:clk_clk, Qsys_inst_reset_bfm:clk]
	wire         qsys_inst_reset_bfm_reset_reset;                           // Qsys_inst_reset_bfm:reset -> Qsys_inst:reset_reset_n
	wire         qsys_inst_i2c_opencores_camera_export_scl_pad_io;          // [] -> [Qsys_inst:i2c_opencores_camera_export_scl_pad_io, Qsys_inst_i2c_opencores_camera_export_bfm:sig_scl_pad_io]
	wire         qsys_inst_i2c_opencores_camera_export_sda_pad_io;          // [] -> [Qsys_inst:i2c_opencores_camera_export_sda_pad_io, Qsys_inst_i2c_opencores_camera_export_bfm:sig_sda_pad_io]
	wire         qsys_inst_i2c_opencores_mipi_export_scl_pad_io;            // [] -> [Qsys_inst:i2c_opencores_mipi_export_scl_pad_io, Qsys_inst_i2c_opencores_mipi_export_bfm:sig_scl_pad_io]
	wire         qsys_inst_i2c_opencores_mipi_export_sda_pad_io;            // [] -> [Qsys_inst:i2c_opencores_mipi_export_sda_pad_io, Qsys_inst_i2c_opencores_mipi_export_bfm:sig_sda_pad_io]
	wire   [3:0] qsys_inst_key_external_connection_bfm_conduit_export;      // Qsys_inst_key_external_connection_bfm:sig_export -> Qsys_inst:key_external_connection_export
	wire   [9:0] qsys_inst_led_external_connection_export;                  // Qsys_inst:led_external_connection_export -> Qsys_inst_led_external_connection_bfm:sig_export
	wire         qsys_inst_mipi_pwdn_n_external_connection_export;          // Qsys_inst:mipi_pwdn_n_external_connection_export -> Qsys_inst_mipi_pwdn_n_external_connection_bfm:sig_export
	wire         qsys_inst_mipi_reset_n_external_connection_export;         // Qsys_inst:mipi_reset_n_external_connection_export -> Qsys_inst_mipi_reset_n_external_connection_bfm:sig_export
	wire   [9:0] qsys_inst_sw_external_connection_bfm_conduit_export;       // Qsys_inst_sw_external_connection_bfm:sig_export -> Qsys_inst:sw_external_connection_export
	wire   [0:0] qsys_inst_terasic_camera_0_conduit_end_bfm_conduit_pixclk; // Qsys_inst_terasic_camera_0_conduit_end_bfm:sig_PIXCLK -> Qsys_inst:terasic_camera_0_conduit_end_PIXCLK
	wire   [0:0] qsys_inst_terasic_camera_0_conduit_end_bfm_conduit_lval;   // Qsys_inst_terasic_camera_0_conduit_end_bfm:sig_LVAL -> Qsys_inst:terasic_camera_0_conduit_end_LVAL
	wire  [11:0] qsys_inst_terasic_camera_0_conduit_end_bfm_conduit_d;      // Qsys_inst_terasic_camera_0_conduit_end_bfm:sig_D -> Qsys_inst:terasic_camera_0_conduit_end_D
	wire   [0:0] qsys_inst_terasic_camera_0_conduit_end_bfm_conduit_fval;   // Qsys_inst_terasic_camera_0_conduit_end_bfm:sig_FVAL -> Qsys_inst:terasic_camera_0_conduit_end_FVAL
	wire         qsys_inst_alt_vip_itc_0_clocked_video_vid_v_sync;          // Qsys_inst:alt_vip_itc_0_clocked_video_vid_v_sync -> Qsys_inst_alt_vip_itc_0_clocked_video_bfm:sig_vid_v_sync
	wire         qsys_inst_alt_vip_itc_0_clocked_video_vid_datavalid;       // Qsys_inst:alt_vip_itc_0_clocked_video_vid_datavalid -> Qsys_inst_alt_vip_itc_0_clocked_video_bfm:sig_vid_datavalid
	wire   [0:0] qsys_inst_alt_vip_itc_0_clocked_video_bfm_conduit_vid_clk; // Qsys_inst_alt_vip_itc_0_clocked_video_bfm:sig_vid_clk -> Qsys_inst:alt_vip_itc_0_clocked_video_vid_clk
	wire         qsys_inst_alt_vip_itc_0_clocked_video_vid_v;               // Qsys_inst:alt_vip_itc_0_clocked_video_vid_v -> Qsys_inst_alt_vip_itc_0_clocked_video_bfm:sig_vid_v
	wire         qsys_inst_alt_vip_itc_0_clocked_video_vid_h_sync;          // Qsys_inst:alt_vip_itc_0_clocked_video_vid_h_sync -> Qsys_inst_alt_vip_itc_0_clocked_video_bfm:sig_vid_h_sync
	wire         qsys_inst_alt_vip_itc_0_clocked_video_vid_h;               // Qsys_inst:alt_vip_itc_0_clocked_video_vid_h -> Qsys_inst_alt_vip_itc_0_clocked_video_bfm:sig_vid_h
	wire  [23:0] qsys_inst_alt_vip_itc_0_clocked_video_vid_data;            // Qsys_inst:alt_vip_itc_0_clocked_video_vid_data -> Qsys_inst_alt_vip_itc_0_clocked_video_bfm:sig_vid_data
	wire         qsys_inst_alt_vip_itc_0_clocked_video_vid_f;               // Qsys_inst:alt_vip_itc_0_clocked_video_vid_f -> Qsys_inst_alt_vip_itc_0_clocked_video_bfm:sig_vid_f
	wire         qsys_inst_alt_vip_itc_0_clocked_video_underflow;           // Qsys_inst:alt_vip_itc_0_clocked_video_underflow -> Qsys_inst_alt_vip_itc_0_clocked_video_bfm:sig_underflow
	wire         qsys_inst_sdram_wire_cs_n;                                 // Qsys_inst:sdram_wire_cs_n -> sdram_my_partner:zs_cs_n
	wire   [1:0] qsys_inst_sdram_wire_ba;                                   // Qsys_inst:sdram_wire_ba -> sdram_my_partner:zs_ba
	wire   [1:0] qsys_inst_sdram_wire_dqm;                                  // Qsys_inst:sdram_wire_dqm -> sdram_my_partner:zs_dqm
	wire         qsys_inst_sdram_wire_cke;                                  // Qsys_inst:sdram_wire_cke -> sdram_my_partner:zs_cke
	wire  [12:0] qsys_inst_sdram_wire_addr;                                 // Qsys_inst:sdram_wire_addr -> sdram_my_partner:zs_addr
	wire         qsys_inst_sdram_wire_we_n;                                 // Qsys_inst:sdram_wire_we_n -> sdram_my_partner:zs_we_n
	wire         qsys_inst_sdram_wire_ras_n;                                // Qsys_inst:sdram_wire_ras_n -> sdram_my_partner:zs_ras_n
	wire         qsys_inst_sdram_wire_cas_n;                                // Qsys_inst:sdram_wire_cas_n -> sdram_my_partner:zs_cas_n
	wire  [15:0] qsys_inst_sdram_wire_dq;                                   // [] -> [Qsys_inst:sdram_wire_dq, sdram_my_partner:zs_dq]
	wire         sdram_my_partner_clk_bfm_clk_clk;                          // sdram_my_partner_clk_bfm:clk -> sdram_my_partner:clk

	Qsys qsys_inst (
		.clk_clk                                   (qsys_inst_clk_bfm_clk_clk),                                 //                              clk.clk
		.clk_sdram_clk                             (),                                                          //                        clk_sdram.clk
		.clk_vga_clk                               (),                                                          //                          clk_vga.clk
		.d8m_xclkin_clk                            (),                                                          //                       d8m_xclkin.clk
		.i2c_opencores_camera_export_scl_pad_io    (qsys_inst_i2c_opencores_camera_export_scl_pad_io),          //      i2c_opencores_camera_export.scl_pad_io
		.i2c_opencores_camera_export_sda_pad_io    (qsys_inst_i2c_opencores_camera_export_sda_pad_io),          //                                 .sda_pad_io
		.i2c_opencores_mipi_export_scl_pad_io      (qsys_inst_i2c_opencores_mipi_export_scl_pad_io),            //        i2c_opencores_mipi_export.scl_pad_io
		.i2c_opencores_mipi_export_sda_pad_io      (qsys_inst_i2c_opencores_mipi_export_sda_pad_io),            //                                 .sda_pad_io
		.key_external_connection_export            (qsys_inst_key_external_connection_bfm_conduit_export),      //          key_external_connection.export
		.led_external_connection_export            (qsys_inst_led_external_connection_export),                  //          led_external_connection.export
		.mipi_pwdn_n_external_connection_export    (qsys_inst_mipi_pwdn_n_external_connection_export),          //  mipi_pwdn_n_external_connection.export
		.mipi_reset_n_external_connection_export   (qsys_inst_mipi_reset_n_external_connection_export),         // mipi_reset_n_external_connection.export
		.reset_reset_n                             (qsys_inst_reset_bfm_reset_reset),                           //                            reset.reset_n
		.sdram_wire_addr                           (qsys_inst_sdram_wire_addr),                                 //                       sdram_wire.addr
		.sdram_wire_ba                             (qsys_inst_sdram_wire_ba),                                   //                                 .ba
		.sdram_wire_cas_n                          (qsys_inst_sdram_wire_cas_n),                                //                                 .cas_n
		.sdram_wire_cke                            (qsys_inst_sdram_wire_cke),                                  //                                 .cke
		.sdram_wire_cs_n                           (qsys_inst_sdram_wire_cs_n),                                 //                                 .cs_n
		.sdram_wire_dq                             (qsys_inst_sdram_wire_dq),                                   //                                 .dq
		.sdram_wire_dqm                            (qsys_inst_sdram_wire_dqm),                                  //                                 .dqm
		.sdram_wire_ras_n                          (qsys_inst_sdram_wire_ras_n),                                //                                 .ras_n
		.sdram_wire_we_n                           (qsys_inst_sdram_wire_we_n),                                 //                                 .we_n
		.sw_external_connection_export             (qsys_inst_sw_external_connection_bfm_conduit_export),       //           sw_external_connection.export
		.terasic_camera_0_conduit_end_D            (qsys_inst_terasic_camera_0_conduit_end_bfm_conduit_d),      //     terasic_camera_0_conduit_end.D
		.terasic_camera_0_conduit_end_FVAL         (qsys_inst_terasic_camera_0_conduit_end_bfm_conduit_fval),   //                                 .FVAL
		.terasic_camera_0_conduit_end_LVAL         (qsys_inst_terasic_camera_0_conduit_end_bfm_conduit_lval),   //                                 .LVAL
		.terasic_camera_0_conduit_end_PIXCLK       (qsys_inst_terasic_camera_0_conduit_end_bfm_conduit_pixclk), //                                 .PIXCLK
		.alt_vip_itc_0_clocked_video_vid_clk       (qsys_inst_alt_vip_itc_0_clocked_video_bfm_conduit_vid_clk), //      alt_vip_itc_0_clocked_video.vid_clk
		.alt_vip_itc_0_clocked_video_vid_data      (qsys_inst_alt_vip_itc_0_clocked_video_vid_data),            //                                 .vid_data
		.alt_vip_itc_0_clocked_video_underflow     (qsys_inst_alt_vip_itc_0_clocked_video_underflow),           //                                 .underflow
		.alt_vip_itc_0_clocked_video_vid_datavalid (qsys_inst_alt_vip_itc_0_clocked_video_vid_datavalid),       //                                 .vid_datavalid
		.alt_vip_itc_0_clocked_video_vid_v_sync    (qsys_inst_alt_vip_itc_0_clocked_video_vid_v_sync),          //                                 .vid_v_sync
		.alt_vip_itc_0_clocked_video_vid_h_sync    (qsys_inst_alt_vip_itc_0_clocked_video_vid_h_sync),          //                                 .vid_h_sync
		.alt_vip_itc_0_clocked_video_vid_f         (qsys_inst_alt_vip_itc_0_clocked_video_vid_f),               //                                 .vid_f
		.alt_vip_itc_0_clocked_video_vid_h         (qsys_inst_alt_vip_itc_0_clocked_video_vid_h),               //                                 .vid_h
		.alt_vip_itc_0_clocked_video_vid_v         (qsys_inst_alt_vip_itc_0_clocked_video_vid_v)                //                                 .vid_v
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) qsys_inst_clk_bfm (
		.clk (qsys_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) qsys_inst_reset_bfm (
		.reset (qsys_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (qsys_inst_clk_bfm_clk_clk)        //   clk.clk
	);

	altera_conduit_bfm qsys_inst_i2c_opencores_camera_export_bfm (
		.sig_scl_pad_io (qsys_inst_i2c_opencores_camera_export_scl_pad_io), // conduit.scl_pad_io
		.sig_sda_pad_io (qsys_inst_i2c_opencores_camera_export_sda_pad_io)  //        .sda_pad_io
	);

	altera_conduit_bfm qsys_inst_i2c_opencores_mipi_export_bfm (
		.sig_scl_pad_io (qsys_inst_i2c_opencores_mipi_export_scl_pad_io), // conduit.scl_pad_io
		.sig_sda_pad_io (qsys_inst_i2c_opencores_mipi_export_sda_pad_io)  //        .sda_pad_io
	);

	altera_conduit_bfm_0002 qsys_inst_key_external_connection_bfm (
		.sig_export (qsys_inst_key_external_connection_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm_0003 qsys_inst_led_external_connection_bfm (
		.sig_export (qsys_inst_led_external_connection_export)  // conduit.export
	);

	altera_conduit_bfm_0004 qsys_inst_mipi_pwdn_n_external_connection_bfm (
		.sig_export (qsys_inst_mipi_pwdn_n_external_connection_export)  // conduit.export
	);

	altera_conduit_bfm_0004 qsys_inst_mipi_reset_n_external_connection_bfm (
		.sig_export (qsys_inst_mipi_reset_n_external_connection_export)  // conduit.export
	);

	altera_conduit_bfm_0005 qsys_inst_sw_external_connection_bfm (
		.sig_export (qsys_inst_sw_external_connection_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm_0006 qsys_inst_terasic_camera_0_conduit_end_bfm (
		.sig_D      (qsys_inst_terasic_camera_0_conduit_end_bfm_conduit_d),      // conduit.D
		.sig_FVAL   (qsys_inst_terasic_camera_0_conduit_end_bfm_conduit_fval),   //        .FVAL
		.sig_LVAL   (qsys_inst_terasic_camera_0_conduit_end_bfm_conduit_lval),   //        .LVAL
		.sig_PIXCLK (qsys_inst_terasic_camera_0_conduit_end_bfm_conduit_pixclk)  //        .PIXCLK
	);

	altera_conduit_bfm_0007 qsys_inst_alt_vip_itc_0_clocked_video_bfm (
		.sig_vid_clk       (qsys_inst_alt_vip_itc_0_clocked_video_bfm_conduit_vid_clk), // conduit.vid_clk
		.sig_vid_data      (qsys_inst_alt_vip_itc_0_clocked_video_vid_data),            //        .vid_data
		.sig_underflow     (qsys_inst_alt_vip_itc_0_clocked_video_underflow),           //        .underflow
		.sig_vid_datavalid (qsys_inst_alt_vip_itc_0_clocked_video_vid_datavalid),       //        .vid_datavalid
		.sig_vid_v_sync    (qsys_inst_alt_vip_itc_0_clocked_video_vid_v_sync),          //        .vid_v_sync
		.sig_vid_h_sync    (qsys_inst_alt_vip_itc_0_clocked_video_vid_h_sync),          //        .vid_h_sync
		.sig_vid_f         (qsys_inst_alt_vip_itc_0_clocked_video_vid_f),               //        .vid_f
		.sig_vid_h         (qsys_inst_alt_vip_itc_0_clocked_video_vid_h),               //        .vid_h
		.sig_vid_v         (qsys_inst_alt_vip_itc_0_clocked_video_vid_v)                //        .vid_v
	);

	altera_sdram_partner_module sdram_my_partner (
		.clk      (sdram_my_partner_clk_bfm_clk_clk), //     clk.clk
		.zs_dq    (qsys_inst_sdram_wire_dq),          // conduit.dq
		.zs_addr  (qsys_inst_sdram_wire_addr),        //        .addr
		.zs_ba    (qsys_inst_sdram_wire_ba),          //        .ba
		.zs_cas_n (qsys_inst_sdram_wire_cas_n),       //        .cas_n
		.zs_cke   (qsys_inst_sdram_wire_cke),         //        .cke
		.zs_cs_n  (qsys_inst_sdram_wire_cs_n),        //        .cs_n
		.zs_dqm   (qsys_inst_sdram_wire_dqm),         //        .dqm
		.zs_ras_n (qsys_inst_sdram_wire_ras_n),       //        .ras_n
		.zs_we_n  (qsys_inst_sdram_wire_we_n)         //        .we_n
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (100000000),
		.CLOCK_UNIT (1)
	) sdram_my_partner_clk_bfm (
		.clk (sdram_my_partner_clk_bfm_clk_clk)  // clk.clk
	);

endmodule
