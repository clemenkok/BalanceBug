��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�!��
��%Y l�׾����|R�bD�E���y"X־B�ZdEy�\��4�YH���G��?����֝���[3�0�&3����v]f� ��d��A��r�I�>�W*�.d��OH?����m�'�;̿�[r��t����B� �m��6��7No'0LvE���������S���
�)J2p��#(�
%�·X��^��e���4�����A2����E�<s,��6��pV�����Mq�&P�\�bB���U������Y��[��$�4g��~�G��))��Q�
9ܱX7%�#�^m���|�	EV��3s)���%p��g�/�&0X���I�}�q ��.�`�Β��L�����/�J�byv��]�3�����*�A��r$`����t8�"�v5����k�m^����_@�e���O�]熽���cN
\�O�63��VH���v@ǽ��R퀰:QH�?���>������EN����%,8^gן$����#�}�Q6UH����|�� �Y���1^�	-����_��, �t�r��[˲d�c��kQU�au�i� �K
����^��kV������W��T@�1�Ѐ02+m-HC����t g�]НM[���<���:h�/Gg�z�t:���[:����4��˿�2��+�(���=�7���W�v$l�C�߀��!���09�e����a9?�H�Td�qGϕ$F=MS�+4DB4=�t����|�������
oX��xm\�Ŋ��Z���	��+�w?�o�ιt�Rj����O���[̍��J�����`�(h[��e9��ֱ�p�}��
'��H��eX��9m�����5 �(au�����h�* 3S�'�=7:��5�0qh-m$0!�<�ƙ�w&���#qj�#8�Į9Էk�0�j�J�/o�nş0�4�Z���ȋG�F���#*U���R�������'�B0Q܈Lu���䊳��Ok�0o��K�1N L�Bp�b�����`) CmI^8���%��L�.�Ձ�{�x� �q$��(��c�ʚ�s�/.q�2�uY�B�/�[�x�����e�+A�ӄ����eo���F���A��2�壍�JG_��I�P�N�U�VfS�x.[&��/�U��S�0{���Lt�I��)\MM�K�Q����yd^��(=wE������wI�A2�;;�����;ZC�oCK�����"VD�rB�S ���"��w�+�{4�}�9 CT�����n�=aE�^e��v;���e����]xT���Q��'�C�`��`}C^�M�m:19�@͊YA�	z9/��xd�V�֭�c'Niv��2*j^V1�e�;cm=p�ZAq "m1���W)�P����w�[?Ɛ:����'�)܀��z�NR4f�أ�X���3�z1B���4\1�g�"�L��dK4lós_�%�e�\�NEq �ח��kA�7ռ�0���l~/pԧ�n{�}��I�_��mp�kC�'߳PaA��P�^u�:|�����M�yD��5��<���U��6.�MlRa�t��`�D�7��7��bۼ���K~T��+k=�/��7ͤ�!��\j�h�_>�<���NUs~5������ lحo��
�K�wQW���X�-� >tis�����?����<E�'�`M?��ɥ�'���������[��֛���vS�?��Y����)�ZJHz�����Cn��ނ�/�����2��԰MH0ԅ��҉�&.�����b��e�K��{���tcҨ{��g\>�#	�F����.(%�_7Dh��h;�l��Q�{^�<ab��+�a�Q����h�=��l�[��!Qt�),֍���W��O!�7�Ϗ����u{�Mg'�Hǩ��&��V���}�I�"�c�\�<A�i+&��������h�����X� �b$����|�Na�&�Kܿ��7vfK�
�R� �y!����ard��d쐫w�~�'���>LLV�]�V�oB�~Q��a�>!�Ň g�'�|���l�3Ӑhvt1���[��3����0�Hշ*v�Ԑ���4��l�&�*�0]��u�{	]@n�& ��b���Dw��&�H�����p8F��&�4�ܡF����!O�����/o��Հ`<��g�
R��a�+�AV��K�IK-f��,����\�'�ۊ�����CP�F|? ��S&B��î��#o_�݅O	Qć>;`T���]޸��S�>�⦃�A�3cƜf�6|<�<|��;�WN�5| g��]0w��3A��*��3r�i��۞'[�V�k��7f{�MRGp�[�BY �uq��,�D���DI�r�(�&&�:���h�v��8�E5�4�y�ON ��7�Q��uс��ѡ��X`�>n�dYjV�]^H����G L�GF��Mh��s��9"�=�1K��\��Ny�n�(�g+�+f��E7{٨Mn��>�8�Ꝝ�9};�g.��a�'�ss4)�`%-ɸ���jvR!5h�5��X���v[���c�C���'�.\�����=�Jr`��_����\u�g�R�{�_iH~z 	܅z&V� �yY3ϫ����c��$}����}���Vh��h����/�����ާ��������?T�-��_��|����;��3@������ݾ�q�_��e<q��-$��#���$ZΤVd��&#ߕa��5OR��6�Ƚ�]!t�,��������2^s�@�����a
��a�ksG�c��h��A�_�Л՜V�W[�Zo&N!�E�O��W��~���]	ڪ�r����@�����Kc�C吇�M��Ōc�}��=d�����K��t�v�GE?���*�/���dD>�6MQv:Gg���$~�������I�'L<9X<y��Jsh�:����N���Z��yy!�iR�Y����<H�-=�h:���Z�I(S�2�y�@ﵚ0d��C�+�kJ-���F�5����!���*����;/�p���({���3��mw��ɝj�V!e-�i|l����Z�T[S&% ��I\�K(x_���eO�G�Z��N)����|nд�iby��b�HK`�1�E��J��VG��U�'o�%��(�3oY��J�(P]Mu �T���A��&��Wd]0�oA�.���L��vہ��V��
JZp��F��CX�!���2x��,��M~a/��ɔ�U���}c�U���N���������U�!UB@@%���
�����(o��\F���:��^E�ӌ��9^�k���GQ�7�ޘ�Bqi�nQ�a�72�h�tx}!)ދ3^E���8O��9�<_�}�&fC���\�8f�'T�:�}�*��b ���p3ñ�#5�W%�L�9�/�iHNs��P�ov�A��#��v��3���c��j�Qˡ�m@��.ȣ����U�y( 1~�M��Y}�����^{V9*�8�X�rk��GX�1e�&��h��e�KDyԫဩ&�<M2��;��_��,��EO��e����Qd�ȨgU:8���&���/e��B���0H	�=W���'�O���R.
M	"d\֞r�w�XMw�?��K+b�����%wl,m@6��1��$r~3YXe�S�Tϊ"������.HÆ����?T�1� ��Dv�4�`?NMw4?G��,����B�w8���$���o����i��i���eܵ"MD1��u�Ds�jg��-|d!���>�f��ʴ9!s\���w�*O݇Ha|'��R�ThY$�:����t�,!~��~iՊ�ޢM�v����F�k�A�J�&����&\^�*�ؗ�/��8A�Ba,���cr ��y�g��LM[7�=c�5w����[:�e'��)C�TS��\���?�
�Y_}�$5.��C!����D)�兑*������:�h�s��Bu��z�`��M��Β�]K���� �Ff"��~\�övյ�|��F������󀁰0LY��ۯ�Z��Q�s��^;݅Aɒ��2,���/��rd�]+����dKD��gg���|���� X�A{r�vH/�1"�
���J��K�0-t���c��?e}��=�n�fkzn�Х9Կ�&����Jv�|~3sXO8���0�s�⡬�����%l��M�"ƴ�f����h�"��'r�R9+#B�[[I��fԢ��̓0�K�Ӹ/���T�C�Y�%�kϤ%�� ]5���:����&_��(�!����Yj�!�L�Zߐ-�)&&�?�T��QU���{�dE�{NW��%�n�rr�T�$M$�-Ub@ȵ���DN$ӘA�&'�	�9Q%T%ez)@���4"��ݙ͑.�5�>Q�g�ސe��e�x��N�u�`�q:_����Ή��a{��]Ie%�v�LGY�:��R$=�kF����r�`�t����%��Vy�I���nQ13�ߖc,�(���u����֑k�r����J)޻S�t�6:��`5X�~�<�r��3&�� 2�= b�Tª�v4�O"���6�ʈ�L{h<��������:\�k�D�P^R֚�9k$U� �&d�P��T��?n)��!�+�Os�� �Kz�k;UbbyG�P�ǥģ3Π��F��S���W����y����t��l�x�����c\�����y��R�!�ԛ2>���a-��Y6�gv���=.�u����!Gm�5~��`]���^G�('�n!ۙбA1m.~qv�C3Ьٓo���RU�����Šj�_(@ٰ:���͒K|kM�|�u~ב%����6������Y���o�Q����"��ޓ.��Ҡ��[�5��%I�f{ۃ�s��m�t�Aw���׬>.^Դ{�2�V�z��h��@�Zj���q}��eTv�&�u���G���yy�y5t��x��aC�����TfJ�AP2�NH�`ٶ�O�>,���اv�Q��W~f�~H�|�����P�� <��x*;|"y�bDM`�#�*�̇�aj|��渨aI������@�C��hT���L	1��7�b��������dA;���"������oP������[�Ӌ��b{�|���O\�O����D�.p�dG�����L?w0/J"��MN�Y:N�O����.�FI:S��&Aq���P��,pNW�pTF���D�s@��Z�{C5���q9% ���-��~�䁓u����ls��G/] �Da��u aY�%
g�_�n[)nm����������S�;lKWp
	=Q�7?�H��f�Q�#�'��!��ff°�C�Q����F�����Wlԁ�l��ս6C�Ҿ�۴~�ɀg��<rHv�����_K.���D��py *�Ҭ_��4�-��(݌�yv���	E�DmK�.�N7���z��,�g(+�tJ���@J���6���O5D8s��יwٙ�[��O{0�Qs��1�n�F=�Ï=�̯�D%���MChj�'��X ��9tڇ?��n£��?�ꊴ��(�xm�+a���s�ϨF)khr�ػN��4 Ř#0xn�;�]��_���?ȱ槊�NYXd��<�q2I�2�r�&?v<.� @������B���O��m��_�����%�ҿ�ޱ��� �[c���-�����p���4#M�?;��PE�
7p�;�?b�AZ,�Y�`�bFAi�اX��L�V��My��G�G��&x���*��_m��s���I)Q@�@1C�-�9Ph���o=#!V'����'�����ݻ~��~-N)+@�G�Y��e'd���h�jN*�zK��%:X{qɭ�DRr�t�Yĵ�(��>���-�KB�"ۑKj�w���F	N闎vc���r���g�V$p$�7�����fRظ���� �^R:��w(�jA��e�6U?`�˂z=��=����*@g���0����ˆtQd�t�B�L��m��?�`-����Cǟ����JS^�T�g��A�v���0+zbs��������o`�琦��j|\	��ꨞԸ�>��P�!�)I�Z�p]Sr�>y��s�)n1�O�Uۂt��@r/7��F� ԗZ"���O��N�yC�O�������Tl��v��JF�ɧ��~��d�Ct�� ��G�%Kq��lЛ��'@��^a�A��t=;8{���"L�'�׀W�)��40˶�+����,��sħ#������H�������F�̀��0�FO?<5#���$=���zmr��=?ZY$�YRȦiT뒀m��/W2�|z�~|�@)q!2�Ѭ����y̫���s��a�r��#�2���*�9��(<�l�w�b�e��9>xDë@w$���F��O3Cלk�X�ȗc��!���z�� �K?��=�.I�C�/����
t>���R�c���ȭG��[*BZ������k��n�m�ƒ�pU���Ƚ6MUŁ��/���H�+ �W|أ���
���S-[����<20�(�[��0fi/�O�=���8��C���8;%�D��^�}���ة�k��M�:���!�^���h��Po�B�����L(���!��h)T����`�&ި����T}�O��Lq��6^�c�O��3LoG�2����+:nOdY���
�!��ܖ�;U���%S_��X�g��kp1Z֗o��^O�56�7>~�:��}c�bM2'_��A ���g&jOe5����#��&x�Z�oXD��Ўaw��זf������љK���`*��#N`��lC%���Q�r�;[QN%��q3��$f5P_�<aظ%��PP͗�J�����$�绚`��/�8�W����Qw7Y@ǆHl K�}2�֪��o�����rg���1����5�m���)�`�B���!p,������(���q?�g��"W��ס2l��(�s0d�s�t
p�h��b�G�0�U�ޒج���v���Y��Ό�T��?�ݘ�Y��y�w�H���簑�Ժ�v�yM���*��h�����[W$�X�+!H��3���'����l7(��0�IA�g�Lr��	��"8C��$����F�2|�]hX��sYy>j}0{ۃv۫	k0�"^z�	��GhGI��~�]�Q�Cņ`}�L�1&'�T���S�%q�R��e�ݚF����5�c�Ws,_�{_���K�y6K�Ay�]��2|��8J���y՞uJ�r�Ɠ�!���9��������@��ם���!���cW����g��<S�#���(��l��l��i���.��`�t[-�T�k�P�G��[���!G�+(e���="�j���Q�l�1�?������)l׿E�ŏ*~u,�YW|�V�*>(n� ��JG��5�6$���ń}��	��2(���p|�2;���Ȓ�i�;��loN�����Q�C۟�3����+ϣ�`n�h��K=�����2�e*/�e��C�Y����F���{wg"!�>� u�l�db��C���o�$��tM�X�� &{i�Z�#�p��+�S���ͯ�́�����;��f����>@9��*&~>#(!�	�����*,��ڟ6sr" ��5�P���G����
���A�	R-[�ٯ�S�pN��%�̑O.�]��U�`gҕ@�x��)TKv�H�<��luf�����i�x����z��X�XçDÜJ�wھ��D],_���o���_,�j����{��]���ړ>��M�0�M���e�I��ή���&�TV�"�4�%.�b�X�r\y�@�bL�������h;8�)����I�A/�=U�3��l�ǚ���i]����꩙�iHR��1�K�j]��'̅���;��+c�]L�D��G��&X"4��]�2B�i�di^j'W����IY#�T�U2`�C,ݢ�Q��ͱ��'_�,�Med�g���uԿ)��K��C�
,�u�����Y�����\$�j��o����k"�@�2���؍���@}[?h�̳ʣ����h�*�O8͵�_O����U���_]��4A��_�A����eu�s^4�2�˯u�^Ȝ���l¦w �J
����ZY��J�ɭ���%&$�/p���������9�Hk���[���؉i�%�ǝ��/��)!NK<�Z��X���y��)J�N�����;?iR��d����0�^��e���%
��?M�n'C,R�h1�n�ta����B
���p��P�|\�	��A\�'_D�@�ܝDM��׃&��w����"�νm��B�\n��~��T�m��Z��nsr�0[x�E���U�*��0Ց �mPyJ �p[��sf��þ9���b���Ο/���^NX����8wr,]��s1q㤥N��Z^"�e_RW�@}8�g�c���h������)ԣ�>;�ߔ��x͋0�s	���[�ء�`�K�6��bP><�Ug	80f�����-��UHA~�NG�B���=��[D3����* ��]����[�)�j���?���g�*<�7#�:��p����t'`K�Ix�x���HE��3��C@��	YC,Y֧���AE�\�/�
إ�ڃfė9K�l���*BhW�z�v����Ii�?�ٯ)\��%'<���Us�t�n�����J䁄����p��XT��P�����|{�KP�XΙ�gDN�lt�ZT�XW��k.^��@��2�86^�_�4-��n����`��n�~��}P�}�(����
i>�GA^#d����+�u�}uh�E�$���M�\�Î�U�i(��jD>�1�J�{�*g��ߏj��<��eJm�V��f;;��̟��e.t���	�lW�Im�U��[(�sa�	|�i�z��g5���Qס��J`w��YG�}tE�ra���f؊�횓I/��.��te�	�?�Y����k��tr����c4��	�m�������]�UN�ȿZ���G���S��D�"��a�f��s�cu"�jq;�3�7�	�3��=�=S�Ԩ���J���� |��}w�3��w�RLP���U�?@_2�m%�é#;o�P,�M^ʁBX�l��z�˧�8�xiA�bj���_�"x+���~t���{f^��aIn��;�9#�����N���^9W��<�t�S(<Pg_cy�Ȓ笀�l���9|��eܷ]��U(�M��~��
rV��hg��'mOb=MF[w�Đ���p*D1��3,kn���{��4�76����`�j�Fa+:�@@���aݹg"K��u��x�n��yi��E�$������ms��㗥� �'�I^"&��gL�}��#	g69
�,@l�:L�~�?ܕ:��z�X���C�&��(\e�����8ܐ+�G	�~T0�F���+rm���a���rX�S!�ND[��}�q|��t"���':/ǰ��\ՖwG�������c�$�L����b� rG/��@c{�����31noUϺ�u��B_ř]�2�	�WC/�-�����G'^ f0c�MB0E|�\��Wg���h����#�n���+�5���Z%���
��N\Q����R�W��d�+B�Z��	U��Rj\kЎ4��g���H�UZ�A����g�Z��o���X���|i�8�?J����>�8�86V*��>�Pd�p(�Z:�Ca Ò�A�1���=��\�m�%�0���6`b%�-�c��~�R��t6���/�N�ڻ���:�&O�p��
�L ����Y��rE<G�f֋G�alr�g��/cݓ���ɱc�K�n!7;�w���'�ɕ׶L�����N��Ѹk ��x�ʓJ ��w|.�wO�?����K&6JK��6��&��	���`�(�}p\��p����fC��%#��	c��Ǖuh���-6ds*�4=�ցZIe�+�Ӌ�7Tc(F��_8�P�O3���E!d0�WP��d�� J겮^��.���Ay@��H�ŰN��BZww	U�>��云��S_M�U��!E��F��\i�^��,��H��\�ql���g�K�_⭩���8�8�.i{��Xք���o�l��ޫ�c�pʡ�*��
[se�A��i�A�m�e
̷���'N�ğQX[���i8�R��~���aA��!�}:�R�+�·;*-}�/���h`ӘQ����l/�>>�1��o�