��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�!��
��%Y l�׾����|R�b�@�n�?O$��5��z.@�ڴF�.�ʇ�t���%Sp��f�/�c�~.�ZI`��}�\�x�cr���r$���g��U���\��x>ٍ�\����{��D�<6�9���V
�r�_�e��a���)�'�����F>V�Sx�D?��âG��OX2�e!�G�~�DwH���� d�qu�>檸�� �I�k���0�i�h�~y��I���z3��X�<.׬%G���!���7���( �n#�N"FX�S�+��� �P�E���P]D�
nx�?�s��A�e�����=���Mwv�ʠ�"�e-�qӍ�r���	j&���0N�jNr���"8���ͱ�\0��\��c�{vY�B���$굸�T�٦�Y���5s���O����V�z�� h�6�����>�����%�#kό�0d���cT�;-_�#vV
2~�����ɧ�婔U�hV3�.�:���Q�.��4��׆��Йe>�3`��KA��a��$�K�J�v�!ui�R��4@�D>5�m���ef�Uޝ��_~����('S�B���3��޺�gH$�-"8�|������O��9�fD1�����v�s�^�d����!�S��ַ+�Ēo4G�ҏ��}������{�FZ�[\�;��Zw㗁�d�\w����?�s�To�3�i;����J���p� ��+v���{4�@�*��IP)�rS�8\ס�����<�	�	B��9xC��A��;<Ӥh�6������n�����x�9㹫u�3M�2�\��[���=��fќa
�i��@��G J��
3��ܺ�K��x�p�	v������C��͜2\M�±�	/��<\�U�X����� N�a�ͩn���D;���]�Bn?ȂiT��/tK��i���E�<XGs����<7o*�U�k���5C���kp�`4I�@��M��u����W�E@���o#'�k�hu����t{J*/΁����6k�Iak��*���4wU�	vձ�*��f���_��浻���}Ɛ:uTt�K�ee�������cn8 O�:�������}�y�t��q��yB���t��m(�5;N[0t%0��gWi��^���1�O3HR����&4[��"����AJ$�4:���n���|���l�/2`>	?�p���p����-�L���?1��K�)9�üZ{�]�cˡ�M�HKZ�E�r7|��5��5����ue�#�32C- Hߚ�)`"������_��on
n����?`?2h2��㼬��7#,��7Dsƣ�b�_h�~Oc�2�h�b!�����a���*ц�� �����˽71cM]_�P�./�T�?YO9*��:y;!��sh�j��$�����'�:���TDm~$e��5o�τ9(�l�=�"3{$��i���Gժ'N�W(`Q�B��ф.쩙��Z�7�I@m�:��a�[f�C$B�s'��9\��V��@b&O�b&���lN
���A�;�Ϲ��-񁐝~]F�^OI���9�!?��]��]�������,K�痊`��Ovo+����MFS�U5±��s�$�;*���u#��a�O1N�3g��H�/�	h�N���g��ʪ��r��q��0tQ��	��2O�vg�Q��]�`�t�|�h�:�����ɠ'�u�~�w6��T��c�%;�]YAxJ��<Sr�e3w����	9c���2�av$\^����R���C�i-�t^�;@���6�r:����r�<��pN�im֨��NqN��J��g�!S�l�Ȯ�7�KȓzǙ�P�M��/�{ˈof��1=m?`T�3O����%��m�^�5�D�����` ��]+�Z%�M�Ke �L�39����t���K_�/�1bKhK�0�	>�>�TBp\F��H�[�ê���HAz�,����$��o��5ؔ��7����lN(���&WAR���iH�8oM�쐱�/V�n-���CW��g
Q�)
�;^�x��2u�g}$�kڳQlC�Y�2>�_r�)�d��$����3f� R&����N y�z��[Lbf����)RX]*O���D��=m�G�^���;�	���G	��3�]�&���^�}TMp�|N�	��,��?D���3j����cZf�SI������m̝ZLx���ZG�����Fl�\}L��ܚB�o+g��Zlcj�Oe���9�{�N���:�! �����v;���@�m�x����&�f�rK=��봈D��} ��� s=z*����ʂ�;N'�ق�N�Z����U(*p�xm��4Oxqv�-0�;�N 0K��'��+����|0~��H�vb��E_�����i�[�S�et��{`�,��1�1>O'Ĺ{>[+��B�ҏ��
�S |[<`�|H#
�r
��q�E6&�c6�(,��,?p�|Q�/�|�;��*�y����bBR	��
�5���	�d|���{��*b��]�(�'���Qdy�{�S�y!�$Pנ-Grlё?��+���9zlC������C!EۋY���������c�Z����{����m4&��W�X�	�܃�bLA�Ѡ����7��7�-``��?󪁜a@̻;UV�U���G����d�Ob�?g;h\; l�*q�[s_��aX��w�	�xn����h�mC�`�p�V����>�eA�#q+��3��t%�+f��d[3����ac�Ęm�@�P�鎀3c ět(}e�~uN�,����\L��`|�����6@pb�+�����%e���9��:���>1�G�X���V�Z��XY`�*�)�G���Fd�	Z�!k�M����i�� �K^���@x�om�/����ʼ�śuˑXFr+2�U_u����R"�)3҄��-.>��{�1WH�3-���=���l.�x�Ib ����G�ˊm69���3g�~��P���$�d�\% ��T�����J�P6����������a����^p��f���G,5��K?b�WɪL�4\��:�Q�0V~V<����ɧe	��M��;� ��x>:���_�7�{�[�l�GQ�ѾҖݬ��`*O�Q�}W��o9�z�h'Ϻ��v@���t7t�4ˢ����u�c˰��T��-dcBҚ x#Mr*�ʂ���M�5��:]"��eH�n��.q�$=.0jԫ��|�f����v88W�o���D�)��Ӌ������ZX(�4<dv/��Q��P�ӣ��AKF���Q��z	�l	i"+T�b�o��x��<�cv%��ۭT��M�8<8	��l� �*u�