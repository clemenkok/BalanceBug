��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d���麍�Ks�%$����+d7��/��������ߔ,���<�E�]��&��z>��>�X������,�){0����E�̾�?�%xJ�̈́1�C,�S��u���7�fBCR=���pE��䠏��Lxwʼ�o��p^�1n���d?v".O�l5g�'����4�Uo����7�5G��Ξ@��/6����=;+�Cgt�ܫ����ߥo��yqa�ĝ!�G�F#{5� �E؃��\il����A�E�sƸ��]��i��Y���i���	��'i�6�9U�x� ��n���}FA3.n^�^�ʠvj��)n)�FPF.�UԹuFy�,�;䋜%�1�F,n��{�v���Q�|/'������Ԛq>4�	h<��9�=��3a�G@;.�vt� ��(�/aM�S�� sX�� j֕�������W��_���� ܹ��uD����W�բ������_o�io�&*y�̀ɜףqK�TN�y�G���Q��No�������X�K�Q,�������)��;"%ܱw�H��$u�	C"�Ʊom^k���=�)[ZyY)�����ĚLI�M�ײo��k&Oc	�����A��6Ua�x�V�H��po������\a�-����O���u��o�W�������G2���{@N%w@� ���u�0v���׋�/���P�z�0~� "DKH��h�I-�1�ŀ�ϸ���`%��th��O|�K8����Ct%�o\�����<&g^�aZ�r8v��߯.۞�=����_
����斛���k��e��8{�l�.k��~���)G����~�lcd�aR/��F����Xa9գJR����8�FC$���̰������ɰ	���s���?u�Ǌ�dq�X��ro����AaZ�l���x�%_��XA�� ���HR��d�͛3��c�i�؆�}g�8�� ��B��	,w�A�n��5�:|����R����L��eރ ���EgY�D���"�H���L��rR4�:��y\�S�fxމ��3y���
c�h�������h�#4~�[�wB�CAh�j��2�������aq���>�Ã�l.�������*�6hԤ�t���Zh0pɫR]�]	���fmt[�ʆ#H���4ei�U�2V%0b�I��K�����2�4kP\�}f�MWސ�j���3�Iϱ���4�Al*W�����L�ͩj0U���o��y�6d�Rc�t&m�X����+Ŝ냡��}��i�D�ŧ�[�}��e/����a�j�MX�Ĭ�9;��G�v+G��`^��iꇎ��oTA>��:�m�r�NÐ6i��${�C�J;��?P��V��`R�<uQE��7R����ߌ��>[���,�Aִv�W*�&�
Qh�Hk��{t�p�
��Z�,�����@���E�ݪ�N��UQ��͍q��3����&�/�$�Z���/�v����	�� ��q�������B�}m��*
zkx$KN���S�ziM�H���.��i�qQ:p����N"����y�M
�D	r�1$�ĉ8�SA�1�J+�-f"h$x�y�����{" ���5su��Ν�����՗	K�v\�`g�=�$7BDfI��%�EѐTYÝ�0N4�G��0���y�A%���Z�[�L�:�W��,	�V��kSrΫRo���'���[=��]f�<��r����l��g��V2�f�|�_��3�bص��G�Ǭ��ϫ�4`�z\9T�B��X]A�.�����N��s$��
w-�E�$������R'_��)j�3)�������p�>Q�"��� �o�Ţ��MH�FFb̸�B߮]�Q�T������5���ſ�9�7�͡}Tu�!��
5���
��+a��W���7ζ|�ڧD�K@G8|D�8*�9ʊ�yޟ�֧ϔ\US�5�R)JV*3$�,R�%3�s�T?��C���T�������t���hdۍ��N�����#_i��Մ�����X�b��d�T��@��3{^zz��	��|��j�=P>�n">��MJ���i�C^*\!�p�x&wAJH�HĬ����z`�N4�G�Ub`A{��뼧_p˟�XS�0z�٪��\m  믵�Msa*�q���v�r�mK�������e�ܝUw<k�c;{�1��K|?��v����!'!���:��8�	m�9�
���mB��ҊJ��ߟT�
��ۨn�sU�~a�h��||_]�5����S{g�I,�����/Tl�J���ʆ���
�U���Fh�d3Is<�oJ�Z����_O%#�g2�D�UJ)���p�����T�=����o>�����֋��LV�c�m�4��lص����Ȅ�Ĩ��Iy�I�v�������Vp7ط���DH� ��)�]��Ւ�(�j�����\NW|�dt.���X9�ev��
	�h���A=�ɡy�c�R�ou� WO�,�:�([��e�uxDˈ�;��~#��L�bB��D��&-������P����������z,9�P��0X��������!r�󫹀$�q��dVh�U���`f�B���V�n�SAP�$�^�pu�bX.�c`��W�د�Cn�"�֞?�{�y%k~����("V�|uG�s!4&O�-Y"��:�:R���/e�Fn�Dz�N���<3�5��뇋�,T��]���+%;��/H�l��.,˕v��fz=�=׉@!�:p/�6��n�����׍3�}�|�d�`t���7R��6q�H ��E_�_�����}�f}�Q�M,5�,g�v��	� 80s��kM�����a��jPB�����O�������>d���n�XȂ���y:��Ng��c�1Tel"��4]����s��S8���7C�R.,ԣ��G�z�6F�Gx���\�pB^�S2�b�=Q���/nG��'�'<\~�J�DK&3�L9���6��K���$>VI��+\e�@�Z��kB�Jy6�j�S��s�ǨWa����ˠ���q$�O*�~�ҵi����a&�O�R�U���t���;~� ��N$Nn�Hm�*f�w�����V�ߌRy�(��U{�� ��܄9X��x�$R����DoR0�.�{���l6�h�q��������]�unC�� C)d1���m��o�)�\�v�v�q�G���S��@��77�����/���v�s�#4��-�l��7�1�;R����`�����$����ю���Y�?!{�z���U8�q���/���#a�)&<�7�e��ƭ|n���F��VN��T:�g��s'\\����|I�,�Gi/�ճ��J�G�PkO��XnB�������! ����Ҏ�?�=gȬL�[Y���3%�Չ��x-��"}�r۳z� ާ��X'�bM�y�P:�����"���^r�qg����F�Ċ)5ęH�}ze3eib75�b�Y�̬�����i�=U�|�5���U�L'J��Yu�xB�nc��AA<�J����]�XNk��U!a��l\3�*"�F���;��E�:NɏoF�I��ϗ��cˮ���G�N[�3������\�g�m�X�F������=�/j�U�̓0������p=3��a��Ը��w򳉲��%S��w������\�>
A�ۆ�61�%H�6�)-%2��w��le6rW��]�v�˜�'ز
tNܖM,%�� U"(�w��T�PzVp}��{i�4g��:к�-�[��c~6Rf7��(�:�_�Ȼ/S))�g�]c�v�<����6E�,8Q�_o�!�&nO*��i�sehp3�,8r0�Y{aj��:H���`���vs��	{V�w�5^���H�|��X�VJxD�.��*J�K�����'�7�V��<�,�ʑ�
���4IU�@S�����'Ko�]��FE�%#.�@���TY�rO{66V�\{&v��r�`�]Ýk��>�xjJ��-r>#����b�ex��V�8�j�Ig{��៰'
9|�SpBн�n<D5�hʿ����ʽ�<eܜ{�ZC ]M�ľ��(���2�ջ5��}��'.[1�U7����џ�f
zVN��YO�����vLJA�=0������а���0Ԣsk���V��zG��s�k��ov4����W��:�"�'��$�*�NVw3z.ޟ(|�W����8Dt���r��k�M*π��La]�]RI㲻�����>P�p
����ڱn�W7{B����M\�?3���5\��Q -�k׍)��C#aX:R�9�Ib+Ȧ�mtl����x�=q"O��lZ�q�7�=j��hC9f7�<��o�=:Y$�hʬP���z<��_��V��+�C��������MW�?�c�0��-�i�d˗��Z�f�jf�}��9�j���Z9%�x����g����5�W�9>�Ui����@{OhlG��;f���E�`��i�hb3U���է����:��ك�O��+�L������
�|, hYe���Qa���WEf`<�B~CP�<�������.J�~�/����9�T��a攏��P��m����u�ng>�}g��C���,Ŵ���~�O�j��b'��D�J���I�g��M-8�PASPk�P���	�nE�&�[�U��}��p�Q�(C'�I����m�xwl��d���������:;���"V��ku�E���H�G�ȸv9�{@L_!/C����z�
�!6� �!Z�q�E�W�����)rC���,o���D�i�P��}ʘ��=��u��Mz�y��Dm"Q����C�N��@�]�3�X���H�\e�pC��l�~��:�.��55w���=^��п�`}��:>Q#J�$F�gu�-�B0���S�+�J��	!,L�.X0��t|�����L۪M]�~:E�;��%�qH�zLe �|����!�ѽ��^r��Ld:u��� ��a㚰�T�嗌Ħ2��j)��n\r$��2l�&���R�ui$=�E&+U'�"I���n��h*L��2��4`{M6Q�S��AӚ�>[#�H�蠁 �[4��Rx,�޽��2Gs���ey�Ew�8����	2#ͣO�A�Ƒ�!F8��:���]f3��x����q�C�5N���?�sT�̺u5kߚ�e�[��<׆Y�FS�1HgRҌ��:k[%q�ު�^a� ������M,��!V��?M����_:A1Wg�5�h<�N٩�;/�щ�&G�c��;p;)̐b���s�u�±=%`%;��	��}[,Ns�FU1/���f{�Tx�N�%��N\Y���Ӗ�)�w�h\63bk�	ؿ֪4�A�P����F�Ճ��z���9B
-ύ���l�	�*,�#|�!�ooW&`B]A��.��[����:dn�6�(ʵ�<��嗁/,�ۢd��!�Om%x\�id�����Y�)�ރ=��G����4��v�S��r����1ʮi�Yٔ6~�A�˩#뇽����N�M�3wi_�شx���$d���ԇ%~��7�g�[;Z��2T����SS�����̚G�ø��$��L����'�y?-�o���9 �:�
������
_2q����58����S��!A�=��e)�ҍ�EBm����3��3��R8L��%�QQq
l�c�uR���;��X���Ή�߲�������t�H�2�A�4�c����Oc�v�"��b&`W&^F$�@n]�2À�Q
�9�ӋOF1ﺴ-���@�NF8�=��t����+���,����G���s������'��2|߶�0���y��� b�bS�� �$�0Y���P��qxH������\ϣ�b!�S��i��(0܁ױ�d�d���%w�����lA�����fѻ3.�[�Hq��������xPc��m���e�4�ΰX���/����ߠ�jY9꼄�"��![vb��T(_�TYs��%����b�n���\{��h��}��&����ȜzS�䙷5j�"���قj�f��5���U[�Ij����V*Ui����.!J�[^"umd+�=�tUnFZ��=@�߀��DY!T񷅏�M���.��w�[��Q%�5L�֚����S���	�o�|�@�����)��|s���GC�����t��6L_Y�A'��[�O�B�&Fݬh�(���
 6g�:]#Ż}���T��e�.�/�&��w��uT	-	���4���t���H�K=�r* XءhP��gs��_~oRűE��Æ����"�'6���Y�tSe�_0���+�C�U7��"=�tV�ٔDx�$�gˀ��3�姢��$i�l�=p�Lx�����48p���&ă�a@��/�~:���	7�E�%.�����l��B���<r�B\��bɡ��a��(��4�f�1~	�s�6;f)P�&`B,��n�v�s�mnàV>n�j�1�7�0�I����w%&�Ml!�!��ċ;���I�>�q�JI�2�6&��=�E�����P>0تu�!�F�h�?�;)5���MMy��3\5��tʦA��N�����`5�Nx�.C(��	՗���-��Gmi,^x~�˰(���/Y�4P��`|H9��M!E1o�M������������&c+q;ZmI��(f\i~�G��bJr�@�7����ś��Md�켉�|�7 ����|����G|;��uF_�)j�T(F���q��9OKǱe�_	(���g	r�7�ޥ�N�p�2�bE��,=���J+�q)!\�.�?攉�5}>x�/8~�ظ���e@q�Y�I�@?Evl�w(6��I���yޛ#��X���'�.�$��%���
�N�Z��'1�f�i�f�5�Yp,�u�;U�-�;�9�
,��-�=���&��ȝ�%��C���L	�?D�2�Rve	f����;0��^:�-�(�w"����ҩ��.�{Y�5�/�?z��_���b�%�fLn� ]�6���c�E5���-�A ��x�S���HcՍ_�U��m_��Dy�y�<�h��� �v�����Drd?EmM0:����S�I|��H!Io��N�i�H�/Z(T�^ |��WB��]�!|k���W*��h�f�����p���i�FG��c@yN�	UXL�#��ՍGr��G�$�vo%n���������!������i!�7�z�^��;-'7�ev�:]�I���r��8#J�)����N�--�kLt��� #-�H&��?*UE5����;����u�:�yT�|�or�����V٧VԢE0��*��o_����N��	�Q�B�өma�|Jf���s�*?&>�v����y}�fH�E:(�מv$ԝ��c���v����\e?F�a#��&�M�q.g���s
dޞo�m�,��A��Ԣ��^0�ݟ���F@��Rb��&_&�?;-;e�/6ר�z�M���k��r�}��gr���:W�*�m���x8�󛚠M���j`<� �3�����C�;:b0С^x���������#;ۨ2�r\�S�Ӎ��M��˄��̷إ5�|�GLx5X�C�Sf��� ���v��U�����!<.i��I���@�nN���i?E*��i�;�Pk��q@�$d�n=J�.lQ/5V�~�V�U�`D V�j���wٷ�4"�M�9��Z^�A.0���c����n�m5%��=T��o�1߁�9-m��#��� ��2 ���������ka�K�ظ���3dD������� ^��+�*#�Ł޴�k�xs�p����:N�*>8Ͳ��hsy/��m:�I����!r7XiY+x� 5x��P��/#��*�̧_��(7���&�D~�>�U����ŉԜwB�"��Nq�13���y7X]��X?���>Y���A���X#�k*����	�7�y��4�3{:�yEaL�?bD^ÔaXx�����Y�Y�+�'jݍ5��]'�m������v(�h���$ҭ��-�s �_�{��b��,Y�x�Ўﳕ�H�6�`RK��XW��:��*���(l@@�4�)�	����}*wi{"��ڹ&�V�'#a�7x�k5wd,r ��0BP=5�m�����>G=t��1ɺ"�ڔG����\u#�%�@��_��ߵ�Y�Y�-�y��)L+4/����[�܎��6d�W�UG��݀�lkmd �*�c_9�L?��6���f���cQ����g�l�ƫ�Z���hD���M1KB9���nh��H�N}�ϐLyh�ar�%"�J��s�J�:e�����0�K��l��~W�TRўPU��
��	ՎΣ�K�=?�z��ܙ��p�LK���a��EA�q��Iz��cTk-7G4-_�xY�BN�>>�UO
�8��t�R����/AI���	`���9��nZsd���S����)����`��@�Q.�c�*y1p�!JDej�uv�L�aE4���)`��?kD�[���Ԁ&������"���K��um�M8����Y�y �����[�O�ܠ y����� ٙ��%�2o��s� �o+[�jY9�{�H����lTގ��#�9���C�����uܾ�:�Em+�[� ��$��XF\s��G�8�����ͭ�9䮎����F�yٞ�����WL��]����5m0>���������l.�#�w�����\�B�.�-�7T]J�gj�JR��m��]"wxlh����7R������:��Z@�[WuzdH���wmA�0�*D��Ün2�7L�>j�N�^�2u�h���Hvr�?g[�f�(d�{x�NTã�?U����{� ��􋅬piWηz)�eZ�>ʓ���6w"Ƕ�y��e�B=C����-w��Å��f5��x	����`lfy�����XRU�����v���iE�{�Q�w��	9Yk�~�}-�˪��&/S��:""���=�^��pH}}��qw`�z����*��g^^�,�+j���c��A��_����v�'&��N�$p�_�G�R(aJ��8<����Xw&���������Ȓ�/�ݱ��
�B;��f+��2>'{���|L� ؼ>FԚj���s�<�{��L�H8 �-\<U���Aԫή�Nv�6���+�6	+�ii��ל�s�^*�M���M��d4l�eczg�r����Ƚ���*��ryNF��&�A�=|ɕ�(�!���4��o��A�����}Zo�NA)�2p��(j�f2M����9���\l�a���83(p�{d���7z��`<H9�th�j,�+����@�����bQ��'���j"��|D����^�{`G�D�ަ�Y/Mj0 ���_�T�Yk���(���n����5����ܫK�(�ђ���\L�eW�|�G�d�KjjNU�u�Ӫ�"�;�mQ�F**���cԌ�NG��˴��H38���#F3R��3YH�:q�����b/�f�w6�=��P�N�ל������I4��  l�0�?zI �mq�DoDz�5fzE��l�2��\�|6	C=
&�<bl��s�D�<J�����A�a��h{d���`!�)��p���$bLx�E���2Tkv���I��떬2'���T��$[����M�
��9��/�r=�ǲ�c��8d�^�V�H�+^��*�;���̷7qGc�d�Q� ������V����<�!��-�N��n��ev��O�+�C�{V6�<y"�)�C�l���I/䰁�uE't«q�C����0�9��~���56�����W<��X���%=/0/U��-npx��4�+�w8��y`� J��X��ηf����z�����0d���U�9D�Oj^E�Aj���?�kAn�kRE�����u�������M��F�f��E\+vA
L�������<eh�KcˮZ�|�5#�ױbD��д�T9kL)x�����
H��!^L�Dp?��\<��pA��
� X�-��k.T;�wBQ/Аq��c��j5rYS$�6䫉�M�Ƙ�7�uT�O����īTXվV��Vt��;�Y0�h˽�?���Kzu�I���̦��W�h�H|`!�U��ˈ,�NQ�_x��z��W�_���N��'�ul7U�	�RR�_z���K�2�};�XR����dp 9��W����q�4�q;�_�����F�Nԁ��&��͉�Vdt�]�<�U���0#���3\3C�l�R�_��;�0+YG��ɶ[��p�t:?�C�A팢�.��2�c����?����T�/��n�{f�ϣ�� �Hb�3��hU��lB��rc�7�@��.��������Dyw��'D����\,�Փ��	�9�#%%���o��5RZ�=]��F{"�D�]�_K��ϭ?9�|�p%Ƣ2Z�mz^���v��|m�Y����
 ���$�,��i��� ���-��7R6����|x?ɇx�w
Ee�7�ّ���7s�����<g���u�i�~I�_j��^�!�ֱ�0yRf�D��a��P
Ӣ�f�l��H��ar!BN�􂦷���VJ�\`���ȿ���V��w�ȯCu���6A=���JL��2�ek	���:�j��X�f��s�*���	�Eo�A�^P�t�wY��$2\4�mD�&�_8�KJ͋�-E��ԑ@j̭�ާ�nw��h�v��B�;�X�j�:(��bD6�FA�ǽ���qM�SA�2ƪ8%�M��ڟ��?�J��Ns����$��k���(�q-����p�����^qE�F^�tS�L�ד%������Ԓ5�5 B����G:(k��U�(a{��kJ��ERe_(d�y��C�������p�8OW�	c�QFm6���,'I��*���Y\�{�xJ)�V�H7���r"q�5��&P/g�<b9/���b&B��<|�2)ݬ�dr�8Tx��{I��BaM%f��^nf��XY�D��
��0���Z̄9�Px]N6�a�k�RO?g�I�ܐ�,Wd��MO�;G�U����**�������"��v��6���o����Ui�9�;���*06nf7EY���v+���F�����S��<��<�Ҫ2a��e-'�2�v��#�`�{/�R��6H<�jI(݃�W,1#	xe�U2~��A��V�j
L����XOe83�u��Î%--��:��5��1<
6��FK|��5���v�260#��n:��ȿ�FB���d�ê�i�3�cT�l}�����wl֏@��O���Lx
�n+�C��3 �����������:�P�}�.�M���Tcl�D�X݇=$3m29{"uEZ�F�iJ��*g?n�s���Մ�(��A�Hucb9�qǏP��O�����Bя�e����Ok�M��U)f~B�\0����_4T�0K
�c�Ti���C{�@9���%��.c��WN8��gj��!8����v|��M�F��������%M����=35���X�~���t6�uU��I������݆3q*�-0B�N&�0��/fv��^3M/*�L�"���̠����/�֬2�������%��%�!))�ٕD2Qa��Zי=�7\I�l�?���:y�Y��u������g��?��#���;�U�>���35Ue�iY�>ȧɲ��6(y3�I�.Հ�:*����fƞU[y�W�z�>(�4!Ԋ���u���ʳ���{Jyfo�&٭2= �Z��xiI��ԗUf��zB�W�	�5R�Z7���ĕ^��g��&	Oѵv�&�a;љ�~ƨ�ܻ�AL��({>Gf��яx�歍/
���}��4�u�_�`��J7��f��cq��nW�ĝ�ؙ���~���@z�{��V��G4�.�����َG������Z��,����!��%��R�7f��I���c�bюyͪ���i���[ez�ɮ�̔/tyT��ʭOhw�E'ib�v�.~����%�Ɏ��̴xZ�"xڂ����hj�x٨�l>W�X���/�7_nA�%�ŉ)�II��h���#�� d�� >��3NA��J�8�Hf����ܞ]�3���f����G�9R� �LE7��˗?Μ&�BSX	5��ͣUc�X��(B9]O+��y؊}G۩��Y���@z�{(Eu���������\���ϛ�vĻ�*���-X��������lL*tz���R��46_��1XٚQM8���]���&��laԹ�u��F?��K;�P����(�F�C��3�����.X���ڵE�	��5�����~��N�/��~��� d�*���b��4�&(H��6N��2),J�I鴾�B�"��D���ۚC�-��*���I��L��{O�$3���A�&ʦ:�@_��W�wH/�$��N܃��yv�������1�p~��ʝ�fpB}
�����0w�T>����*�c��d�o�aG��� �*2g�@o�$�w�6@���p`�j^�ʡ\�4���5
��W��(G��y��~��T{'{H�>���ᩦhOv�������l�3��,w��^���\V�5p�e���P�b����(��IE�lw����:��p����ޘd����f�?�c.�[�VӖWN/���N""��E�ڂ1[=��m��9it�%����\�g�n=�l!N{���y�T�ΉY�Χ_���?�ʪ�ʓe��N�'��I�9׼��S�-@%/�	,*�-i$EA,�����������w.�Qn�q,����U�mw��Ӂ3�A�B�$�3��`
^�`&c��a��NP��o|�e֙<����Efy���g`�5MdQ��Xg�i�?Q+?��p0r�練��~:@���*á���6�}��z�3$���V^H��8nQ���p��B�����c���_ʉz�}��T����u=��0�<H���Bs��^!>̈́n'%,��s���\t��6i6vba��᭐�=�ٵ����*�ңo�"���U�5����|$X����^�F�����. �Sb��7 O�`�=�FI{Ne�yax�C�U�T����܈���,��l#���{�]�6Bom6����?�-z����RG�������oB��>h���k���<�)�T:L��ⁿ��1�ϵ��пL��p��'Տ���l?�iO���Ε���h��OD�x�[-n0�_�mTH�;r&�.�܅7B)���^�]rCR3X��0V��WNP�NCK-�u��+f�K|?��!�� ��Z�!�0��b$v�.v�d��H!��s�($�0��2)%��iנzn�ҼB����/�Zo�?����}H�$���2�u��1�r ���L��4U�\��u��q�W��
r_#�u֝S��Xs>�z�P8����ֶ�S�5�^�&�/� �Ȃ���27���a�Ӆ���ޟ.�8�]E�
L�#\��2���<�z��'$��_ƠlR}��Ǜ!�&ÀG��	b
�%�q,������G�<���v��ւ�x���ᅂ������aL����G��Jy�B�FLG)\�b�?�2Ś��0�{�X������U�5��hϐ�b��!��{�M�V3:�g�En�n�8���y�%Y�����-t�h��2�dDw��_8G�˅%����[���$Z`��L�������֬G���
�z�����3M��/�lߣ�Áxǆ�v%A�X݄��M��c������#.<��n�S,# A��4�}_��a���U������$ ������h ��Z�J���_�T7�f�a��5+�ұ�d�r)?M�����<������u��>��7��`���T�[I�]��B5���:F���$v�����|� uQLՒ���z��+u�9��x�'�q:3��	�J)��(Z�S/Ă��76� #`�<2�&8 }�E�s����5��9z؛�=����1��e��BE�Ѕ���S�X(�0�2�bn����%{ƿ��ӊl3|�݊b���¾��̂.�$������+3��(xc8b|���%�ES�>���9�����M����L[[8nʦ��:~,���Z١�JALxA/�ԜM�֟z4�����6Y%E�8`�ku�^�O�}�|��T��(�-K$�Oj��	���z�}�,��ڻ��Q��vU|�7���Y��r%���~���eV�vIx� a�\��^F��[b�_iQ� x1�  ����d
�5�n�ҀIu����N�.7V�����V�7�)���T��f݂���1C�3��J����wT:�9)��\��-z�+�g����I�`n���,���z���x�Ϯ$S\���1}{���+=?vV�_iBLT�I�}��I��j�����E��IN~A��m{�e���V;�w���R7�͗;���э�yK�qX-9~b���IG��~�3�H([��+7.���rd����i��1������8j���l��=W(p��V� �@/���Fݧ��³r��]B�t��1�����H`C��Q�=��ͦ�*waȜ.�@��פ��L��c��7.�u���Ɔx����v�7�[�71
L�fL��Z���(�?�q�-����|�Dz�u��P�$��I�4�����lvLq[��?�r�n�q�a��P@�V-2-�)��c8���ؒ4������c!w��}d>��DȂ:˱,z�|9���xg�e'�KD�H�.I����3�8��Y�lڪ�+';�2���Dt�6�}��L���j��q6���n��X#=��z�]�P�>F�$+U�Rf;����c�F�|�z��a���0��X�P�	�=�rj�4#��ƣ�bS,��	=�)ew[C�1Buj��K�W��(Yˍt�l��'ȫ��s?��h"�U�ri�
N�)z1�~r�`{*Y�ʘ�@� @_�����:Q8����J>G��l����G�-��N2��S�0"�����F)�ye'��HL��}vݵ�^[p�"��0۔g7w@Ż��f@i��A:���a�D$�=ł�!�C���j��x��~M�Yj���?�����65߱�2t<��a�˜�fՀԟ�R�%ߍ"�Á�-��X��	���e��f�y�G�v:u�9l8�$�m)�4&ꡳ{I.X���8�;۽iZhx���3l�gIzS��5���v�6�F�eVk�P�`k`�\��B�|X �й�r��퐺����b���QL�sz[�_����M��a�8�z40w_�*}Li���@{%�$6@��� j��ؘoC<��j���-�q��I�'n�+���Œ1z����h����kJ���t�^�73'�#�X����-N\&����<�:�4l�n����-2���~�)�bj�!�ڑ��c-@�D����!�"^���� �p�
��j
ݹ�٬���TM�#��^"E�+�M1��SQ�Gwp�DGhk��	ni�"��m���I4��8w]���̗ I�r�T����f�\=�2�6�t���K��"z���7�+(�m����z=r¯w�t�AJ�2�Y�Tս�b� _X'�[:#��a�t	n��#�5��3Yw�'���X���2�\���g�*�V�"<M'�}�ZcL�7��Y-���'0�\�|�sOv��f��d�c��;�>#@��B� b�;����������TNi��ҞZ�iM��O�.�30����"����y}����Ju\�W����c�����A�h��J|3�H��]�����t6�}S�H�.�& �:��m����_2����"���OICj����R��I�P�w��k}���M,V�rv�'i%���P,�� ��LM{�$��+�4�9	��<B����^�}��}�=���+Ӕ%̞ڭg�2��:ݸ�����^�����ݟ��^+����ҩ&0�]���"q����~�	��U�/�_k0_xF��g<�0?Z볩"%�}�2��_�m�ҷ��%�4���'�p���T����( J [���.v�d/>�k�"����}��dT�b�]����
�����҄=��N%?|���������ȑ+��6)��x��']�M��+�ooDGC�>�{M8|Tq7�Q캳��bEllA����z�n蟝�G�cy)e���������I��u�FU<C�; {
9��!}������k7��/Bv��Y��E蜜�Dy.6�sĦ�>��;��ei�U�@����n��5>F��=��7<��6�)5�X�.0H�/B�Yf
d��� ��vWg�픙�ܰ�3��́������_K�i4�H���B�Ks����n�J����U����;
3ZZ��q�HS��\��$�{濰[���z�����E[9�C�����_����p����ӄ7�^�����C]��,΂���,��=�S���U��%u�W��[6���K��J�*a�mG�֒G�F�7ኩC0aթ���,�>��1D�	��ڊ9�PπL�$@eR��[�+(���"�9��+?����ksN6�@���f�u�<��+Z9���c��w�M;�fK�p"dfv9�wMm� 6�j��E�������k�G��E�:E�^��|��M(<�0x��9Yߩp�إ� �_u�p����hԙU[�=4�$ �i���[��-�-��U�!ROs���=+x���>2�yaI/17Vw9r��E�)5ҽ:C�)������^3�y?���B˗�Q���W�&���&����ŪM�9�:)�����wC��Q��:�e�i�7?R����b��)K��ɷ�8D�=��π�Tk����e!W��{��)�^XgËn�d���]��b#�2�{;c@�>n�+�䊬����Ϲzm�%\��e!}�O���F@XSt�LP��Cmz����e ���
m�YJ��(��b�f�sD+��V)S/��W�d�=�Y��f:H��\	��[�=�"�Mp�����<��)$�����q��vF�-h^����aZr�:��p�u4��b)��h��6w1eƛr�c^J�qo�o�|�Z�j��*i�����}�.�WG���dp��jY�i_@�|Y �7����%]1����\E�����s�vH+<њ�>���a�����+����`�����ܒa��1��H����l��[��r��N��in��r���w��J,�$nF{Y����䬧?֐�ߢK�`aN9�-�t�1���	
0��)���G��g��Y�eX;`�	�:ZRw�����0���L.�`#ۊal�hC9掲6<֤�=��ĩ�ܽG�=�˔Ӟ[UU@�|�{���[�>���wv?���.��>9[4�p�V2��*�:S��ӑ
�Y����v��`���4�=b��5o(_�,�/B� W�E��:��Cn?�l�����y��mH^/R���PUf����[����ʉt�i���!�V��	�_�Qs���(����3%�v��h�{�:���5CG�1iD�p!�_3����0$��s|PA�'�A��?U�^��a��}�ೕtט�}Nb��A�,V'�L�
g��q"��xhM��*%,�u@iF�E�L7Wn���8d&B޴а��5PPv�&���� WT�ma8*���>��C�;��ٞX~���X�{��ij܂=J��T{FPVsWQ(;W|}wu�I|�(����m��q���$����U �NU��ǔ�&�k�~IDY/)a؁���z�����V"VQ��m���giGeM���II=���_��<A��_��W@ ����
��>I%f�n�^~�T��2����}`yۮu9�Z��Mw6���!!�O�ǹZ����U�i�#��lDo�Ჶԕ�3#?J�\�<��F���¥Ejf"Je�9���ݣ�?%lDa��I�L+cC�
������v�#��Td�|I}g��2��&ּ_A���J�g�PL�_����=s�_K V8֥��^Ȟ��Oo���i�8��R����5y��t�xZ66�/�f�Ʀ֗�}ieZnҋ
9̑8�x$P@LA��"K�m��Y�#��TuwεB��Z^S5�P���H��^�3�f�NlM��Ha؏E�N�>e���c�u��-���F��@sl�F$	l$%��]���Z4�@T���Y���v�/��P�ݔb���|t���[��Y��%����:^u烑&�wK6X�����Ѱ�_I�?�w�#LJ�a��Cq+}�����_To�P]LȐ_<5� <~o)s��3ap#�
���G#�,�A��C��'��1��F�:,T2�7j�����:�=+zB%� �os(e�݀s�ȣd�&s-/��	�^]�aIm��?�Z۳���M�(�D;�����cq)�4�0	��-g3]WM�K��g��%3����Ո�s|v�R�A�����e���`l� �#FW��7�a��0�9��?��ӿ+ ��(��*�5�t�	ZJ�A)��bRe�e��{��V��f��E�Wk\�nT�#%���ت����E�r��������4�݌U�~��ɸ�ky,��FqB��/{I2�,����	�4<9���N��{��{Q��p"X�R�s��r��~�0��qbZF��m1����@�B��b��Ŕ��ab&؟��8��MJ#L�Z�R�%����R6�@IW�Q��1W�|�ܐ�lcP�p�����L�H^>gP[��|
o��������g����J�����R�e�z4v�Gܛ��>s'�hE���v_��i��o����1��A���2z�7��'�No�P����
3c��J	k��V�v>���I�;ı�ܯ���z��W�c*dk�9G��Zt����`	az��vG�X���r��y^	y�v2������^ؠs+���5�@]�5��Lݓ=�:����Jn#�,Ɉ;�)����.��|���#&�[�e�:��	�Ws��s��m�����d�i������)�Us�Iۂ�)��'�����(P?%���,a��+"�/_���c��n�Ov;����乕5K�8�����#���M�_� �N�9�W1�?H�z�^(�6s�c,�N��-Y��'�u�a���H�,I��!�M��-��%�㟽-�����4P��M�����:8�<[�^ẕ[�Y
P�L6�c!�|�i2���L.a�i�?�ANe�����P�4Z�����fs�P�\��`�X�	��4Rv&��t����9��a�����g�y/�a3�CZ�]�W�C�,��33Ě��х��k�C�i�#����e �S����_��N���oN4C������ �+i���v6����}!�S��TD�21dv.����74v�)�XÊ�!�0`u���}��d���y�O����A���ק�fe4���`w��	�c�<�
�4���el)��> G�\5��q�-*�ght�m�#��~q�g�v0��f^_E5e�Gño�V���Z`?]�{�!.,�����Y�]=kzt��|�� �^P��^$(��� �pJ�廋��;�ݭFkF�]�Ŵ��������@�
 ���r��|������	�8�X��E�Ol�Cx�1�'d���a�l�4)Hsd�s�&z�%���'����v�b70��ayf�"�RG>3��K�9J?OC)�Ƅ����!-^�PE�����������k��c+�*x�e�b.���z
O�Q�l�ڍY_�cNb������7g�TW&��zO��]�$"UZ�*�1QL�5f��'}H�۷�k����b3��R�5>���6��Sʔ�,�U8_��&�V���Қ7�b2�;&L\��N:�R^��
�~���>b������YG��2d�[p/�9/�p��P���qZ�I���Њ��}��3���u�M3��$P2���	�AV���n��i�[�1�=v��J��&������C����0�J�7<�w�mꇧ��pٰ\�Or�"��Č$N�����Di7�o��Ԩ+k&�2��W�3/K����?�N���wϔ�`X��$+���A�#�3�r+�n�ʅ�����BO��/����^��2��áKU�	ɐwG#��1��)�9�H#������c�.�5��F��/ 5���_U.�0.�A����0�h��b�7l���m��O#����K����#*e��-�C�VQYO����/���O�o��*��
��L~{,���iTX��@:���d�F����_L�xYssp���nm�ccQ���

c�~|�@�lC~t0���;3D|�b�Q����DY�9P�X+���$��uw"9{�&:��\���k [�}�/�U;"_D=y�A�>ǃ
k@�;A��'��g�혏���Z�4�F:y�$~g�:���m�E�v���`?�x��!�-�P`�ۗ��S�~-�7�Ua�'��H�a?�.�!K�m���Vd�@e�D�fjOS�7�7&���N:ݲ{���S��5E��/"����5��n9+P_�s*���qO4T��T/�S���Rm�#�D|�-JD+֞l�� ���8S�$�%�3�~��=�k�bM�6:H�z�1��P��Y
��{鼷�J5QI} yטo"	�I�ɓ z<����#����3�.�U��hkq*�~��CD%#T��>9��������X�v?�t�f.�t��?K2`�ҎDU�� Zb��bG���K�&��K K�Bw�E>����B��s�G>�L�ʗ�foM}�c���TN��zQ-�v�zy�<`�*��C��"�>Iֿ<_?�Q�:sh���(��`勋��?E'��������I�7���ۺ���o[ЪfnX��3I_��	�s#������߼�ה+b;���	�bpRӃxiB=��{��.*..�*���3�;Y3��T.�"҂27��#�H�ʺ�ZI4��l���r%� �Y�!��#۽_��ƨE�`S9.f��~cHY�f.��Iv��Ԥ�(��id���
q3� �O�%��Ӱ݃���8�ǩLu_}d?��qN����b����KM3y��p�T|��Y{���@��ATkU2�l³���a�3n�Ĵj�W-� �ڔ�Lq_H��JS�p]�\<�3s<Ol4)=Z��r'�W]S�?&R�':�4��%�x2b��3�>��3p�ф���i=���<��bH�g�6I�Z3%z\OE'�sl�X?0�,m���hy�4@ ����%�G۟��	���1����L��{�~&,n;�R���&��@	�&� �S�`:y� �� ��-ixs�a[�"��NR�l���靡��*bw���sҚ��|��,X�
Y�L7ҁ��pB-A���ų^b!�s�r��h{�����8��<��Z��j���I��ꇉBj�R�Q���F�6񪶕{d�#�Cc�����1�jP�ݿ��*�0`��}� =�H�aϕi�T�0��N��?p��9:z�Ӱ��gm��v�1��u�����;��������T�V��aT֎R_
-�����F��xK���Z|C=k?�0!����ExF<�W�g,�y����.�
f>�-*w��Y~a3����Q��y���H��W�R�L5�[QY��5�Bi��h'�����-eDǹWf��)<3K��A73'A�ҳ���G}�(U-P����`2k	d��7J�Y�2�h�W�ە]i6Ӯ֣;��k�j�G@�b7��l�sz��d�9���2��@����P^"���Oǜ�h$YIӜlud�I�;C���@��
)d����@d��� �&��|X�^�����K�||-��%�J��y�<;
,m��w�?)������ƾ�<V�aNĎMZ,� �Ds��*���x�j���<=i��_
����}��y�)�F�)�ȧc �t�U�S������[�N���RP���[���YVa������Q����z8�~�U$�-�;�˿�|I��<n2~���`�9����m������o�o��������n�m�[�7�򔐬���
+�Mh�����&�n�&�N�C � 0�����?�_��D@�$Vz��ZLC��΍s��?��`��J�:���*���2��J	��2���~�)^ ��]h�d��<�\�2$�A���C��%  �\#��bl�0�_�u�"��`�S�*�x FECw����La�#_��Wr����q�� �P����I��������[f_nX�����l��5�ui4��OC\��@m��(�3���Bk7�][��|I���5��C��fER��܅�$˷VQ6�A���$�vhUB����Bg���4A38J�i��*�����ߵ;�#��TF2��馝f��{]¸~��FYpO��ɟE�7�J�\N.�v�����E���w�����s�l6� �pR�}ve��Ķ��!3�c�dh��F��[��{钦Y�'x~
��H��b��U�����*=���z�+ф�Gl4�Ye-=W'	��� q��gf��
R�1ᾌi��ݻ�[���Z���^M�l?�7�@e[�%!]��V�v5��]�#��2]�6h$�㚑^�S� ��}|�����fG�����g�KL��0�P�S: �x�>�wY!LtG�À{�����{�Ř���~ ��y'��ʾY��_'�b���F�G��!�\zw�7OXԂ@�cLi�k_	i��E˔Ѳ�/ڠ���@�\ؑ <�w3Ⱥ�?���q���}�4Ί�X��cu&1h"�|�����{�ͬw?�bfz��>�B���f��j Kҷm�w�=)�Upo(��୰\��pU݇%�������>l)�'�@s�i��i�b��k����K1��x-�a��ڍB(7���g���r������*�M}������R:�S�\��{�o��X�XkZ]�u�]x��\�6<G�B�C�4
<�������&�kgll�����=���	|Q�$�L�����?������}�!��gÈZb�	5��;��hNg7t7�{b�:����ͮ�޴{/��C�}u�e����o���-馔�H}�ɡ�������-�]��	N#���_���%�
��E��l~�	?�.���f1K��#���
dW��PJ�n+�n��NuQ�i,
qz!������F�j캀��=/�o�B�V�dF���=�������;gJ��6�s�2!�K�|��:���5���ږDbDbV��ٺu/mո���vk�e+)� �)��]"n__�*Q�8`|4��"y��c܍�]��220�<~��^0���QϭV�;,�ݱ`o�5v#h�@p�[���o��@��G�����G�~5��<é���L���kcM��gBɔf���J`_�࢒�q�$�yb�xH׋�0Ox�#<~��u�9�8	��JF�-ԇ43�}��2������9!���f󰍄�=�/�xz��J6�u ���L�7��EZ�ߞ�W�D�Xz[�sL�]::BQʦ�S�����{p]�v��:�
i�OP��pN���ik�:��DVHH��S7܈l�bn���h���i"��Ih�$=Ey��@��Tn��ɘ�	�)�����v"$O2)�W�T��x�@!�P�@P�HJS
��z�g��OS��K�n4ѱY��nF/`9��OsE��bm�l3�0#��Cu�ϛݒ���u�׏�O��"��q�k8L:��nꋪu�-�a�$ ��
�7|���$�Dǯw��%v���Z�w3��G<0���c(�����':
��6G����f���蝹G�,��5z�g*^|�*���T��<jU�������qkp��s�?g���8��莢�y��-E7�3{U���iG��p�HYj��f\���h�<&���b����L��8����*�K�a������;�;dk��N݊���YU;�"��&�\���6���K�Ǿ�����TQo�i�R������>�(�C��K����ؼ�c��΢0j)Z0p��.Ө��`���;^ޱtTdw�����'} �ضf;����xΟ~~�]w�A��F�U�u�ɷ@�/bM�!)ӏ��A��d��*?%"��!A�#&�����͹�V���	b?�b��%F�^N\&o�#�<�S�U�~���K��)	F�S����L��ע�x>��'�0��G�N�"�҅�OX�q�&$��}0"�Ц��g�@��!���-ـb핟�#�)D�:K&g���\`�Ωy�<8�w���]�����ʒ���v��m�����?G�W�R�f�H?����)"s�a�͘:�(4�H�&�+�\$/;����ۣ�#\��	G��T�>>�,�F	V�� �,n�RAp6��W��?���8��KLR�h�RM)�m#_*�/�j�>dG܃Cߣ|���9�������Q��D���ً2�����~i��Q��r��3[��+���Umm�)}���F�G@^��=��ql�ȱ�Y��1/@��� ��*�~G�@���l'?�b�KgG�D:q�Fb�f#.U/�TJ��B��|��O��������ɉU������<����	�C%ӈWqz��KT_�ō�=�_U5���I&��q���Nf3x$�Źj؊�R"(���
�&�����m�Yk��H�e��(��~�(�W�r�����	9u�s��ˮ�×��QԣRL�� *����s6��:x����3��iK�<���uF�{�{��cu�!�D,J_K_�1��?�^�y!1�A�P�ScL��ߗ0y9��a�b���Vс�CޏN���B�I���.G����_�����`<����5c�;J_�������4��W��r�-n�g�&���UZ��@�Czf�_,�"��Ƃ���W�#�݇x�$YR�:/���)+~t�'k}a-S�/�lm ���=b�9^<��t�m���mO8��,�/��Y��:��<[T{�.����I�F�)0xA�!�^3�<��R#(���Ǽ�+���ڲ�s'���O��qs�`�ѯ���N�*��I�U�E��8Z�L���1Zwކ�Pͧ�Dv��*�g�g-a/��P/5S���c�l��]:~[��5e���יw��(?Z�s�v�?��l�+��CMQ��j��*^(�x]*Y#wN�?3�;�v��q!�&����8DSM{�;���"�$�&�p�����2i|5�2��YD�#���Ȭ�鷆Ғ��<��y�U���AF������ot��U��4$m;;(�$v+H2��8½mn�G���`N{Coe�S�~J�#>(����K�2n��0 �p����ٓL�S�i�mBv7�S���l����ԁ���*�8�g�ҎÍU�k�]b[��j�yy��>����m�6^��Ə*�ñ��G��"�X���ա��[U�"�t`�F+T�s0M���w	MJ8t5�kK�З bהyM$ʸ@`���%h#����u���,I�T��N)���M5���
A�7������zL�OcG[�
:4��kh ������V��)53��*ѥ2J,�s��*3,���9ܺqF�b=�즫X�^l��ܝ����y��q���sY��G#8Ê��(?�˄�::�Q��r��G�HfK&�iO�dM�Q=�Y�������J�	Vͤ���Z�&R����7a��*��-f�':��@�'�Cm�A��aM�!��<Ek��>�&6:�,�n��2&�Ǡa�n�p��d�^y(cu�g��8lg!�"���?�.��O|[����� ��3�t	�G�3���a[.�&����m����X��7ǖ�Ȇ� Gu���������.�rmq�x��!f��'P���"����@3��Q��d�����G��5��k�UC��g��x�T^�v�DId�|nl�jAN�}���z��v��at���cvT�!�oF�)Xu�鿝�Pl�tl�=�^�����ռz:~�)1�)�x�/r4b죃Y���;�gI]-����J�u��ԙ@���X���4��f5�A�W;`� ���M_��g��=��Zsڀ;kl�]h��p�X]�Oy���rH�mS�I�Õ���A�;/�d�p��B=�!��8����sjj2�ǿ�k�J�%r�����٬�;�Zx�Ͷġدld��%�*�Z��bf<��}���+2�X��BR�U�z7(��t�߱Un�����Hl�������i���oK�=�Π��`�H~�(���^��2蘃�yr!U~� %Ŭݯ�sC)
�)��%�9����?�N"�{� PUF
`֕��Q�!U�_��6՝,+�l�r����ㄡ�E*����]Y�E�aN�}AOzt�\��8
Y��}R��f�S@�N�P��x����U����T���8G��m(/�����$�ۡ��*7��9�ccI�1ڪ���Yj��3����,�]i�������l��� m��#�M���@XӅ�q��B�0�-ViBp�3L5 j�^z�܁`�)!�{
/x�!ꋹ��^��:�w����I<�� �r�UL>N	� =P�؏��rڢ���0�"�(��/6�1�c_hH����)���o�2턦��������+�dg��}JF�L\��~�'T[åTI�R��l�3�v�@έ ��ͰdQ�)O�߃��/E5|\��&�:�zLF2z��i@�@X\���&��ADP�,:���4�H�2z-���
������x/�<���������!��W���<�@�-���D�@{c��Z��]�$OvR_����ݨ��W�Rs.�+Nx,b����X����\/V5�����ܖ�(e5޽Dg�lN��8���u|�;�~b��������ԫ=(uPe������>\<M��2V��k@��$���yd�1�?�Hl�$�x�K!�p�E}���n7�b�T'2#**�9E7����=?����$6&o-tn�M�GÄ\筌;�c}�Sbe�l�.>��O-t����X�VujH21��b��~ۼH�(c�"|=ΐ��V�a �H��a*pv2��d`�ʤ)�9���k<���sH����BB`��!�J
?yx]d�NA}����1E��P��/R��uo���̭L�Z��+�X��!��.���cN}�������"D�BC�&[��Sx�- ��/)���wڍK͓���E��"�F�a���~�SA�u0#����G��鶇J��]V�"$�����xp���uK&���� �}l�.��n^���̩���+	�J��h[/4'
/�G<����ϒ��*�(�Ye���s9M
Rf�󎽢�{�(��XGFQ�;�V��	�.b�A��H� ����*��RK�2�7�I�f�gv��'o�y��6�hNW�"��ٝ��*�8�Z<�张<�L�jj�J-ζ��я���m�D��2㤖�X,�T��y�K{�5x�^�3@��X�9�}J�Ek���ֲz���:�	���Ւ�oX�����s:Y3���'����4V!�����A������Қ�P��%�� 'F�W��N�*��9Ⱦ����Le��Cw=/�/�s�ն*���dB욡����SŖ��۽y�1�����[���:� �5܁�UJ�V�)�77���м����]�.��'�E��S,� �QJbN�ڣ�#?���BQ����#u֞�frC�f�O�F#���N����ʩ?�lV1<eVa,�m���~_�����$3�H�\��2 ?���Ph��^���MBM�m�i���$ER�R�:�/+������4"�/'ӣ~��v�Uާ��yk�f���a<��p���Z����L�[z�\|2�J�cl"Z�E��}��:��L[C@V2U�V�ZH'8��$ȋ�>��D2� ˔��_F�a�y��-dC�%(�њ�;}S*��;��28�����jЖ����H�~�gPO�"�zb�(JF��p�-��~zQ�c�	>�����M�H�F:��jo$�r���~����d2?�-m�c����r��hJ���82�;F��D�Z0�F�(���q�5�-9�����d/6lƵ�\jk��|�)�T�>���QΝ���L,s4����I|���)�Y�v�,x��u1�Q͒�J���P��
��)/=%�~�ڸe�xi	�b"�9P��[�ҏw��̒�7�zI%���YƁ��[-��"Jd��©����UwK0VZ�;Mei��.���%���a͎�zvʟ���H�]G��x�U�>F&��Rf��Oy�;
ـ�q-��h�,`F'FZy�\�ZWr�^=���n�2h��0�GԀ�����w�k�p�<q\�O����c�w�Z����1N���ՐT㦻�V�}p&�|֒Z*c��Eݕiÿ��w�s�f/?/���c�
�GP��tS⯐V����I�3� {���_�1�s0q�"x�����Ьu�Өr	�0^v-�=tm]Ԣ��k�N�� F�}:hVom�t���g8ua��0Ӡ���f���3��:����-�����a�4ϨI�՚�QBL�(���(
ܝ��݆F^8�	�Ur�l��4��S�;�_K09���{��
Ԍ%�w�������Q@�)@QyǍf��Ǘ��[1x���U�����נ�#���kW�HA�#F|@��<��}�F�e�e��͝(�>�J(c�(n%6���������j�i���5�;��6�>f>lo;�f��yNh��Sj�V�6�x� )�
�bo����<�4M�;e���o�
�\H�Mj��碰�
`Qw�fF~��S���K#ٮ�_1�Q�pK�=׳n�n4{#/�Ӎ<Y�I0�n���v%K�=��ׯ�
{�^%J����2��E�Sf��#��$I0�L��Sp����Qa�y�~kti�IN�<����e$�<)�#����vZ�?$d�~���W%@n�Ľn1��~�s XS[��(��b�j=l3>��(\�uL�lWJ$�4wD�n=�"���l�sbE���y�)˻��L,������)��a�,$��͊Ѯ)F��^�a���Z��Vk�vk[��(��W��< �Z��; 6���/���E��N3�u.
{Ȟ9��p�y���I�i)9�/�a�a~k��`�)���1�Hjc���$�2vFY�r[),z�YF3$�hŕD*��ĥ�o�7d�ι��ژ���҈E@�vV�e��d�x��=" ��Ѿ-�+�q?A{�G�r]��q�9�1�\��s���9�K�7m&ޛٽ
iќ���	MO*<��w_�ŢN�#ƚ��I��k�ΰ!nN�H���5����#��!���{ϻɻ�.�r�����\�`�z�zA�J�NXn�����z�/��ׯ��T_�֗��~�ɫd)`�����r�*F�HP���D�h��bO�xt�#kF��0�i�eh�i_Z�404��f.}|Mb�í�}�=�"M�����X�eB�����YX 3�/���W���GϺ��Cpo+h�v�an����a�,�"�9PIφ���N���ݢ{� A�J�ړ����<�t�� s�\��cso�k|{�)8L�gN*Vb|z��Wy��7%�=oϘ��m��/h�Mӹ<=��<�8t�˯����b.�xp��#�T�(�ʨKG����o�j�\_i^�0I��:;j���ie�o ���������G�Z円Z+��"����w�r�� ��.�Vb#�6��Θ��é2�P����)����AAo��V5�����c'�� H>�H�q�h��N��ƚu���KŖz~	Dg�Ү�ª}��=��tCY!�g�@��T�c�4��H�O�)�������u	��Z�6�=x�{�s��w��D��G|�{�I�lB\�Ρ<)��b&�֕I��c���z��T��:���Ҵ&}{
X��]�K;|;P<O�85��|̼�����̀�!��%F=�r7���ߗ��K�5��84GK��M�Un^�u�1��㨠�&O�?y������a���|(���DqT:e#�y���6�1�%�`T˴��{B6<���MQ�|��zq�������t�;D<r!8��?�}d���LJS&ѫH�>l����⭝�=,Y{j�Qȟ�]�).�W.�����ބ���\V]�%hC�Z�n��&��}�����\�}.Z�C�H$j��X3�M1ѴC����$N4w����������nKW��:kC
:�~�H�� �x���0@�ZH/.�f�ܳdxm���!��[�:kբ�K�-����*$�ҼA��nkL�׷+x��T�vQ��U�N�������0�Ei��K*Q"�:^�ϊՐe�(ְ�97j�T���������E	4�Wm%=vHoB;m&qABO��h9-�%��._5�7I0;��vn��^��J�ٛ����T�ŉ�!ڲj�E��Y���C���[FR��~>>g1kT?�������2��R���?.�K@sm���֫��&٠z�C_���«e�t,J����<[����N"zG�����J�E�M�zx�� ��o�N1K��}V��4�
�V>�J��;�?����z�f�ض��W#���p�E%�e�4)�0�:D�3��l{�{*�}	w��c[*����z7�>W=�l�M�r��W�"����}�L 5�9,%2b> � jd�����x��a�-��	��h�&���Lݻ�"�_!5��U�A�O25�d�j�b�(<B�$�ØG����ǫ�m���
9�y�h)5<;�a�Hr�֬�3%�yF�$	a����Ü���a���z��v�)�$#Kc\T؏����h_[��&bW�ĵ`N ,��,Řf�O������w��rQ�؃��aQw~�o�_�`P�a|�M?�x�YF�(PB�2��Q��1)�2��3����kM�(�_UIerN�c��+(N�8t�����,���xזdJOńԌ��}:�
��G6M��6J®E��4+����Bv��}��ʄy^r�N���+wZ�!da���&E6��5��y���V���W2�?���G-c|��G!�pPg�A�-�C���H��)v�ѯ�����dzW�&�]��4M��y�¾��7$�d�Ь��#�zQ�����})��=k*2g:�!�
�h50{L�	�w0�K�nKN���$�Ҷ��N`ԁ��=%:_��bh߳�R=�4.��Έ5<s ��~��7;:�6˿ �=ؘ1��K�Pb�팸���.6/ �&R�$	/,8f�E�cT�|~�sO���ط�:v����0��5& �:Wz�P�Ӣ�|��Jd'�z�'�JV$�<�#(�E�_�0F��9���F/%]�?5W=dO��v��==��`�מͫ���$�xTw �+-������K����qs&�� �G=0�BH�*�z��������!d�v�i����l���<�2�Ƨ�q�w���&k��.1� �Ì�^�)snXJ���)��\%��n���w��8tEІ�(�cz�aA�EJ�D��ۮ%wVt>^���m%��͞]��*�@�9�d��T#�[*b�w��.󁂰�;��	���(�й�� c@(F������2��	0[^\�p48��q�e��Ú�7_}����G�v��2}��"�����8��Ef6[�������0�vk�^�[��.Ǆ��c�t7b���Ӑ���V��rt���a	I��\�/C�]�Bԁ �սX`+��X�ܼ8���eѪ��G�?k�}�{ɑ���4I?� �ne�-�us�hK:t�3��	�]��*��;���V���N6d[�1���8�L��􎦠3۸�d��b/w���j��w]��Y�δm�{ƃ�@zT4.���'�M����䃗�v�����\S��S�]o�HP��'� ��Z�݂�!�9q|*��y;9��,>y������jG� g
�߽}d���4O|�޲s&��L�X%K��+��bT�_T=b#ؤ��:��:�bK%��G
A�g!�Q�?Oh9-�$��wh�ey��ف���r�gi�{I��X��B��&���10����Mu 8x���Y�/��`��8�Vl��pЂ��j�wH��BT\������TYs�e���q��׏��ہ�ۖE��ۻ1k�$�
�r4֛[��^%��JB�쀻�J1Wf�	_ݻ��n��<r<�^O�FG���*��dv�s��y���3�X柦1B[�5��	������+A8�9���ZRo���"$b�Qx)�{���g��n�/1���溗�PaYsB�	�����}��\sVmQ�?C�g�J��A��\l���k/�N[���I ��+|d�����{�������!Y9Vt�u��j�q��[��k��G�$��;�>:S����V1��Q�/bC��W�n�\*s-p�[Hiv'��2�����;�������֫�Y�_w�>���L���w�Ũ�u�>!%Љ��A'�0	�8�'oAEDzgY�'B@��&�^|������]ɘZ	6�1Ϳ��>_U��ٕ&wEe ��Z��ЕzN���a�ÿ�9�� �~��H)ֽuk�_�h�'��9��D��%^��P��<�WI$ǂ��BUe23�M�8ɶX�{+6�;H��D�G露�Oq�5y�d�g�w �7QŰ�[�A���p:Xg3�A��c�ܰ�^Sn�V�P&�߼oO��Ѻ�Bκ��|�/w2'�C.�]�#��TB����Lw�}�&.c'��>����W�Dy�|*Cb��u������a @͛2�{`�5 Իjc�؁�/ʇ�Pbb�p�6�Syhh�kq�+ktjǺ��.<����p�/�9j߃9댎d�"3���2�� 
 �g|�g�"fr�E��D�Y�)��h�,M��F�j]�#{�7�e_��z�Z�ښ8��26Ak+`�R7}�-�np�P��R�K"��)m
ȨThsX���廃,����3/vl���4�dGƃ@z)	z ��nYV�K��PB;`� [`�;���`g)���o�?l�%��0����_4�?n'���S����Cl��M��L���	E������з�f�����|2�2�POwN�����9[�P@uUY	Q���_iו�^�׎8���u	Rv�	@�z�G8�+\�3-��Rr�.��+��Z��]<�݄��M,�(�<�%��/sq�m��P���C��>�#2??1��H^#�1�����`��6z�/>��&�y�B�j�h� �5civ�Y�'�0Xkޮ�t���o�#�=��
��x�0Y&1�k�(��Ir�t5 �u��u��4b�XLv����y)s�[̄�'$Ȍ�DD[�7�C3�D_fߦ?��6N�� ,��<j;-4�VJ���2�&eF��EBL$���4���X8�Q��UQ&��� Aa�?_z�4i��ݑ�ωR�-��d!|�B!S��Z�Ҕ�8C�-&��Ś�����EpܖL���^Se0 �#�w�c��?ܙ����^�	"5�K�� �a���E� ]7w"H�y��-Gڨ�E:���Ӄ��q+�Lhp��{>�F��*�)J�:Z�mjD�Z��Zw[���=���Y��E��UȗX����+�	�U��_����be[��|�v��`(�nfK�IOc7���E|��Q�m+P�H�?�P7�
я~��~N�4'��N�y��ep�+@`�&x�#W�|^�#�Fa�AV�4aҟ�Z�(����!�;äl�ѿ�I�a(&�iۜ\�OX���J?����5�vOS��l�&7�m���AИ:�+Z���vGXb��	!���̀�'��9��z7�te>�G�a�C�����RQ��#}j���#Kb86Bu�}ה��(:�l��q�W����"��U�N���2�=�G�*K@�11�7؞{q�_#:<�;u���/R��UÔ��Ѐ�QE��v3�Ża.�6����ek�6oЙs�4�#Ӡ.���!��M��*=��9�O<���7�����q��S9x��F]�π1�AC꧵���<�%�n7)�Ϟ���@�lb����z=��x@�lO>���|�������&	�\���-�2?R
>���Vo�O6�wx�SY�mo�S�&�o)�`ζ)Z厧(I~�y*�F�zkhnsGA�sՔ*L�~Z�(�e�x�������Ԏ�1jն"�,l����ű���!�Z����m.��Y*��m���|�
����4u��0A�%�1�u�r!�����&���>�ɤ:��'`���E48òjy}l­d��l��t%��2���&���˩!��=pk���.�\�_���KA�P���^�6L��
B����W��*��p�O[pfo�%|�	�^!Ph�.����*Q�Q��ݤ	��R�/J�\4����:7��_�!��������e��QO�܌ˑ�,N��!�~�	f�c��O9u$�i�+�n�H�c��IN\ �=��!	��a4A0O�{N��U<+���,�Zk��p2����u7c�f�Ҏ��T?"����O{��ܟ��ȣ|��:L3���J�(�%�������CBXm�M�7����W��`N���)�������@��YJNf:;���M4E�1C�� z꘽��G:�(eR	G�s�,� ��)BMwo��Z�	�j��f�d�K�\���T��8-����X��d Bi�k%$%^�$��W�@@���N�g��]��z��@���4h K��ގh{/?�Ո��N��al�鏣i�]�����:�+�z���8�M����{��^KF���Y��8%�F"sQOF�������罦�ˉ�$�)�ɳu����-��q��L��m�e�
9/��t7>�Hm�5u���{�<s�6�Hp\�3�n�n��ǰc�����;�'J^�d4�*K�V�@���0�-7�J!�Z+q�rH]�d�om����/�Ҟ\-�=��$$s��m��hz���z*���g߸��n_�M��G]��t��#�/�\=>�J�ňq�f�m"������k�K$���E�-h��&P�C'f�Ǌ�`�U�G��҄�f�Мfpk<��4E�3��>�gq��rbxJ�o��t�⻇���u*V�9�?�9�O���E3�l�P�*��#��vf�
9ap��&�����������9H�&J`-�o�,�ބ�b������;���V�"?)4r}k�Ϩ׸���"�X�3'�����N�c�Q����;���~��p�\(��ī�"o�P:��a�ѻ�Ê�mPE��aJ�(>�0���oK�z#.+���$
���ý4H:�e&�{��ӐO	p�x�FeC_[�A�7�DH���09Zk���r{�h�rҏd�nL<�>�\s�hz�}��!�R���!P���C���b�q�a_]��. �����_;�n��X�Z���ʠ�׵�����-	D3o{Ӧ��O��J��mz�![g9Ϡ���CW�E���	�$P��u�%��|} Z�4��u����H8�����f�Z�m�����0}�`�������.P�6��@S����@�o�O�$�ݍ/W��v��x�(vE`&�&�m>FO����7.�=��=�^����'kSs��{K����P %���_�ai|z�(���[��6�B����Z�T�����N�ޅ��pZ���6E20Pq9�4pP��\Y��G�C��;ſD'6#F,����{�B�ҢWR7�}���=��f�O
�N���)�5S�'m�Nù����.d�y/p'�<���� _�Ѩ@g�~�;��|hSa۪jkj�����onNy9���u�Ʌw�*���r}y��o�L*�Pxl��<2{ֲק�rY�|��i�\���*�o[�FbܥܪnM��ܿ����ZO�1��Z���Hjc�<�Me����`(�/���ob~�N r�s�.->@��e�i�2�M����o�N�M�T�ŀש�te裉@�C�6����5���9J7�%)h.��'m�P��2kZ廒��F6�����0o���*u�-���`���6��^�x�L�P�ce���X�w���S�����5N���N��������`���ŀg#J[)P�A��f� =np4Ғv}���,|�6���`�y�ۧ�>��6z�.)��a#�� Vم��^2����Tc��u�J˭�f%�H#e��2�3�֍��I�Y	����R�4��t�~�v�y{S~@�d�"<�I�O��F�G:Vv-*���d�nU!�ګ�-�a/�T�.��
�m�E��09����f���u���<��̒]gX��1B��X�~�����3G$�c��Ln�ʅ%l; =�X���B�j�mڲ��9��]
iz�u�x=UFDhR��>I�z�:xK��J)�)Iٝ��2[�:C�-��'�+���c�xkBCB��IF�ܸQui�*�^3�e�U�9#r/�ű��O����IpT51��C�RN �����N���p2���fYh�����f�Z�o%�<u���3����A�+����XY��m�	�i�sp�a���"�$$Z��V�OUO���F����ΝiÏ;򪖿D�o����;���u����jd����I~��/��=���t�Ȑ���t�-i��!�	�6#U5�si���Щ�p��~�7D"�NRt�%���c��}�!m^��Gw(��WR�\���4�7Z����*�{�	g���,���cS��o �*&;�5m�y�[�7ܩ���w���vF5h#��.J'��m^��]���	2gK\��X�����.�4
�����􄇍�0<�A@�zL`���Hf��Ԍ�[�鹰��台ũΈc�k����,a
�H�u+;�:�pc_�]���������#M�����γ��LΪhFrr=��<G�|�@��Qw�0Hi�,����.�fy&Y����-�$��[U�s[!�#����G>����w�i3@���~�-��7���I�X.���OF9�܋S�[U~CS�6��P��3�AƤ� �ꇪ����L��!b��x~��y��b��)�!��1���?��v�mbk���ߜj�^^��˷Sb���ʡ %�,�J�x���M�y�k����4"U�\dvq��zw�uV-@-+��d&�fv%M��t��G��d�E���� q�����1Y�Q[~�62�q_j�.����L.
:5�_o�&aQۺ�	�8wa{��0a�}\)��G�.���F���E��G��w�c.��u�o,#`��X~�ql��W@#�(1?�>�عOZ��_p�RZ� T1� �?2�M�ô_?~�@�����-���Ӈs ?5�<�⊺H��`7���-Q��u�k)}���� ��n��f@/ꩋ+�f:_�~��,m�!��l}���!*-i˰�ג��/n��(u1Y���(���)�%�3�P���.�d4̌�B?�z�*|�{�D*���a�:輪f�}�~o��1�6O=��߁(3�3U9����F�G�9�f��g~M\���3'���\�c$7�w5��^��xѢ�x ��j�F�2[���W2cB��j���<.'�O�#d,���O!xp��9=:crVٷ�d>�;��V�{����+7����	�60Q���	S.�M�:����U#�Ӯi@89�	�KC��WD���!����;<���/5!�z*�pC����7Vv p�Ϣ2��z1&���#���E*욡������h��_���oo�(C�I"�f���=:Y�b6��WCޗ�}�%��8U�+ۿW�%�wH�E�t��{���̕]D���T�؄/��\x������ݑ��8oU�V��@����<e+^�j�\���%$Q���6�&:�2�X��\Ϳ�B�-�}���̎�!L���sY��'z&x���N��e�8�G`K@����]c�9��Q��~N��w�q�{\2T		v���]nZ}YO�~Jܷ�3�m����6.e� �;��t}Y��G1!��퍍���
�P�����k��7�)��v<�P��!=��M��-H.��E�>Ȱ�j�j�F�4B�.�P�m���Q�ތN �͉��b���X'� -&����u:O�ש���*���9�PG�M����;���2a;|����ڪ)��{Ǖcsڕ�⤾S�O��Ġ�/hK ,�ޭ	HVT��R�_5K���◠RY���ɫ��d�s��_�R�/�2-L@�],�)N[T�
�v���{:%k�M��;�����vԐ	�֜q��ՌsFK0���E��9 wD��1�YɆ�i7��x����t&�q�aK�
4��<�5�|6kdw�X�H@QtDHsO��d������4��$pc�5�=���<���\R����6:���3�j(�x��7!�!Ǉ'�Tp��X�#����;���!��@}A�Fh�3YKibE�L�J`�u沓��Coݮ_�e�GwC�`��2q�H�e�ͥ�jU�51Xߧ"�&>;y
t�2=���y�g��1s��m�glJv����rU�(}��|N�4r����VH�ʱ��R5а�n���;o����J^�NSTn��:�������w�36U��}Ͼl.�T�y��_���41�����G��+������w#�J27)�F���Y_D�Bm�4Sq���+�ف��&4�����Y�!ύy-�X��J@��*��8�����&���)����|�MХ��g�O��q�.���X�@�%AFjyU7� 4���5s�N��u���Ddg��̺�,O꧸C��������]$.�#0[u�����n�
�+Y�L�	��h��g�$wY�\�07�P"��?}m�Eɣ.�v���ƴ�&f�:�@�������WU����2�Op�I����Qz�o�%��6����:[�z�w���%:/��5����G�O����;Z3�:Α�m_Bq��~]]��܆d��3��~�O�����`�@L�?��T�t�b�-G� �ha�;a�P�vlu�u�l"�ӶM���M�+#�\��)8F&U��g#R���ԑa��]�7���������e�������T3��{i�J�z�{�Tyn3�Q�2�W�����-!��OCS	�iw��i��-y2�ĥ_����|7�`[X5؞=���07�$��"��SK`���� a�iR�]L���AiR�'g��,��koY�=���O�v� �m{m�/�#W�T������mI.X ����V�ߣ8��O�w�2ocr�yJ��*��F""D(k�kR��K~+{t$����[*-T7�Y�����|��?k��NC9y��V@`��^B�,�M6z2�$V��㞴����k��kC,z�4����xZc���/~CfA2:U���LR��4��_��0SJ �rR	g��gH�����O_W��a7�]��L���`�&��JB��H�ݕ\��Qw�0k��o�U?�p$*i�ԏ��Tѷ�C�㪗9�7�5Ѧ�bx>�X+>1R;�E��B}����]JA��RkU��nU��5�#�2.����9��4'�nWZ������ �g�p���
$ʭ'M�{�,��W�z�D�?۸g舸!��ÇE�&+5?f�������b'^#�Y�+w@4�����b�i��m	鼚$h.9Y(bD�:M� �Τ7���{t�|J��d[�v	���ŕ58qh�'ؒ\1�)�n��=�uO�4L-謍��E4b(���ᥩ�T�z�#+�@J��XV%�Q/�r���/XO~�)"�,S�1��X�e�,��kj�I�V�'�H��Ɂ��D�Ωq)�dv�5���*�&����,��!} ���"C���������'�֕��yY ��m�n#r����^�J.i�(?��% �>Ń�d�NB��'���ꈱ¢�ym'8�9kpr��4������YME'l�j�i�`����G�.����z��Β�Yt�B���fN|Y^\��Z�]��j4��$�Y�|���+�ƍ��֓���v����T�!hڔ��&Q�ˈJ�~0G���n31��h�9��eݺ&# �DK������r��Pؘ�i���m��������:Ӈ�tF*��]`�[KT-�(�'��QX�!�n�=��`r�K\B��������n�_��bd�l6e�Ld�V���|�~z��n�H��o�'�[Jר`�Fϼ��EO+���	K��a^�E��c��Ͷ��\��~��_w4_�FmU$q��jW�/+Qc����Ko�SP����,M�d}�
9 )�|��n1!��e��V�ۧ�¢Р��ŰI�*������m*�Xz�!��0."�*�d�����E�Y�]7���mQ�`Ǵ5R�#`(��`P�h'b��X��A��W���t���O|[H!����HP�G�t��_0y5ׅ{y
�����H������?H m��W(��F�f����Y�a2�2��|Ӏ�2<��������6�tQ�y�8��~UbB)q�q�1*�f� �!����h��V�ĸ�ba2�U]�\F�]�0|��@��l�1�"�������j)�z�;x�*{CI[X3s(~S��� @T�C}��� F;�E�o�4��+MVLe![/�m�\�6���~Rg32��!�@���?/jG�s�u�n�ԟ�L����A�؋��5-V���Џ4���}b?���������	�8ʩw��2����w�[Eb[���z�χ�7�����e$�7+��izv��(��Q�4j=AR%�i�e��h�Vτ�=N��z� 6wPv��+1�WP�#���oչ����>������;�l�@a)����1����!?/�*&� �̴����~���m����dQ�z�(��u�4���H��9�2gh],���-&�̡j*�&��N�H+3s庁�=�X�P΢>�^P��@u�*����/X�#$���C�έ��MƋ�Ĵ	y���X���>���㦛֙DHaE�d���X??�]?vا�g+gs���=�~S��0��K����5j j��4
n���!,�ڠD�qP���bX9�)^��㔯A�5�w���}�]� #?X3VۏaF�iL���U���q���� +wqI��˨���r_�a�5=Ge֕J9��ܴ�c˄ �-�F�7j~�~v'��e�q`�Ф�)o�hl�k��;�Ϫ�z�1r�vȃ��%f�m�9� U6|ŀ��E$��h�2$71��%��ѡK�tO�C���01�}�G�P�gwJ�֔ ua��1�|UL��N�����0"#6o8}`o�T���)��SA2_�aJR��3���{�[�a�N�U���s�0öO����������4]���g?w���5������ @�� ��3�G�/�}	�J��h]5�/Fc�:������Gn�#���	���̖��w'��1���Z[�N'?fz�Wl��[�ve��8(�E��2�K���;�:���9��R�=�1a����Za&堛X/�tndu���:C�೫r���Vg��,JrjS�x�8�i~"}�������>��I{}����hь��^}��L(p����6�7�7���c�[�rz	N�,쫸�ŎJk`SX���>ڸ*�H����V�֬�J�ϊ] g�s��_V?��������M�h
b����딸�(�2��V'�w��ES�9>��X�D�I��3�?l\Pb#L��������6��[��8�a��P��IV�ni���IW����<��%����֎�����0He	5s����t|���a���ɰg�x��2�Ll�v�h�啼2l��͕9V
kA7��P7�`㵝��}]������p'c��B*���������8�'�f�rU\�&G"����[��Xȸ��^^y�|�ex���.�k�F_���-a0g5�#�B�25�e;瞉�|���a�3.�J/���t����.��+��;k��%�`}�^�l���̮�,��^5,�A�J\��2�=��dG�n���ݰ� �j�&R������-GաxIc���Э7{�<��I�y�6�Bf:%_�\|�c����7�N��>�t��ҧhV
�u��_y��K��*�ѝQy;f�0�ɉ�Y���j��*=no�p�g�W�.��e�(I͛Q��%T�7 ��ԃ�=%�j����KE��E//��y?)U͚*g3�!�EC^��,�ݢ �X�c��9;>�L�-(mt��"u+��wq������U
��d�+�L�Um��F��z?��$�hM�7dJ�\[rA4cױ�e�+6���D$.��Y��5T����!�|F��wN������1��-�\SNj[N4��M�*��{��e��)�潰�0��K�_+v�� t�OH�yd��^��'� ����U�A�3'v]���nx�@֩�n[bn�������>R휣Q&�!��,��s�?f�1����=��E�}Y�C]���p-�]�)7���x}�<�w� s"H�{���WI��Q�����$4]>�Z�l[=�n/���S�{D���]��S�?���;`�=�Ⱥ�^\'��^m=�M�Noڦ�6�4���D�n�����g�S�B;����tr|"0lg���?���`>pc�ӟ��t�GZp/InD�X6QS'��m�`��K����+�Y�o���E,y��I3�?��Cg\4e)�d�G-!���m�����W��fӻ=�?�T�9�>|ZSt�8�E��z��"��GjZ��}�,�/R�y]��лc�v�L��G	�T�Jl>�%@V��Q�[u�?#Z�1���
7�@�[V��6� ��OA�����W������J_�	�C�����B�rǇ;$ ިw��?���r��r=�#�D�������kt6��эJq�����o�C�5In����F�kPd�?�fI>,=��*~�ސ��������Xkh-��x���>����(��-��8����f�4��s���z��e�;&+F-R��5�%)�p:��wY����f�1f,��u�;y�n#�t��u�x[_W�Ͷ[s�Jsu'�s'���5LZz�s���8�F��30
�
f$�̺;/�c+���*e.jhn�3��W�^����ol�<?=+�'��o�=5�"��=8�m~r�pJ0f[�%>�yj(�_�Y~j���J�')�
T�Bʊ]�.�cl�N�������l�`�����61w�s���SA�i�Ȫ��MZ!]�D�ḒEu�C��\�@��L�A�����:�:.ى7��c����
gַ�q��Y�O�5�`seh|�|��o�4�4�f��(��~���;��� %�#
�����0��;Y�B�6ۈ5��[S��V����9�2X�ܽ�=�n�wN��uK�dc�ڒ�l��a,2��q�����ea0j+B ���Ti�%��c�A�W�[�}���}�?���u�ͩ.���{��|6�V�d1bke��@i���<(�43@܄����P�%����o���v���w�#�;)�X/��ҮB<���.�!Ż���jEL:�Y	� #8}8I�yP/�,XJ����Cx�c����`��� ��<D�ojd⡵����粇q�1�Ĩ�/�p�ۓ���n�b���x<)ir�%��3��y�b5g*��4�G�o���JD@|,S�~��ѣ�U�pO�Xq�Vxo?������SC0��.,�<� c�X���*�Y
J� ��{����!���z�_UΔ3���ԱVgP@CE�"�i����������C��*:[�J�%6D��J���?���"J����f�
�@�ŅY$(��$_�>��T�ϥ���|��� W������pv.�U���+������A��8N�tf�lfIp�����I7F��;Wj/�kT�J௎G?1�y���s��G�{�)��L��Q^��� oX�N�1(O#Ja�&3��
��㄂;Nao���1Aj����w�Ҫ%4�C��i��������8 sƆ��D���{�8X)���˒���.��y��-���w�����%����+{s@�a����[��d�A>[���6zaz���^������ .a���M�5nj�vJ#�+6�\?`ϒY�~�qu^�-��Ȏt`9��AwM<������C�����f�d݃�M�T�h�Y��;���O��qwY��]X?^N7y�Y����|��T}7�������`�<��	Fhk�m"x�rh{l�9�e&��fZ˯e�M|�e���9�l�		��Z��OS��g��eOzG?�'���ڡg��`ϸӱ�kXj���7�jCE^bٵ� |�"協�-�#�k~#��g�������UW�����B��#�Bɻ��C���S��o@KL�IC��&LN ���=p�+Cs����j�S�|B�
�a��v����ml��n4�Ra��欮�:54F2�T"m񯏽��1���#�#��q~�Ο ���6�;k��5��O�6ýw������'<y�D2���K}��c�U��K^�Ō�DZS������N��.��5fQ��0����sV� �o5��Ї�}Z������[`�`�?�Z��M2w��df?���F!r����s�_O��/Q�D5��5�#��4��f�ز��}1���O���Җ�^^�y�4�� Nz�@�K�� m�F���z{�����+��_g�Y��_���䨑�����ɰoI��"��bDjΎ 
�P'�bZe}���:��D����=���1�QS¢�yw�@I*�b%[��W,��1�}�%�M�΋�]ϭ�I��z��i}{�m�Tm 5K撴���v��ֆ-!Զ;��:�$K��
xE��*a;
� D�1q,mO!t�G�%����R�%�$�v�kXK	5_���u�J����YZ���"-�f'ƭ����m5���q��Jo��yD��r�Y�<��"FzS�҃x�zey4��G�>Iz���Z?Dp���Z�C��ڡ�����s���[@�k�î��9������[���Z_{����-����|�U�?%�+tQ=_6�c�X$����:ٶyM�����!�Qp�m���+V$̳Q ۮ��C�B�r���|��5ˢ�݉��ɿJ�F۔Q�s{)B ]���&�k`F��"�X� �Fl��K�3D���U��2�QM׷��'�����=��W0(��О^$<��珓 ��`=
=L�g�o^$P"�W
�Vų�Nn"��֫��8|H{�n�(,oRP+�� ^�b�W�؃}�D��O� 5o���z^i����8��/kR���y��;܋I	aMn��'��ac�l���L����wIX��k�a�]�t��6�}o����{����C��E����QyH0�::���]�/���~n�Xg���D�_������Si��ȑ�^� D�ʘ��7���L���[��
$x�Ȍ��7�	�:f
b`��,�̉���4�(�%��ɺ�ǕhCC�Q��ۮ��#1LVw;�U��uo
^�I�R���),���0p���!�mG�IF!�0�Al�(���Θ1�iW9���;�3�9^�c��%��S�X����0t��A�ba)k�0R�ay|�L!�e��|f��b�������JK���M�>/�:��\~Ñ�qL�]�Y����}En������лz���UN�Tw��'zʻRz%ㄙ��H�l����9�j�N�iݽfTۇ����O���^ꤙ����Q<�!�6�Ϻqƀ.b��F;����+���c�,�r��e�ɸ�~��C�C�_�3*���R�l��&0P�K#g�M��Tڶ�q4d������b{lw[�&���{3��ʤ���-o��0�<�X��l� ��'��"��9Tm8P���nl�ZI̹�K��
��H�TǏ_+MlDSs�znZ�7�ж�����m&
����*PaK�`1ܢ�{����[j
u��˅�s����z��t��V���f��cx,�$� ;��O\rv��^%��R[��p@���b$��m�����)�3���>��C1�\�b�<�<���+V����{~��Q[H�T��0����u�'���,�&��J�öޢl/]�\V'¢��8�삺'x�iBХ�� �¨FVx��(���Ij�,�"�%�E��ZX��5$7��L_4c��0�8��7�bV�[�Q���I���R�[p�!�
:~���iN�3�Y9�7�R>�K(�����8@n�Ph��"�%	
�s� b�+��ʆ`2G��%}Nz�Cs?��N�O�ȃ�}��E2O*P�'�Gzh�� 0�������OS��Q�	�5��NtWh�"Y��W<�J�7�
=2�~ln�bnK��*���[��T?&��^q��4��)�qF���T�횜%DC�x=��m�'��U~th�o�;Tq�����[Su4kNل�VX���A`����q6ؚ�T�6	���ֵ�z��Njay�
�v]Y�ւ�y�FA�I��P��ɶ������.D��9_y�@�hx�D�5�J&�A�	b����У�{���{.�O<����#�_�W���!K�+T"_����F.jd4�Ƴ6��߾S��,��u�h&բ֩��vG.�s+�\J92E�nLy��
�G��p,pp|a������4���Ԧ������9�N*��|���PFK�D0��h&H�<��9h��>!�R'��r��9�3,�:F���i:c�a1��4ż{tw�����k��r�t�g`��k�E��	/w��B~�:mOR%��
�(�ڔnH�+`�4tg���0�����kR�A�Q�r��"��cG���eu(���:�����x�.4���I��Oz�Ѝ@_Z�e߸f��1a��8����f:Q��zasj��EAa�".��"��>���CVq�u������|Cs�q�W��#����I��G&�!U�����fg�sǻ�_LBz�=@�������oȩ�i�Ü� K����V1���˫�I;�@h���C�&.rW#)�s˻���J����Td�L��'`������j��E��ā9�ս�:���j���P�p�4c_zw�+n~O��+�H�� ����7�;,��${q���*�N77�^
�T���@���������^h|�� ��s�>(�ٮw��|����䜟l|�3�K';p[֑�Aw�>¡VIX=��+�e�'��N��!�c�|.2�i32��%g��+CZ�����)T{5c�-�FN��Ľ�`���It0�D�X�F�p��HTR�MsyGH\�D,�9R$*���,(p������l�4؃3�v�¨B��Y�vw��D���Y��!���Gz�Q.�����[�X��XkA?f�&;S��}��{E/�C����U2��1o���n��+鎋᷁g+��+ս�U���E/멃��xqؿU��W�����b�%�xK���\��(����+0��;�o�U	���<d]��}Ĺ��kx�`ci��A݋8�r{�l��)	L�/>B����w����-��&���$���׼���ٯq�&f�
W]agqG'"��+@����G�o$�`(�a�n��������@{���F��)PAG�8i�YB&�s~�z��q*A������W+P���ʯ���2���Qn7Q�
���IH���373n���!�8��Q�v�u N@���;�Ԍ�	2Gp�n���T��~��Cr��j{^**��i�.79�r��cz�Ƚt��g�OT��k�#��D�M$B���ew�m�~c�`'�8�u?�t$�O�_]��*{�;}	i���Gh/�z���O
cш7D�4�̵�T8��*��j�1&��я�����ل:����妢�Z+�ҽ���b��2E�S%%���f�$�5�Q?|5�4���V��W5�\�	@ع��%�,�3_��QM�H[q���g��QR���U����h�z�Fw�GQ�v��lT�d�n|�W�����[��$�|�T��?�0�[��a^(�:�]�M�/?L����ZV��N&JL~�_u�'��������O�	��x ���07Y��`/�g!���k L���t�)L��S��֪suG��ؑJU-=�\*V�"��d&g=�,��(���/�&a����]J�H�����X\XQ��Q�����K�LU��n�� ��Q�O�J��m���-������T~������t}���2���=4M�h�<�b��$�ǧ� �SGџ�7H^K3�=U�WõQD%�ӓ۔��-���l# ����ε]e�+��Ppr+%��mb�[�e,������l�)dތm�X��	�:�T����N:ii��<��J�*Y�H{���'H�d����ԭ��YP:�bKn�����K��õ57��� �-���}	��Y��^��>Y�c��">��'�#����2)�:����GFp,�.S���\���zA%�i�9���+�,~l˝���5���x��8���W�b�h��f�|srݜmmQ���T"ߋf=�]/��Vp�8E�*{a��^
b��4H�E 4���(�T泽`���M��S�����"��(R`s�=���l�֙����j���	��f.� �����+��R2�E����f��pg}J��Pd��d����9+q���C�ʟCA(E��;��j�\ʅ���/r��l��h4�/G�!D+�̉j�a{��u��~W�oh��������]8'm��Z���K@%mO���S�7�9��C���\��XA需��K,Dԃ��י�i^��c���٬U���_��g>���+VS�nj4~ǅ�Nժ9�6�?��q�J�FΟ�����<�*������{^�6Tq3:����$z���%(�y�xBg�Ι�|+d��ZL��	F����Y�C�u阄+ )���֯�w�>�������U�T������s�W�"��t".LP����#��w��B-T� .�[��>�+bUjz�?ֿ+�1�8i��m1/�+8����x\�)��(����t�ʤ{Xot�ʪ�� �r*~�@�QtO�U���T�E��&?�tH(�;"L �� ��^�KE��}6�/��������$}C��i�f��w^�fσw!%x�.�s!���$�h���%VƑn艩��+�Ԛ��q��T.C��
{�! 3Dڮx�xDuD�������i7n�7�FSU�W�ﵲ �u�N+�-�A��q��וoR}#��y������/�Ah^)��k�ŪE����B12}D�>�/��ə��k�rW�8�4{I$ɻ�?�1�Yd7�?�	�U!�~D�,��$��GPK*�r7��I^a��X\#�S��¹|�zSuu	�_�Ք�{�1G��ዥ���x��[&EӶZ�K���k�K&ם2�fO��nQ�I��003ri����8K��D1�^\NRMT� x&�QK:$�M���ʹý�J�YeGϒ��7�Ć\�g�<���pO�	Ԕ#�uzN�_��o�y;��,?W�rC�X�FE�(4��.�hm\n��%���U�+ݺ�cV?�r�卻u��BT����3y��c)�"������x�w0$�k��b[�N��� �Ы���)WN�����3 aμR0ە���L�	X	�MѶ�<�v�Ys��=x�8��J�b_���������^Q�����oO�Tf��t��"�0���Hu��������(\���q��PQ��c��}i�s�K�/������:�h��q�<�^�K���k�ZI,(ݩ�*�c$k�-�]���K}^��ݎ�ܠ�1�u������8�m%x) ��p�Y7;�	���2di�ΐ#�$&+�x#�~��μ����S>I�f�I��8X
��,�#ϲ�8�O;�oz�g�Ê%���(�n���_z��_�p�S���L�����}x�yvu���#4�`u�Ll;�ᮕ��$� 2��_5$�mG��[l�wN�[�� ]�JK�,I��~M��^<R�pt�C�����R{�6���T��'̮"$ Nu� �|�4J˟���R�ޠ26����d~So|���Q�s���'`�`6h@o�������*�Ț?Ɣg?�&Cj��h�/�w�U�'��&�Z=gɑ�� =�E���Su��n�r�q�X�6&M�	Z��Ѹ�^I����T.E��o���	��S�� !x�K�ǹq�Vo��������\Qh~��Uư����bL�o*Nj=�}�l��Ӳ�h�UB=$�׶(j��1����E2�Y�r�N�f)�c��j'�9�,�gc�Y�M<��DKP5�ƳĨ<�_B�����ɗ���ww�߼�
$��u��(�(d�Q@���g߇�S���n�m��{���+d���z�ko�{���\U�9d����g��qYL����n����5b��g�=��/��HԈGƂ��H'����O[��
y�)� ���b�������&�m�E�����V
�L鐅���K�s��Ӿ��㣫�z9\ਝ�?�A��2�lp�'F7R|�GP7���8�1��f�&��4'�p��8�ݨʾY��OZJ��D��ZG�cl���K�5_��O`$�$ɠ������N R�7��O���|�U7_LMi���s�CV0�v����֌Z�Uǻ����H#�h���7��L��4�V���W1���n��c��-��Ԩ����iׂJ�j8\[D�x�@�*��wm�v`g6���k�V7�dP��<�r�~�6����Z1�\c"S�I>��(�Ȃ'9����]���������`�y�,���ڳ<`�̈�^p�u�������.K�L�<�[)�v5�W=��ϭs�&�e��sk�w���&��w�=�_G^�v@����4��Q�G��-����/i�3x+�� ~�pK'��<�y��/trh�y�����k�P�/L�E�v���l1�z��+��Vj�B���D�yV��Vv����ƍ�&��R�����^���"�.��L�5��:k�0/m�\��Q�M��k��F��+�qX��9' �gY����a)5X�I�,��N�i����}5 �p���\F��~ o���p�(m��ʿ����S����PLT�"ƫ~~�ְ�y�+0��H݁���*������H+/�@��4~��+,/4;��8�=NEu'��yļ����H�"��	����H�n�a^_�H����BR��;�x:�g����JmCR� ����f�N0�3�8-��QU�);?C��[�q��Pg.�T�"�2x@��T��'��n�j��5�3���1`g��Ee�їt�'�C�g|�����ڏ��WJ4:��rّb���WZ�qV��qI]��t��[�=�T?7-9T�������_�М��D��r��o�]�(S)S�% 4�����=�������x�o��E<��¾�9�ILK�jvN��+Eɻ]:�Ĺ�VٵB����%"�*`� �O�TS:@G���GK,��+��}�-X�lv��_�F���>�9����-}[���3�c�a5\���a�zw0@��^aK���3�k������2B�`&|�h�ĉ}��(�.:�Y9A�WD�nD難����d�2���)��l����$������Gtm޸�7���e�s�$ij�	�Ĺr�^sCa'�t�����T�av
ﱹ�z_f���W����n�\�(��Iͧ��3(�=�g8�5�ƃr�H�a���oz��+c���� .J�� �	����l�fX���z��V�Y�V��h����n廘g���A�����ޕz��n��|v����]�<&���	�R�?E�ǌ�|%�	dm<!�ǰS��\��VQ8��
����.nrRic�,7_hl���9�8ë�?@y���w�\ܴ�^�@/�ǀ���=:�	h�%Q���X��7+JL>�R0�r�}CS�r�&la��@�UК�����W�|�������j�H�<��W����ɴ^�d���9v��
ݨi�mS��A3ai�Wܕwry'�\,e���-�-(�ph�2�|
w��zSp-�D��
Or�>�l�� �_k<\:���]�$&h�t�F]�ǹ�a�����AV�i�d�~�X%G�h�4�0�;
F���t[P$mz��:[��*�<���gZ:��zg
&4<��v�_��2v�ch�dn��U�J��:w�_�.���_�Y�=��E�U����l~(t�Loy�ֻXT�$jo��)�y�ifzP��	U6���j�T&��y��6�Xҝ4>��x��G����Y�$�*����=b�'�&�� �Ng=���ʤ+��Q�,�!���lZ�N*k�}qt�7̫)��!{v�Pō�9�W����$��3��l@ �)&~�1��Ih���Y>���:V�"���"oLw�3.�>��Nк�\��낄G]*5H7�;b�������w�9*_�I���I�VM f�mA���f��u��`uv�>����քc�H�bI=e8�r5G	�u��]ŏ#�K5�o����m`7Z�����T��1k�V���؉�,o�wH�,��<�Z�8���h���A�5P����]�P޹dA�B����S�T��+�.���Qhf���s1'��K��a�w���,ڨE�cm�fҡ��J/���q2��]�uɳ�{nk��\�Ԯ�	+��S��&��%�����x]�Q�y��)�;��<yb��lTj�FF�/�-��c����0��Q��/��1O�����6���L��D�'�6��qS���5�rU������A
��+��徭0�V��,)س�I4,'�DO��(�j�r��g�'�b&�(��t�o�V4��s��W	��_x�n� W�;Ng����*�{s�Z
n�|���*��)����d"➖��z��}�_��9ge����=�+�����r�{�G&a�� S�� �:R�R�	k�/Y�)7�&���]ݨ��n)�
8�"�b�y��L)@�c�	�����"�E�&�ݎ hf�L"��i��]
CC��^�b@�2�`q��r0��g�%*�Yg�?檱���`�:}��$��Ϫ�ӕX��*-�S?~�kl�׆K��>˶*
Ms�7�7�2$�<�h�ݴk�p��3>5����3�9��xY�bPtd�49��FO���o;B�l�� \t��vBi�];q��磢<D� "'C��T����ަ[7���=�4a�Y�}��o�x�a����R��<�mȝT(H+4��wi�y�U��t��#�^w�_y��]����>��v)?��_�Id9�M��{���5����R�x���w�$Q(�w���>���||E�hc��p ��('V���1��"-��Ԅ7ky��G�sl4�igz$1LU��I7���Fc�`��BeX��X�a�W�ڕ���U�;k!J ���;��J��-#�HB����D�;9������ܭo ��?k%�dY�9�e����%_Jlϟ�X�j�ofB���Of��}Qi����Y
����:�ym�:]��\$'J�o1��u����6��X|��*����V�]m�;f�	2�2�� �����s�����û��n��Y��P�4���J���䙒��Txp�xb����K$b�P�D����N�\[��<��>�{�[(f���H@��. ��
쨵�#������|i������r��z�c��*7��\�玓f�$Pz���h��B�b�}"��/tE����I�e�Ds�-���O����SE�	z�z�Q/�k��4���Z+�o���۹�L�U�U�YX���j���S��;d)�`O�u�an�j��S�i��$5�`B��]@�5�ˈ�7.F���ޟJ
=y�sy�J��$F���������&��Ԣ�Н����j��/�0���CR����.�K�͠�˦�R �	�NT yS`��k؝�@�}��$� RHBl���_�olj�(~�T�}�oׂ�C��*��N���Y��B�x�X�����Iv�ZW8G��vq�����刢��E��:�d_�.wW)ǞZ}��ػV����iFG�8
D�!��k	��<eMHi���^�Q��ǧ��Ծ�LS��m��Ѽq�Y������!���X�gk2�}:���C����X[�!�~�&^^�3z0�#l�At�ƈf���7������
��6�T�v�E���sRx����ۘ �2)&����D�E&7_�S�]E��w�h����.ơ��.��Uj����Ȓ�<���d?��[�X�^BM���]n�A'�s���w�Q��$S��{�c��,|$K@+xOS?ۧS�l��M}�R����C���Z��vnK��ש> ;7�#&䕬&zW�'
�9t*V@�j�%�I֔ ��b&X8O�xu|^Y�qVd�m/��=����r�L�]T2���`S_�B^V�����Wiv%^��c`ϕ�W���1Y�2K��${oN�gX:��Q�?�����H=��ub�l�Q+`r8��������V����꒮e,䪬y����H��W'�xӥ�,5ԟ�L�kKֿ>?X>7���&��]C��9��3� �F�ǻ�O��6�:�`bp#B�������#�8~o3a9� �%Aڸ�({�����=�?
�6D���+��3%���a�ZGtp��N��ta��Vqn�"����XLUu��J��h�rC�G�D��s�M�
��3���Z�u�1��Ț*�7���E�d�,Q�>T�����
r�@��%[]'�ՌN�\�{~�+�E��I`�Z����-�WÇc..�E��A��#)�Y_^Z��*�X���uӼq�=�8�9BN4�$bz"4:f��)]݅(��B�9W۫	--g�o��z>�ۅ�8�ͼy�{ D0�
�s�`�L�ܕ���Պ���cWC������z�w(۬��?�Լ�aJ���6��.I��Լ�?����[�Q�}��
�G��E1]kF#�d^X(MM����w��l2�� J�&'Һ������-�MFӆ>py��5%�U;/��'��5\z3���Ɔ��@ȝ�z��}��K�zyr�}�/�� �?L�UQe����|�ȱ�`n������=y�8{��yt٦�9�#PÇ�?�;������Ԕ<8O�+��S�R]�ğL3�[�%����")��5Y��Ձ�gc��6n!�5a�����~���8m�G����>�
�)]+6U5�u��z�x���a��2��h����s��;���<*��tJ�0�������RW4��T�"a*
b�`�׳^w�֬�{`�{#�s��Iw��_W
3vtU\{����XOe�<�I1n�Î�M0��_���d�!��[��\����8g�rm�B�[m�:=6�@	���7iS�d�M����v��MŎWN	�n7]U��pX8!����c:,�Q�E+�o�[�������W���t:LZq��y3E5��m��(<�o��냑
Ҁ8~+��!Mt	Ù|lT�?>�����1 |�A��l{ye^���Jy�:{�`%^�љ\ ��K̺�1�0�������k�����Π8��|&'�6��0����\5X�i��.�gv���ga������!�'����/�i�L�u�B$rXOQH��}�I�ۧc�]g7��o� ��&�1^��c-�6���C�+)
������f+#�b q�O��%��r�
�ktɅ����RQ����Y���E��,�}�%�@SR��u��\��ʑ֘]42m'�E���,y�\�b�e��Z�(����.{{MS�L�L��|�����"��>���C�~J�&�n��z����bť7��hv�Mau�_"$s���f��O������U�~��:V��s%&4�
1�|i��� �q8��:�N�Y���(iy�7��(��� �2�@7�
��2=�L,��~d�ȷ:ʜ�'�/�'��i|\�����4��Ұ�Ƙ�o��Tv��T�s/��|6s�`B�R�V�l���*��a$�WC4��%X���N��Q2	�>��N��vi()�_�ˈ�QG�[ʫ�'�Ҭ��R��J�߂l8!�oJ���f�m,r�FJ�,�Nd|�c�w�Sߓ`��2�]�)���;�m��rFt����l�37���=]1��P�8���H}+�ށ��;]1��)���|o��
V��lق�$�dn~�2G��t��L�~�g��|j��<n���Q�V�-g��>ƍ�II�-If�a.�I�r�鄩�C�]�����֒��P��8H*�uڭ^
�=����W��Zq4�B��H�ҕ^��O�1�����n�vZL�0Y�sUR�A+�������(�Cfv\z\ؔ�V�7��_���E88ZΉ�����#O+μ��i
�V����8���}r~g'%�wǷ	���{�y1���̶���{�]�XA΄����_�Q�%�;2�Գ����S�B��YĖ������v�U�/����y�0HM�b�w��'��Őb&q!�Ӑz���S�h �6@����io�JpvN^v��'��/�BqN���l{�idâiƈ����r����1b��!�`�P�ߪ������&MV��3�i)'��Æ%�Q����1�=Y�'�5|E�o�9�nŷ��'8<_%x �����Pnܕ�+��ί5��r�.�V_"h�ml�BV� �:"쮻�o���|S�գ8�7���f�M��'C$؆Q��q0�A7#����!�-d�}n���i��(��7bV�7i��J���kQ�#�׳����^��$�1��2�{d.��E�2�zձ�LPw�����N=
B��$�@t��gd}A��(�� �S�A�u1pOqDY���@̍k���B%��8֨
֎�6|1�.V`k�����#��� �(n~d��u[�S��p�E ���r��L#]z=�L��$�qd�(8/ncQXSB���"n�����Ux��3)T�V�/B��Ё���;i��9����<����d���5��
ޜ�FW�i{���D�6�����ыw�>����݊\�5��BG�T+ ����)�s�ǃv�	՚���������6�asH����Q��rܔ��_!�=&�b������]Q+�˲ˎ�_X� �x%����,�Hff�踢��I�.�4��* T7K�}[u�Y}�gc�0�곞K�ʁf{
]����]8j%�9[�ԋ���k/�l�a�d�	䨷>[̆�>�]�F�_`)=���-�|Ԑ	�Z���&UY�\������Ը1
���������J��{B��FS$�I�'�����`�Nab1k2w�3Q�lȠ�bX�c�=5�^�(�5]�+�)3�j{�s"mif.���
{�Mb�&͐	
$�[9 .��v�a�b�Q�{U(D؎��j�S�Oϋc�-�������ї��5�
/1�0���������0Ǜ<b�D��W�ΙF�&�a�6=�?�ԅ����5��O��fϬ���}E�]����/)�r�dӪ�����(�D�U2*�9�[MDH*,G���	ϗ����9)��QB�Z>��GQ�<
^���b"o�΢0�m��+���,����0�]\D��E��N��'Q�?ڀ�����(���0�o�����:�3w��ճ��Y'$bnN\�F�:v�|YX]���ˣ���wjm�5��nP1�|��d��-�B�jA�ww���O��O]�)ק6h����	�Z�'�t/ZP�Y+��s~:�A�C��M;�GQ��E/A���ҙ���-@9��>Mrl0�t���� ��|��胙�MDi�a���%`ew�U�NwN+yxj��̎E�[��0D,y�5��0A��ǿ4
5� ���Jy��X�#Z���f�w�Z�rf�D��e��?pxd�����$�R��a��E6�;��׵�]<�==
� �X}<�����L��@i�9m�Ńw�1�c,'�sn
�����mn��+�=�-�����p��}����܇��yZ���vO2\��(��yU����R���rؐ�����o�16<jNP�d��u~z�@����a���pJ9���p��#�l9E���Ė�#r�?
�!�,�|qǲ���:o[�yq�2*%���:십mu�����.�pY�Z뼽�����
��+b�D	�/G��?��h�.Oݥ�͠��53�>�-����2r�a��GV�4F�Ц�a9�G��*��T\BuF����t���������J���Y"ʷG>�H]16D�*�e+�Y�ˤ��П�^D�|�CM��&��[�f~58���d�f�j��ϟ�����0'�ph�d�
������_f�H?=�3}E/=����L����j�����	���������񁘣�1x�Q�ۅ�o�3"�Ν}�A�h����C)��1��&�}����
��YwC�@^%���jdJ�-&��\��+K�J�c���0���R��`Ȍy��O,�O?��\51;��&�z�����Q�H��,�3ʞ0���搵�/{52B-�� �Yx>�4Y|쐚2���iv��<	�z�n��M�l^P`���&N�Q��X������Q�s;�í?�\��[�����P�{w�H����A&���d�N��7��dm�K�=Pe� D�$To!���(��.���,���v+� ���@{y_�`��PVv2����#n��`�X_*�;[���6]����Ԗ��D/�T%���4�2��%�D�FP�"���	SǤ�_�����c#�.���ΐ�*.�܄��^]�Zk��<�$l�!�N&��i<2`D)� U�I'��̹Į�nbg�jJ�����>C:e��Q�\K���}��F2�u|q�ʔMf�`@�_R�� �?�K�,_���sb��)���I�tJ���宽tʻگ�*�UC�gʕ*��������O�V|L'Tp/����%3���-~K c�KT�ʛ4�ݿ#��k����Iڼ�9�|�z4N�D����H-ʜ��?��K�d��i�p5㨓�[����?�
X7
)m��-����޸v̝�M�Xm�ݎ��&I�j�L��K���ެ��9oܯa��޸�Y�}���.ׇ?V���/��L��5U^x��7<��9`�4/���,����G8b"e��t�s��$�/�-��U|]�h,�!ϘB�bfe�?�[a�BC������ƙ��TYS̟���K�^&���1d9 *A)�U��Թ�s����-�V ��Ͻ�[��f��dm�Si���3�9�NZ9�B��"0(fXbT�K�-f��(q���h�[j������~
ڣ�4��5f���Y̦�n��X��7��9"�����VK�jZ=�;m�� ܗ>�T�\~��E��#��W��cZ�z����WdnlG�>�- <���s����Q��t�ȶ������w	�]+>M��]f%"�<���ذ�8~�?��e���>Z՘|)�
���"ǭ{	�+����w105Z���c�s jx�C��"[^޻���,z6ǯ�OF��pu>��!-ֳyevs@��`�/W����ʰJo��2A.i��v#F��Q~�%��Q�e�߅P�`E��k�����
����2����:��~$Yr[{9�s6Mj4Fva���C�.�	�ق�Vk��Q�)�J�ݲ�] ?���M�o�9�hK�}X��������*Q���aɝ[N�츩P]x���jeiu�Ӆ�:��;�Z�$]+�r�;�(	%8�MA�>QĞ���/.|�]M�ܶ�~aȬ�-Y�cy��i�Er�:�6=ֲ�;�Q?���z�ݼ]�֌�;L���`�n�M���$b��6Y&�<�V�|���|g�F"޲���o&7N3�#v�|6A�G���C���,P��;�j����5j�݋��$� x��ʗo+wC"d]h>�Z@%�o�ט�!;�7�����
�|G|���9���wv� �-d��;J[Z���s�E�~g�_)��;��\Cxt	�� ��Xn��͋���T���%�S�==`���L��D��@���J�F�̭sG���j�_t�boo��&�����!c���:\H�oت
F�t��s�@Yx*�:����=~�F��;?�8�О����;���nX��nWqʾzp��,6�܁H�e�|�h��(��CL�
�s�7��$����ܱgݞ,���>k�<,n"3��_��T�����H��rp�%O �}�UE�t�򠇲�����D3#}�3"�J�T��$��q����}f��7M>��^e'v�k"���-���NKصeN]�����2���?�D�����ӄܴXc)]3�Ч��y�ؾ�iܿj� ��$��t�=H�CU��ҽO�pp��)��L��=#�|-�wk~�@�Z�z����|靕AݤPÙ�VK���.Z	��R_9�I�1��'K~�$Avr�T���YL�rA�T�-i�5��_ޖF���Y���3=���c%�2D_S���ܚ�m�D�O�	�I����Z��߰����3u�m�fͥ/��j�jğ�|Ok~t=6����l �x�M�*BO�'3�l:��˨���~ۓ�P��v��7�Fz�Dv�-�VY��2�8�@Wʵ�ņq�\|nehqdNݝ���~	���w�=XY��,�l�]��u��U��|���Y� ����3�l4u�z=��(�w��8�YnAM�|W7�8"��YJ����e����e����A�ܦ��wU�?P����J��w�v1Ȯ�y� ��������:�`9ţO%�#\N��b�{h��%�/A�!���,���dxE�Ƒ�q<����%�/*]�=�i���E�B��\�{U�o�,5C$)�ǟ�|��� �M�&���p}�	�دʓ8	5��2�,kb�
�F�3��i�:r�Q:����T�>���W�����L$�K�e��*H��AhI���z�K�1�A׬��
<�J4��$CU��64�?���9�?�z�B�K�z.OpȵI�BL��(�L�]I��v�}�� H��#T� .|��,4c�z���M��;������� ~��{�Eb3\�Pz${�:1�;��R��u3C�O��Cj���k*+�)]ǘ���k-�Z`v��/�O� �U\#dK��L��	�}�AB!��ӓa��`Y�[~2_Vó&4���^�]Z���H���|�]����X3�vF�%!�ᬍ��e>���$Ft�y7Q�v��0�0/S3Fz�>��~�u�����
��d��%��d֜�NvE�
�s-LEC���#N7]c���
���E�N���A�	KrVh�G>��ڿ���2��ϰ���Ǔs�1������̷Pz3��g��u����4�V�qS�n<MBn�0ّ-��!2����W����bs���c��k��Ci{Ӣ�Q����]�6ж���������?�ڝ�Y����������r����jzN6Uc�w�4q���F��r(e�Z�b�*J���_�A,� ���'���u#)�-R����W�M̒G�n��n���c�f�¥b�S�x�'U>�'
Q��H�|�|骯@�-Ot�ʸ��̒^�N���KÇhD��9�S��N�Hd��B�aL�oH�2�:�ǹ���0��A��i�9�1���t��!_9��1�Y��������ZU�t�N�b��=���0�u���'v�N�S�1�-[���^�ǐ�1�)S60�R�4�$�CP�;>����ȡl%@����䉦)�c5�޹��������BC'�:�?7��5�؁{/^������@�J8Nr^�W@�cq`��x�=�b'Rb���?��@eĦ��� l^ �����;4N$ݨ�=��{A�l�l� +x�F���EJ�{|~1_��eh����z���V$<��e�c�'^��Ht��k�i���R�=-��i{_*C�^���|	w�!��r+��5U�H~]l���娈����z�!����"�f$�َ�M�[�wP���˶_�Y&0o���N;`e���r3���7��z�j��tHk�.T�]h�K��kv+�FQl��Q���#B8H��I����ݭ�?����Z?{���J#���`G�̌^G�Ń���y���p�Ci��^�WԽ_״uuq Σ�\+Y��b?zr�u+�
�Z ����@��%a�������F	���O�n�P��Cd?r��A����+}1��ր�����dEOS���Kr�T�����r)�8���J"<i���F����)Y��V{��@�=�-c[F�B��_�e3Q�X?mB����1�L�ą�81��P?�>c
Y��<\l�-1����8�q���֎T�Tc�^�X���iV{@�x�8��U������>ؚj�7D���I�K4���C	�oOԖ
c�\��Uu��Tz(��	�#���c�F&���x�m���V�u}tZ0t9V�ڌq����U~���D�L�ڍ��xM�{ �7ִ#�kb
{qb;\k�]��tS�?�ɹ�'�I����l�z��hKy\���o��98��)�Nk�i,^N(�W*��(�G�OŬkߔm��@�	��f���;��Pמ�=�|�#�׮;+����ge�N:���^�.r�w������6fN��f��`��	>�X*�M��~(����$�x���鈗J��OO���^j��GD�� �U�}�� 3�~2��d���w��R���$N�0�A��9��>9W���6��\f���������sr���5Sʦ=o���c�5���˳Y��)Y�[
�=�y&&�>���΅H�sX���Tt�Jħ��6��q��P���&'C_��h{�ƿ��U�~:�T�^��\��!f�<;��f¹���k�g���#�:C��m);��p.��i̢ko��s*�2G�T@O���B\G��7�Y��#=ݑ$�C��7���	�M�u5�s����Ql�������)�U�f�	^`�@�x��^����3e�K6���ВϝL\��Z
ӧ������vo%���>r���Ϳ@3C2��d��z� /��������(��la�S�rPw��yɬȚ�ʆ����N��3�LIؠ)E��,6ƶ[��c����Y!�y�xi!���	R���?��V��,�C4��ݐ�_���[�8Ėc���(�.a�����3�2G�z��Gh�+C�m����=�j^*\rI='�X�[W��~�����Uq�����<��SDT��p��a�A^�?�Nt�X�l�W��t���&d�Iq2��	�	�N�qwIRj֛��-ȐB��!�`÷�o,E*I��W?�d��Y���}�
���y~j��9��E�Kce�=��A����#SN���*]��c�K π����*vC
�h���P$^h���2ȃ�_ ?r��э%7��4`�R�-�����	��]�bh��f�Vp]<ZZ�=w@�OiHu�*#����t���Τ���q��7l�b֜>'�l_�|�q��7I&�# ���[�/w��SPsC�3�kQ�Ds^�V��
F,���:-vK0�N��ZĒ4M@���^�nE�YxL�>�-�N��uo���Qk\n^���?h�I��o�7Jy69���Cwf�����q�m�w��-8Zj��s�P��3�:,��O��K�]�][ׇl�W�X�d�A/VkW��B`��w��!!-��4K����3e'w��昏m�?�-/:�w�UbO1TQ�;���R�I�y��!��Nwa���d�ה����KY*'�8G9�C���N�	
���Tcp��������~[R�D@��5.(JheK�q�y��upQ�K��� ��8�JF0](uY�K��=k�X���pZ%18ǜ=I��޺�!�v�?�������Iq�����r|�I�J:�OIz:j�������٧~�F�h�H��8���zs+�k����;JX,%�Y��g�t��=�Bū�v^�ԭ0�"K�r��"@�?���	�iֲIǿ�wﮎ����oj	��RB�4�ܴ�a������K8uZ��D��+K��(�O�l�!�'�t������*Pd2��l.��I��8/��W�")bUm����M7lA"����x��R�J�x��&=i�Ņ� �S+�[�Ю#W���@\��X�^����;��1?��GK��P�����:VU���&d]���(��u�Pd�$l5,�g�z�)z��r�x!���})`�oJ΅{����aL����a���<M�d��y�<�7�ly��0�#���c/�\�$×��E|�	;3}����i!;�G��4�8�p�~�bi"������"��B��qN,]@^�}V$	X�Z�5Yl�D�d'
7%��$�JCG?��	��,@F�eY�N�<eG���f$hA���R��rE5�Z���<�M�&K�BK��xP�u2@������g{b���P���g�
�g�C�2�lnd��aqr���)�>9tpBBm��:HVth6�}|�Vmt �]/R��S�0"�:�3��x��T�G	�f�n(j�̢�k[=*���@�_�[�@���V��9Z)ݠl�2:*1����5������-�O�X������zq���>t�d��H���	g2���Ą���hC�ݯ�Q� e]�K��j�x2�;�ʒ�5�jŞ���.Z+����`x�5�d��A�B�
k�3#R&A;��y�������0�l+�&<L7�뵃����+Z�0�A���~P�S3�������_�T����F��^���ꡧ]�<�ϬQ��:��e�=�_�~��~�_>d�jz�رy;&���V�J�XN�t@Dږ���T�0��Rγ�
�:%���<���EB��Ub�@3��A�8n����46�}n��BI�&�S,?� ։i���m�*��Z��\�8#��/p���K->8HK~X��n�e�;���X%�Us˦��M���{��#V1S,��"�ZoW���?{l�\'����}��B���c~S�}#�\�x�Ԫ�k��}ᱍr�5��!K�k	!��@�E6�.��k*�ة����W�Z��p%3��I��I�d���X���SAzN%S�s�O
ǽR��[L�����<P&^:����X�����˿�B�H#9��}��w�a�C�PKZ�����._��<�OB�r�;R}���&.�TX�Uo)_Y8���U"<�i���;����e��i ���*�̞6;g�C+�:
��Q�C��#��uLG?�[�R�"Ո�p����p�gw=]kp�8 :�I�s>�ƑV\5�$cdo�!F�����T�s�������e���\,W�H�Ýs�k$"����}"i��$z!����[��>��#p�!� A���F_{�jE�;*��V=�J��Ɉ����U"���\�H��ݗ7���(j Q�ک`.#Ɛ'�汒�|�|�u4�]��7�����rF텒��:��4�K�0A�/��*�Fц3�5�Axyl̨&n��`b��ǎ�K<���{�X� �ܾ�rF���F]��7. �DڏN�?*`���Ƭ$	�D�j���ګ:���lp��b���ߤ�|�7�J�g�]�{�<�5�Pg-���ωw��[,@�ܬ����d�E�Ln�-��tu���`�)Thw[�Z���>�����j���O#[�P����t��2�Rf9R�H^�n�3)q��iy��	)�)�]� Ѣnr)}ۆ�i��W_�B٥�;D�-�ߘ�-m��L�]�4�@aq��ԑ��2�40�a<I7CH�{�o� ��v�R�7^kk§��!����3$��: �d,}�,�3߿��E^��"Z�r�ۄR��O�b��}�ts��7�e����b987n�n����=>��ț�YӮ):/M�/��mB_�S�n~[G�'�T�e��ɧ�V��!M�"���^˚Q<~c��ػ'���M�]i��B�<���֑��'3q-�U���Hf7gQ���e^���l,z��8[h�a�#=�#J���#�;�YA�"�����4OZr���5;���j��;][����Ff��L��#Q3�̢ź�h �� ���>���dm�D�U4�z%�`�s�L3�p:���D�r���4��6!ǥy��F�9�a���d�y�)0��_�fPOf��P�~��/`@Jo6H���/�5ꯞ��gq����K�4�[�i+.j��N���Q���h΀� �������$��^Ij�s�u��0�qX�q����r�듩&/t39#�or�EV�O��2�n�܎���B$����O��.��Y<�@���_�{YY�VG$����B��t:�����[�9Z��B{|<X9F��,�l5��_EC�51��+��>�
���hc!?����ddǻ"�T!?L:v�З��n���$_
���X�m�|Ye��@�K�g�j���PE�+�v�W��hN֑�,��dI��| ���s�T�]��nx���Rp�r�v����hB��lqƴ�/2d��h�iwAC���jDf ���"H2V��f��yY�,7<\��]p��}�J�S��V���� b��W��
�~�m9�'b�`x��rb5'lV|8��rkly�Ա#i��x�>Mo��De��v9-��|s�	s�|��/��"C� ɹ�_�1P8�1ᇋ���H���*��|�Ʒ�_�/�#�膴���Z��}�'K*�Y�����#wq1f����ؘ=���S-�4�68�h�^���[�̳Z;�t�jQ�]NI����ե�,T\�����$�'����ߋ�C�L�C���ζ��|.�*[^�d.Q�6B�zC�Sf���a���2K����h"�kR�RL�>�$;�+��Q�~���P����7������l�4�"�5�L�c�q �L��}��3�WE�������KJoF/^UeW"+��	AZߏ�9M�����0&+�]1�<G�����~�*�˗�J�4\�T3���FD�l�&�k��Ѷ���ۡb%9�5�D�q=�c���҄Q�y�j7���1��<�j�t�|�Y�#n�X��Z����'��#���5+�'���g�`���K�����BH� WV(ѕ��5m�l��B���x�>I��g�E��]�A)�&��~���U�)1*�ು:q8��fx� p�Y����mDA���]�o�J�ӎ�Xe��Sb� "����>#��g�ЉI
��Cz �:w�S3�]�ìrSG��#󄷟/	�:��! ڸ�<)v�F���6B������H��{�B���{���V����e� 2�c,���j�'ի����k�mL�Q�rF���v��o&�VX?�NY��.qyDs��̋-v� M7B�Դ8�g�>W֭#���T��n&�0�w#s̛��|/I������A�}�F���3������dZYp���:������`���ء��&`^
����=r�����צ�Y6P���9�n�5L�^�KR1ԥs�q �`�kW_��:Oe��!��R��@*<l�y��D6gʷ�仁M�]	t�y%�8��Dt��z�Y�����������Ұ�&5�����Е�z��<h��O�ek"#�L�(*�BBSE���q�m/��ŭ�0�x�Wm��@�cсP��,1�ӈ-O�[]�ٜ�7�[��S? w	�f�>A��&�-����~�&ﭦ�U���g"��D�L����8��y�i�����ZR�H'�4��@�)���0J���u��d7��NS�%i��q����?�g����|�t�Qn�B	�I
`td-�,�;l��*T��4]l<F����CA�����e�.��Tg=*���i{�����+,VT�7�`�̆"�i���'(We��`;�1�ڋ2?�u6ӡ�z��q��14�e���#�wS�E��1d�F4�pE��S��f[t�4�W�2�F1��J��۞c�K�3���5�zq��l�OI���u.Es��]�ٜ���uٽ��Z�з�g���`3��0�B����D�G蟂��c�z{J��r���o�r���/�c]b���=���
�)�+��<�*������������0rn�G�NTN��aҨpƿ���^�^�AЦײ��~l�(6��.�9��n`d�a��3�)C�ָ�|���\����	��?圬��&�A��v��a��_L@]�~��P��H �4����:�0\�Q�Ip�(y-2�Gs/��m���bs�&U2�7��-c�o��z�Uo�YM(,�h���T�h� :���Et�6��p��^ri�X7�����ߠ�/s�����G��sj����A�4�q3Mna��:	b�f��\ �>��C�`9#2A��C|���I�o��0� t_Y=��p,�����#qL����>.B��$����34�Fǹ�z;��
�)Cw��̽�9��;W'��]�����X�x�U�R�ڐB�Ҙ���Α3_T�p�o|t *r�o�#��[���"��8z��hZ\�@�����f�����	�<B�y��P�y��_8C�W6gǇ}��'-�-���ɤ�r>�=��R���r��#�Ra���|-��w�#mD���}�JW�����}M�g>)Fm
��Z�>�t́�1��S�$1N��q�VJZwlBx3�X�yX���m�&���Q��%����K����E�G�
{\K�
�/�D^�1�?@��	��c�ZG�P"�8�8E�b�	�l>
d��Sy����I�E:�)�<+�uCc�~���ҙE\h�n�2���G�{l�4�}�3Z	Kv�ĀN,��T����&��2eE�㐝�?�"��Do��x-�:�3�Qɑ<�P��Ѣ=��Pӽ(Cm���l��"*C�9�� *��y���#��{����.�Ǧ�@��А.~���bg��&�
zD
���;3�l8T��|l�//1����*��D
h���Ŏ��noñ �(9���w�ǻ�uFR��i��5'Tw�j�� q��Bn��="�E
��t�j�E$������dre	���g�-�C|�r!D)i�FK�+���웨�|��GDѿTlB��g<fr��P��'�� ?���l���o�l:��d�']�/�J	?�ԁ��0�Ԛ���
C,����o�|'��_b6�x��낒���^xu��Uiѳ?�;�Ok���#^�����ho�NWQ}*�)=�[���E=�YER�ŧ�0�dދ�;p��� �p[��U�*ky��G+,�q���I ��7}�썓�r�VvPP@@�F�A�\);N�7w��igV몥xxMۿ�/���f~��9���2�8A�
�2M�UYS�g'���_�����2��gg�%����'�� ��h�M��3�x��yMV�&�����W��8�����Z;6�>$��b��&=�~�А cG���Ε�¯�:�H��5��㼤�l��;��x�M�'���	� ��k�jF�p9OAU[@ǔ��WH�W��n�?�
���o0�>���4$PN�vk9���ǚ��( M(�M6q#ٳ�!^ �=�#�A'�F���a��xQ��d��i���7�*Bd�_���&��y=��a+�d.��HdI�ۡ摃J�םH9Z1]Ƈ�x�#S~��6�������7:��8�|��-�D �7s;J9z�hu���j0[c��D�M��zW���p�]�n�?�_(4/o
+�>���}hBS�Ul�_ k��>��$����=����:e�kS�M/�5�YZ���ւ1s���l�>�>�J�d��<J�h�,+ā����׀��8/��Ρ�M�5�����N��NSk�a���C�g�+���,��l��l��k�����j[�Jƈ/�,���b�E�����y�"�
�k��������#��s�F�U� b�|�~�0JH �7mR�7f�����Pr}G2" �����%��۹���"ܬ�#���$���t	s��6G(S�Dr�W�;*/}�.C��U�.S�v-���m}����7�6�c�~z�G�����8$g(F����8��ZEN6�b\�Bo�2�K}��n	v"�Q+���G�������%�lzw���F�<WC\[�ZU=\�y!��2w�7jJ�����֪3f�NW��vC!^y�q-3mr�9���U��2{��? ��f������z�:穗�P�tcb4ξ|�ۜԹ5C�tXd5:��S�����)IA��h�;�҆O�>39�9���X��m�y���f�ѕd���=e	�;W���^�ς╧/���0��{�.�4|���L�CPZ��/�Y�4���?.���,/!�ӡA�����Z���r P{��GI���cIJr�${��ZW��A�h,�(�7���zaZOiLv)�#;6�즆õm�aj��H�K";?���#6:�ȁ�i6e�����!Fu�zt�7��[�Q8[�i�i�b�:�H#&��l%Pۉ߈� K]E��QҾ5����N�0Vʥ29��H$4k��M�S��4��Sr�|��n�vB�2?W�i�$M��~@#��� �C
�T��������i|fʴo��Ě
[�Sx)sE'�����߱��$�1��ld�1pj:���h�g,Z>$E6�py1U���w���~7[��$?F)�q�� �^�,�lZ�q*�#����@_���T����fFi9Ot�*}zAz;�u0F�嶠I�/g_�O��`�t�X�W������1����\��q��%��K�FI_������g�>��(�$����Odb�Om������:O��i3�S�1��}qy<  �\qx8�xwn���ѧ�_�~����~)��[�(�#O�����0�u՝��6x!�6�N,�.Y�����ϗ�͔��{��o_�v��_� Q�����7��p����<���X��[��
r����\��u�aa@��)��*�O��I��
6��Z\�;SWl���`�����fUc�� ���T�M��IsE�6�9���ͱ���/ J:3^��f�rN)�=g�_�!JP�f֙r=�3ⴈR�K���'��.�dJ�W<Z�<fMK�W�'V+��L�X�L6�EN,]��I�����hx�u)����|���KF�C�JO��e�i
���T���ZdCR�q�D<ε��a�1J�zְtW$Č��Ꮪ$PO��O��f�����OU�A̦%��n�XX��$~�����J{�vydL��o�{U�	��>�Tx�b��K���G}��,j{e̡*�08 >Ld+�9����/��b�U��ZK;�����.ʟ�*����&Ž� L���?�c[���A��F�)
g] _���Ȍ<\�y��0% �4Rl���Woԇhf�?Gߛ��k�3� (�e�̎^le�F�9�UJV�r�[���M	�-�(�U�ؗ���E8����i�)���]i/�5��H�%�A$(��K�X��8�����g%@["�!��E�O����uA���H�0>w��J#�f�M��f�g1�(t%�P�W��;�#:�m��⍀�����!/�z�&g��b0�����'�m��P�\�e����"�\�m�n�˄��`�TB�f�C'����X��ZD3��Z �CQ�Ճ�(��Xv?Y�97�]�{4��2x���!���f#X'��+�9; ,>o�:��ӧp6��_R)Wɦ8�Ѷ�����������*�N�~����-3�Z`(5)�����8�X�©ruK�9_y>��_���S`��g��٭+Y�%Kwl������?��E�G��@�*٪6�����g��g�4����� �	�3�G��V>�'�N����5��u}���{dq�� �0T0^�9_��#���L�9�Ǣ*��P{9w���X]X����X��:�b��A�����S�m�	�u����o������$Ƴ��1�t�7[���?�L�9J��Z4J�j���X�}��'��M%HK�8>�s�@�V�Yv��n��1y����#�eCr�[���:�m���P�����T�51ġ�)�/�I�7��}3l�PLNp�lE�*X^��+gp�6��3#������r�>H+�n�IcL�����l�>�l�m��{�̜w���%�{�
h���5§7OR�uV)�E�p3O�0��ž{&K�:�9k�j��4��5.Z>���wh4X��ƶ�|�w f����Q�龼0SW�_9zz�����x���=Ch��OZ��M1*o�J�%2@	�\J��!�H�z���Ə\dfr9ʈTS�S���?贎'�I�x"�cqb.7r��a���D��0��_�"J)\T6D<4~@`�������未$i��������ڂFp=4�$�[Q��0���>���[�U,����Q�B1���N�?Ie���� |��
�&��48l��E�xk\<wV�
c'3l�y�G�e΄8~TQ����` �Ig�����'�'�����Tv�A"q@PM��-n�(���}9��d���;�ta'��n1�wIؚ��X��Y�|�4��3򌹃?��\��<�N�c�;+�dE�K��`�<+�
����F�*�!�J���@6��C�3�-��]�"�c��O{!����qK-�ޘ�lE]^4o}*�Y���OK��������zMg���N�4��mkv�o,Ԃ�Z�e�8����#B�p0՜R��1L�����^�HZ�0�������|������_&W�}�C&�u���~m��F�`-�U4tI�΍�?����7�(oI7,r��ؔ�ϗ���Jl�M2��i�_;Tz?�a��b��T}�)�C4�̄0�cH�f�R4"\Ŭ��.�}�u�歵��@h�����u"�0�TM�?E�ԁ?�xt�UeLT1=�aE��Xfox*�e&��`8^?��ӆ�/�}����\��&Y>��q�L" �7�7b�cͳ��$-xTԓO�eZ�����{��j?d���	Won��	`��R�.�F�g�v�`V��T�!�L&6���&�,_b=�Ty�.?�
��ed{���ݼ �16�p��,Ȩ)�?�IQ��f��(�\D)���ѳ�*䇑5�!(�U2o��5�D�Γ�j���V�m�#�s
��? '"��&Wq�52_N��~����H�11ч�_�쎎}�p�Q8���F�9�E���ɺ2!=b�uAK~��>��w�����|1��Z����:�~8�TVbjLr	�f��	�1 G1W"M�_��J�bRO�r�M�	{���a�Quf�����aS����#��I�+-��O+�K�e���h(b�2b�CE���Wd�@����B��4k>'�� *�q� g}�a��E�����:"Z�����:s��%�9���"���EumB,2�Qt�ж" �W~=�2�.d��i�a�y�#����N��p,�R��>=^X����+��\; D�2���S�*��I㾱�c���L��*��_��@���3��vpUf�6����rX���gH��jDΎ���1�Ub��ۢyP��a��Z��������U	��;��	�&�y9��Y8��"�y|]kO��j8`Y �P�Yd��إf��&fv�iz}��'1&��n�����|u���Yǹ3�����\��=�Ȱ��a�A.^Tȝ���=�G*�+��2��ӄ9oc��R��� DU]�Ks�����I>`�.rS]�k���@eoT����\%�K��]�ǥc�����/!�����@��i�Y)T9��L�WXY�%�P�7�[3oA���h G���x���R� f����_�6��\1K�=�(nv[�C�%�����!e���,�*0]� n�d�B����ɕ(K~:u��L!��kS�l�){a�cʉH�'��m�}�����ZRY=���+IL�
/Fg���dr�zh3���=^�n9����Y֞R��*��"�bCE��%h���j�6�3|m5��]�����o�A~����r�-��:�}���/8��Th&�i�+����=��*��o�[�wU�X�B,�BƝ����c�l~>_�N�y�B���y�$��u+X�w��.|�f<�{d��Fj���O�IMo���2��n"Җ۬��y��˙<���.�/��{Պ���7�Nh�!�u�M+W\1��C��0�-���c�uv2�/N������/��._�\��Ƒ�����'Y�ЙnV���pGLg8ڔ��PEn��*o0�A�(,��4�2"��fHqKM�'+�f�z�<HtR�]�{Y`������p�z�AI1�\�dg��:�^^�ԥ��'B�(-�%Z�����`�E�6�2�ۂ�=c�U�~��w4Ek�R	��`&���Sr��°���J��}������t��q{�G4����)Ui��pX�CN�㸌�=�C]5�<⋓C��Z�s��{�2]�Q�љa64��e�|�~dcS�~���\��.Y�_O���ҹ���T�"ڭc!�BE�xaMB�?	��fI�r�{K�5�昌�����Gp����C#K�ڟ���
� �[Z�0מ%G��&���k�\]g^HT�b �d��]E;����X�yWbJ��<vг��g4�9�wS���j�P�Wrp�P�s'���ϣ[SE�FqX�AB�	���5��Q&ܓ�KQz����,�����-�d}�uk�[Q䗀�a1�y��1t�&I>Ȅ�=�H�x!�����M�`kI��qئ�����b�����Oc�#��)�x��gN�&OM��cm��d�u���]�������l���K�{��Oj��n�[�jͯ�zܹZ��������I�G'WI�����TM�￣o��Al��>��*�$��F#�շ���S�^��P6à�~��UC��Ӓ�	|j��AH�z�� �������oGB���ϥ3���x�?��8���[��*�pb�v�������Ċl7�HCo>��k�K��Dђ�.���Ї��EfI5B�p.�͋�d����q�t�E��S��BK�i��^�@N�(�u��X�+A��&��ݏv
��RAp'���}~���A�U��*�#5�܅��N��~���x��\� lJ!��S{�w(�aK�ɚV��Y�P�iށʳm���[��Zr���%���G�|m�O¿ǯ���3)�"��B��C5�6�a�v�&��ΠC
�k�Ǣ�C����vo6O��Qrl������kG:� �������Z@!u螆;/�h����/D���N �]~6?7�X
�1` �h`�e��O��`ְ�yK36!��a\NA������R�2�F��8�v�xDO�j�m�b\�JG��#��"��� ��'mL�%K�Xw0�u�L�Syͩ����9?V����Q� d2�M#�7|�ɹG^�����"���$TxT����	��&�D�^G��ׇ9a~�,
Ɛ.�b)�C➲_��ng���	�Q��24�t4�(=�$nX�3xQ�}-~	���|�C/ҽ��@D��D�e5���kI������&oob1�!<o?�4�DK:��í�>�ֿ��<��<4�X���2UG�"NU��E�g��?u�a  ��kԣ{���=u��+��>��.�t�Χj�k��xl��X<h��D;�ʻm�φ�*~�v%�g�����0*ۣ����E%�Q;�hZ��F���|���T�����9��\��	w��w)d� x��a��`�mSu+�Z�V�K�����o��'u1J��G��q���K�>_��j�;4��ڨ}�]��	݄1�B8G' �^��α׃�&&q��E�ۥ_��٭N�A����������I̷pQ&dvO7�;T;絋��:�{��qt��u�
@ے�O����C��x���L`:�m���{��	�LC�S�ER{�2҈�N�;����q��"��u#��!)��7�=Q������ Qq�:�@���uD�ϊ��c͜�G�G���u7����C��Zuz�|Pw�U�~S�b��|v)��$�����y��?���6ӌ�q <��rKl�	�*�G+B6}rAq:��f��h\��#�H���^�����=�����8�bɊU��-�_l�aB)qR%+��������\F�8���w���5����K��E�-آU�~B"z���J���\�x�����ј*��S���6�3;�a.�)$~������M�~�jԃ �#�ۂ�Jb�4�a���,��q��o�pG�����b}͵`���`Μɰ?����]�c�t��ᏪC�L��P�k+�>@��
d��!h�t39����N���cY��@	��+vw@^˂d:COr�	�*<��#<Q�x<^��`"�(�q��M�r���±!��L�Ɔ�]^�}����f�Q״1Zy�&��ɱ��� &�/5j=���4qB	�$���:}E�y2q�ŏC-��_>�ƛ������@Rxˀn)s�^���0�&=�)5�H[����<c�� �)B@ ��|���U'���S���J�ۉ��:*١]�q�@G��/�ޅD?���\�"�oܠ5#-3t�j���	`�W�&H%��N����k�Q�E�on��6��S�Q���(O��6��<��
����L_�R�;���p��3��i��Q�Љo�e�ц������m���T x��J��������b3%o�<�����3�"�p���UC�.���³����!��W�'Ȁ���C���������wg�v�w�ٞ��X������EL(&��.q��m\u��X�#r@�D�݃�-�|����ݍ�L����(���~�P��(�DZ�g��g{�����nO�O%Z�H�c�N�T�Oi\8Fu# �(8@u+|��;T�$����K�<`�&��8��Yj�^�r��8#��<�S��\OD+>A�)`YYM����Si�Z�"��T|�P�gY�`AX]�ц�j��-�!�m˻՚C��%m����r�A���IJ;�{r��NM����?�r5Q��N��7p@��W��A	1��Ծ/=K�aAy��6X��_h�!6U�R�@$�6�V�P��5O�M�${F�|��a{ghV�dd  C����b���zַ�2K��i���Cڤ���)9����pe�F�Zc�����������p7X;�l��0���2y���z;$"	�<k���$& �W�!(���Yм�3��Y*dɧa�r!����D��zG�Y{��i�L�����E��a
v��-VF � ;��ߥ�=	�u��Dj96d瞄%�<ϮD�-� ��{Q���L��fA�܋�+I ���V�.�3JJ�+�jO'��i}�������b�w~��o�l5v�G�
����NkgwZהg��=�S�u��B����բ4l�����yT��r�
����s���9L�����#>'�=��5���ʬ�VJ1@P�$��vAj@-�/�G6����we����TM���It���4���4�\��i�-�Er��&R&����{�_�U���LØ�_3�0��<Q���>2�Rh^{�ʅ�w&kW������!MY�1uQ?����G$�U�ԁ�� vI^SP`r�IQk% ic�f1�U�����h�
2�6��*S
8�!��'����^l��^��'��&N/�V�e���3�T���i���d��A,9��`D�+Y�$���m�D�V�,�V���M�vV}?
KVW���H��j\�*�4m�[���Z�Y�kf1Ł����s�LϪ%�߈��jA*�߯3�tY2���-~C�4pp�J�N_�Fg���3s��#R����PZ������6!��;V�G�C�#�n=W(�d��^�}��QNh'�#P�X�5&���R��Z{O�EhЈ �&�'P������+�0&��i���5������Jb�z�홤�f�`w�U,�|)[I���P��y~(f@�]���?�[f�}G%H[ 9�4��t����\y��,�.B3W�(f~��	���5D�K���}?Dnb�d#:n"%چ�VI�k�X�[�j��\�N�?�7X��I0�&��'E|ra���w���\a���J�p.�����L��@!�-w����g��[���ŕ��u?��+wG?��?y�2W�%��`L^�y�l�+�Iw�q�J<P�V� h�)����û����
9�jEL����AJ�$f��3�@5�@�N$�q~��e�ى�>"Zn�.�MW�&��'Bυ��*���jz���Ot��n��a��6���ےU�\��A6w3���a����'E���9qr׏;=�k��P�SO"����ViiH��*]C�	X�	G,�έ]m1�f'�LMܹ1�_wm�耣�h� ;^�ѵ�0��v:��<H�J|\.�f�5^���E�t�q��
����lG\Q�� �2!�Q9��R��tnw�a���TW�Ҥ�x�}�h��L��v���	G]�t�Fk�D�n��'�L��f�UH*��1B\��u1��q������R{(��z�����*ǝ��TQJ)�m��t������&}�L���[���t��zF�`����I}_�������Tva-�"�'_��K�d
�,�ljTѵ���,�&����.7��E�Ě�0kk�b��>])ĩK�A,8g�t>V�x~y�\`�ҝ��T�[�$ tÖ1���Mx@8�.s���Hkt;©&���2�B�����as����Ź�Ω�t�9M9����%5bןź+>,��"=bO!��v���^�l*���&�cO m�xfQ�	-_��5�q�T ����/<&l�F� jLA��@���%���(��_+&q:�B��	�x�-�eVX'|��3G���&��->"|����-T����5�bw�5U7-�;���E�.���$7[9g+�ᷙ��"���O�;���9%*20W�l���~�!��C��
lr�nj�+P$C,��5�(�y�k{�6�<�<�w2,������D��2�%
y�W�L*?��]�b� ��7�܃��x�]�?F��t��r{��QV�{V��{p����"a
�$A�7!��̘h���J��|�6r�g�����3D��u�M�ʙƃJf�X�ZqM����p,{�Xs�%�I�a���n�!�sѵ̍���y�(�l�<�I�Ma���w�l��f�V�F� d`F�S��A�Հ!�8��,@E5s�0v��x(��;�j���yJ&�N���|�_�;;ۄj�8N.�D��.5Q)[o��X�$�o��V�����E��d�rc���_��5sH�c�|(����m��c{�jP|�D��FْΠ?���T6%#���c�����45�����Zq�`�˻�4�� �<9��ܢ�<��F���tQ�J�*ŵ~�~�x�u�L�9�o:��hg�S�&C����ʓ�/�|�A��� fA��蒨�6]>j���n�j$�C�����>��g��*!vM#o;h��Up�y�h�%;t�q��6��fdc�
sQ�	k�iattQ��EEB"Rd�Y�����~?�;X��|�O�6��-��*X@�]�o� �IWE*�a.�P��o1 �ؤ��^W����`���N��A��;݈Q��_+�ɽ����ޢX�gyc�\$�e^�C���`��Ч�T�:�%���My�Х��^s�N����b���|�3�ʰ���q*�<����x��:�������wz���
pgP~�.����2���V�*=�����F�W�r��Wʔ@�6[�ک���]
�>WC�W�j�m3	����N���#�G8
�-��Z:�P�K�v�L�tqS!9�U����&S���]+�2!<���Q|�͎	{����J�¹iR��T1*OO�iT�^wm�G��!�b�;؞����귽�aI�/xtPÛ3�o�F��?���7~�d�:ލ`'�`e_;
]p	[D]��	��	E4�Q�m�]f�L^u����ZH��4Y�k��w�@j;�wZ[fЈ�&X�a*=aS#�V��r��Yj�m��/xl����k�*�S2}��>Ȯz��ر�,l��q��eL��W�t���.8f�qJ8�.�`��>Q�����I\�j��q��n������>����n��.��ٍ/��pkL5���T�C�V����RÁ��u�:f�_���!3@�[�e_1��=�h���{�ݢ!�rDn��(y.�� b}���Y���H��6�'v����&��� ~*>�a[8_46�K��M��o�{݋2F��މ?�B3�.*z�m�:�?
�dvm�Il�8[g����S�u��b��S�W[Y�=&�ov����~X��f���a↼K��ѢPl��	���s�3�6�5������F�g7f���Fz>�EW�(ޚW�?=X$?��~rh��\�����-�؁qu���W�,���ٲ�T���']��{�(�m���y�]��)S�����A�Ý{��tK���D�8�/K�s��U5k,#�~��f�`1cO��u	&���jN��⇝7sLI6���^po���/��8�D����zu-�<��iʏ�T�iy(-6�Mo�Ͷ�2P��b�ݼ�{T{�m�PR��PĽXvhe�.�vtF��l��2{ՓEgP��W�𜿍ɐ�skN���,8z�*/��¶خ�I(ؼ\��E��A��(kb��U���h+�I���n*�^ZK�-��dǆ�sKO.���a&%V3t�S	��ۻ�!��-\����r��D8Š#!�x�,���:�Gd�"�_�� �k�"2I�  �� �u��f���q)��
�A�Lp���o�"튠�`�('.��ϐֻ��S%ޫ|�B~�MkT[�?������;��������V�� C����w4��XA�k|#]������S�_���,��E�� �q��~%	�P�S����s�� w�v�q	�W@=1����Xq��\
��p�Z�vP�b�:�a��ĕ�#���F��\�P}��q�~�t��m�Y���U_���)�k���G��EU<1/.���Ĕ��	�N!Za�Y�@�2B**������m�=��q7�h�qf���R� ��WEm �m���&V��Sj}�]�e��M+����moڶ�i���#� ��+�]B�58� dF+3 �W$H�d��hWG��p��ލ�V��d�M��DY0�\�M2_/��%��g�!˳�q~������s^'��&�\�ww�R_`�߮�����s:�W{0����6#z~����q�|/1x�	 �����O��I4�QફO��Z��~�~@����^HB>*'��e}Đ@L���%Eb��B�����q�4����Űn�9��pT����4�g��
f���]��I[n'�܊��̃D4c�B�0�ge��У	���:�O��%���ڲ��G�=w����t/����5S
b�څ�� �`;�����',���5���i�\g�����h�w�ý��G���^�X��c�G1Lj	v �k�����f ���7L�M\���0TQ@x&���k�ϙ��WK�J'_�mX�V(����ϟ��@��J���u)��Gf����|:LϘj��"�m�[�lg]q��㻟Q�I��&&��k�o8zq\��Fxq���k?�si���r]Fbf�U坯�p��{�o�*�*&� 6GC�m]Vk�B��������K�,KXf%).1��?i����K���c�f���b@��<�i'�e�܋G��:�_�jR�����O��e[���-��%q��1��5��ܸv�������z���E���E荔ӑ�2&�H�|�����Z�a��rn��t���#��KC�����.FQ�[�2�IR�n�v�Dk��	 `�i���y�5�S��7�lըa�g^�]�`��^x�)naDt�V')������n�O�R|MV��+�)C>�����f�j�"��e�Nȫw9�KP���*��k�#ɱd��&þ��u��l�J<)>n�!8�vf�2A�S�c��OR~^M��(w������g�H�3���1�y����"�&nD�#�j�F(�6��凷�{�XY����3�Q��=I��;e����W�A}�DIM���K�9(ET�#���P�����R�I���>������.Vn^%S��V�T�r�Z�/(�����$Y���a�CeR�*İW�a-�zսW����{&��m���V�Vq�	Њ������;A*�WC�«V�`!��5���/>��\m�*�+D�%i�:�N���>�$�s���
��#��)B��Ρ��i�4����m�h��8�7O�ɬ�ӭ�=ȻY� �_Y� ��6.S�1G���U5�^��$gF�����4v��?2$ieŏi��4.���k�_�oG���~��yMZj�6�:PY�꘥=�����{���t*3`�7����W�j\g�?����Ss͑�Ή��u�G��qC�c��h���q\"�9�%}���CO
���^��X��5�E$}'х�z�[�/������m�m3�ǵV!�ǘH�Jz�;/Dɶ��t/x h�������˘ ���)7�O��LĎeD����������|�w'4���ʚB���M*J4:�=�~I�|�t���gP�:�&���ub2�ͺҾ�[c��J��o�!K+�"��W�Y� ��X����P�9u���.40O��錡;P����ۡ����խ�9����U%���М�r0L�_8���.>R9�d��O}�{��Q��Lb����|s�l*���q/{6��L�][�����D-&Q��0wu���-�y/VuQ%���AA��4h�"�����p�����0�dp_,���8|vH[R�BJ�Hy���9P�ӕ����M梷�έ�X��]��L�伧�2�Ȼ��j�(&��R��W���\=`B��z�9�mb��.J۳� w��i�ҝD�0��;ߺ���b)s���S�%ݻ��[.}D1�
�V�BI�¹����}�+�񎪋'�>̲i�Xv���n��a*��
���Ô�pF�l��߅���g��Z�(|M���38���M�VG������D��>4 ����B�ܰ�T�>I�:ÝR�n���}�?���[�)��|t����>���X���HE㟶���s�m�2*�+��6��߻�x�:���k�r(�>dch��O�^q�=��5�~��������@��{i1E8P�|����t���QETF�%����%_��}4��?���#Cl')�2d�w�a�F&�@y���Ɨ��Ï6������I�wBR�&�jG�뉜��� '�m�g�#|�31.�Q�9��
O�2iy��+�|�����b�7Gm�0�狩�~ؤO�r6�}�-�<��+�����ܽ�y:>��+�7��fj��	���B3����`��7Ym I��LUo�+��~V����U�	�*r��f^���U%d삏��f�$��z����bX�8Z�b	#�m�EM�a��|=�����<(č}fR�����^A���##�K9���%Uv��M4���=V���c�J7	��9��vXV2����t.%��n�f�Y�y�-�HV�N�����#�v�S�n�=G������TN��L���Z��墄��NI�8�MA3�~#�wc�f8ɂ���<�ǭ���#�,{d�0���Sh��7q�ch�m�Sf������l=?����(2��ݷ�d,=�s����̣�2]�J�8���p
����sX���a�E�4���t��E �g��xTi%/���%t���K�c�}(K�˔�c�d����c��CCJ���4�S�rQ�(��Np�D=e�ڲy�] ��N���\����jC"*�tv��>���JD�8�����	ߜ����E{`�F�+�q���޺3���~=��;t+�5������i9�U򭘘j�K[}έ��ݘm{��,9�:�{�xX�V�65����KԵ4n �m��ʟ
fxQ!|�|qpV���	Չ�@�U�c��ł��}��1�&���n���ɦ�����j�4�7ڝQP�(��ΒtmkS=L8
P�h��k|ƹֆ�"`��tp/"K��>S���������k���7I�p���gl�9T��g�A���[��x�aj���|#�������<���Ζ؄v�����"���%B����c�:�	׌Rk}ȅ�LԊS���?%�v�(�w�'\�!�#�/Oh %\ƖB�X)�h��-oZ9���\p
5-�u�h�("_���)E����)ϺruA=;���;�O̛�悧�� ��*(H2	p1咡�7-�.Y���bTFp�Q��,��w;`ǜ�p`�� p^ �s�7"h�Z�%��
i�@K62���2��!y�m�������r$e]:[-�D3�1�&@��٩@CD�X7^u�1j��xKͥ���`�?�/I�U��&���ݘ�x}�y_�<U��jߦr�`��d.��Wd�������C6^��� ����Z-�N��f���G���l=de�f4!P�`��I3�y}sg�:������)*ډ����}%��5�؊����5�u�K0�&��Iq�ɋ}��4�J!�3P��Mg?��\/�S�)M]�n~�TU(V��r � ���!s}��,]W�ɦ^�F���x2�>RD،B�y?i��S=�_���F_w
��z ��}�؃^��t
�3����&�g.��L�b]� ib�
+����)6o]x �&�c�&�ܰ�SN y��^O'f<~,V�5�yQ�	�uN��c~�V���
pJq��|��d#U��ޕ�A>�k���v?���F'@�����z��`�i^��S��5���'W9)~�D�t�wR	�OcZ�:��#�8��}PV7�#&P���q6��m��TaZ�*��H HX�`A�����.r�Z�⠯���h�C��S��>Gb"�*��_��*W������?�ҡW/�xMCTb�ԯ3@@wLss�2�S3;͞%��s͎���`��>�3˜$��`nN-���8���V4�O�}�t�~Tv\�S�E�e!5Y��i�G=i	_�����:���P�l|��2mL��..��[g4Ρ��J�p0X���L��ge�ie8�sJzH5d&^����äY�aD��w[v�7i ��|ϩ"�?�a�YO�_?��c�j9�/h=�ֶ�d��}E��F2�R�36��Q+ⶺ)��A����+�"X�Z��U���qO���[
�E'|梻���X�j�ɩ�E)��V6S9#�%�������E����)�(�$���p �a�^�pjM��[ׯ��u�ɨ���/G�	@�`���Kt��M�#O%_�k�M�v�C��C�S�����|7%�rO�`� �8��'�8�,��q�]�Ӑ�0R���x?08TN@��cWCx�x�#c�EV����\�&����.� t�ˮQ*7�P���194�T#A�L�lo_��r����z�1��L�3��l]���^���5���6IF�E:S�`��2�d#��'��d����@r�Q���&�*Ȓ_@|�!{M��3" 
���r�![�"��CNG����g����Ĭ�ge�Tx1@�c�JS;Ĺ�'Gv��z"��Jɿ~�`�� <�)��A�K�;����6ʒo�\P�;�0���Y�'���d�Ȏ{�p��?o���#��h�Z��~m���o+��s_���[ұ��[)��Wy�]x�>|de�<��9�1��B+$A�4S��@NnQq��\�YJ�
+��R4bZ��de��k9��%T]J�U�nzڈ L8������1���N8�#��h���������qX�2B;XՇ���{��j�K}\�Daγ�ES�)~H��v3�k�V{+p��uPt���Xu�E��YA���΋f��pz�tU��_��i�������w��|T��a>:��-/}C��,'�Ѧf� �s�?uV���Q2�۪��6x�C�2�?#�16X@64��Nf�������Ø� S7���zoy��sm�ݺn
��ՠ���$|��z5@z�H��*l�<�,����'���҈��	����`�Zu-��7P���*�I�^5��Z���M�P,Ŋ��/a`�F*/e-\�Jc��T�,�цmi���_�6��dj~!_�f�,T�7�b��e��?�aҵ,+H2O�l�?}5bA��Py����,ر�ip駻i��R'm��c�6W��`�e;|�Q�V�m�U�3 �k����EH9��y?vZ����1>�ic���k���n_�[�P���^�b9$���	^P�9w��B��ⲵ8��R)gi�yc���i@ԍ�LP4�s�>ܕ�b{�W���r{o��0���NwrK3�(t d6����	I�Á�^�����94�ȑ&ʂ���`�[�N�jyEzh"��N5�l�����Ll�~;ЄU��7�Y񜿧�E�(�0���Z
�����UP9b ���K��}}c?-�Hx][��w��/2���ZVa��6����V�n^��&�31=C����c��3����q�u�Á�g�B��k�)l�N'c�Y���}���G�]��=8C����H�%׍�>�|���^����6o���Rt�� �g���<A�J��N1kI�2���?�4�ˑG���xʿ�yXݗ�E��3�_j�b��_�w�s@�����_kG���lf
���JKS"���R|K��~L��(<}����2N�r	q���6^�*���I�^��l��K���d�Dd� 	[!�T�JP&Qq�&k�#�@d�	A4�i�@MWQh� ��9��#M�]��:���b�2a���&��%6r"�2�$k��nAr�JB���<�n�zM�-J�ĥ� �����Q&�t:��0�W���C=~��Z
��8��6���%���%���`��v���_6J%�N�����JL+�7{�a C�#��j�W����/J�H	�g�`m[�83���\T��;�,w`���;��
Ǎ�H� "�� j69m��i2O���;禑��iO��w��=�]����<N>9�3�����x���2�f�ɽf��o;ͺ�.����!��J�=���7G+ֿ�:3Q�G�VP'�I�${|�X�t}��Ӟ
;/���q����*�f�N���U�~��.�G��8����Ł
�<3C�і� ����˄���}� ��L��PQ�8��LJ���*�=��|AN}��	.6D=���)�/�](n�i,w����zZ��t&-�eD)�������.�������>����5(�|>Z#-2����)�]��� ���#�6�7cR1e�[�Ӕ��|?M� ֋�ˀd���(�/�]�Rd`�%c6I+���z�E�� :�dը(�����M�������\��[����TTgVl����.u��x��������}<���,��4Ro�R��(�U����a�x�'gƝB��i�~Xɇ�,(D���s-N���[%��:�cn(N;x}��{������k�rO�rkm�+E����`�Wn��� 瀡�;0��pu���ɮO�0{����g/��Iչ���\�qdgyPG�ҩaWE�"�A���y{@�<�VTh���Q��z �T�Y��7>R'ڝ�Ȣ"J�{�D��H�Q��%s��zp\!�A�=%�ѷ�\$Qc���1 =
LQap>TǗ�J�H���d}[P�KNK�h��%���<������P]v�]�!	�dd|��_��&�#���:מ��5�*�Sa�d���yy�ɠ�%�*����}�3Й,�V�h�ŽK.���|%����������M� ��4s�'���cmMeN0Q�C�=�@M�v�~�U����{hL))�
�/�ofg�=&��E��q�� �;�N���V��g���o��h���B̕X�N����}���Z����b���h8�*���D�������"�q'���p��}$|��?�qh&��נ4�r��>}|3�SJiT&D	��J�C>��X�3 ��ɂtV%�V@C"���,�*��ޣ�����q�3ka��\1��z��|�ێ�jr�aQ�A���	�`<��wX�e�bc|���R�b�r�O��Kv�ٷ@��Å��k��B�3v^KU1SS�	U5D���#�X�8�<��i��~����h��겷A
�Cy���F��W� X>�����	�F0nT��<������A��Ίx�(o#������ju�j2I����Je0���	/N� �/}K�����W0t"�%�
�X#{~O~ml�|l �+=!�7q�B��./�w��K�N%�'�d��cj	!_�'�k L���e&w��D���n��>����&��o��e�(R���w�u���~Iu�;�o�\L	Uyo7jLxĤ��-���4}$��T�0$��A>ZBT)��`�An)s����&����}N-��9��;��6h�e�.��֮�ChhJ�I��>膶��JI��>̫XN>jT��j��B@�ka��k2��rA:�v&$�;�Wb+���{�wC�D�����Qv�O�k���M�E�-�E����-F"��##1��q�sYK$]���;���|��3�B5n~V���o0�gH��8���Pj�<;_�³�F	��N�:�����C�=��y!��d�
	3��p��O^Q;��x}��U�)���}#|��Cb�.��8B�~��z��s��Q�v�<�Abq\CX?����"�Mȅ�|!����&؁H�U�0�9�WА;�~6��
qP�
�zgqu(��7	7��jD�!P����=;q�H�a,��S��#c�=)3��i��P��ݙ���\����`�d���`���|�T�쵆�^�T\�GX�-*��T��b%N�r����B�� Q]0	� ��/����0^�̀]�}l`F����oxS�_P��Jt@zsOW��� ?v�g�~��/t�(讚�xĆ�m��`[V(��M����T� T�@+�;Пq���|CA��VU���ܮ���g���Q��6޳�JUDr����R�4��D���6;?��jbsn�aC��*�f�/��^`�{봍w��'�Dv߆
��6��s�<�_b���׷=�i�Db���=�c�8�\Fͧ0`�}��a���h�����P�]s)��d�C��f��{�y^�����B�b�4�K���=-�q5�"#�lQ�M�{�P�O!M[��]T|��\8#�.��>$6�Ti|��]��~�Qӝ��Ξ�grx:s�<������`��L����(d�?�V�����mm�d�����?�qv��@�s����M�ǵ����'=�I�(���_~�e���E�����|���V�&�9��zo��&3N��x4n�c�5���]�Oh/�����s-i�?� m��g]Q��J?���oȈ<:Ư�^�1�1h
��u�z�V�ù�K�����������?�񱦮�4���e�����P��&fɸ���3�Mb�
M�Q�D�^mM����]��ՆW�1�L�G�^���YݒjH$=�t�o���>q��\ GG���B@��9��@�fP���������l����6�f�褈:+������K�k>�؛��P�ʗ���!�i3����B(���ǧ|6�D<��5�D�TFV�o9�ëB��%�&�?���'��Kw�w,Z³���6Ho�_�'?Vlų����5��'�����X����o}5J���F3��&ezDVmI���i<fNc����F�#�L+H����r����g�AT���?suG*ßO�j�΄zz�gi-9�ƊOs��B�M��k,��Κ��'�P~�.8(�r�Ug���9���KIN�S���3�7����j�&*��I	 T6Ȃ�M�3��PI
�x��]�i �A�� 1��r�;�9�2��a�O`�G-�+��:M���ߧu�����<-��(?.R^�����[R�<�'�xd�T{�3� �)5����1�@���~{�^LX��/һ&6�����<j�	��5l!I�qe�6Y�i\�%/W�z�y�pz|h���Ϩ@QX���0r�+���,;ø��p����.�e�$(�J�qfd]FC���ʻv$B����pP���k��fm���m��,��L݃�KR�U�U�yj�<���x:NmXV�]׿{r��_˴��y�n���3_)O��w|L١� t�,�Av��F�j��s/�� *��҅7��y� �Ϯv3��c�7�H��Et��+��]eHd[����m=��TXҝ�y�l�}���)�$�a\`�Y��Pe�o^�"�
p�����T:r�:��7m�f��=E�� rd�f3!��[!+�h�:���lVx��l(�7�r~�����gh �� ���Z���"�'W`�tֱPL�̻�`�h>Y?S!\����#D+LE�Џ��F�i�����+����j���+0.=��"F	H�dHy�D�I�g���6��&ݎ�|���/�x� y��_r���$OK���g
���x���S���z�R{s�H)Q�Y�
 N'�&�P�A���^�I�S��pO�Q�\�)jQ�,b���W^
��) ��fq8&�L;�����%C������mVpl�� z�*Y���u��lφ)'�sq�0~����5Ӳ����H�l��t���(,�~H�=!�Hrȫ�-�]ՠ�O�Ά�?�T?��'bs �G��I!�.�2VZ�OƉ{��oM|�W�0��Wr��R��:V=��n��4]3�p�$D2����	.$|�|��8�?���~�I�s��ȃ��*��׭O6�u	� j�X��#���z���rЛݝU^ς�B�d頎��-�[�����d�\�C�!q�V��/{��ظ�]�/�)"~+���$O)�_�}d������E����x��?��������M���Gc��ӰqDUP�|�q�{�1���Ӥ7s}'� 1>�b�5eV��G�)ժx���݌}_@&����<{[�8pn"�`ijs|�H 
��:(�k�'��iǓ�@'��<���=�ʉp�^��}��E�����z����	I�`f`�L3���{�CL�����#�=3F�[����%�����tY*��>��A�{��}Nc���JEKo�Rg�%.68ͥ�x&��O�|�"�-˘�׭8�̛�@R�i$��[�gzt�МmgX�t�0o.��ߚo�ⲡ�-��ݣ+�gh��yö#����
�d��H0:T�x9�%��!��R xW{��m�m�ה`�שǌ��7�<�=�׬���譐t���t�r{���>���28TADH��%�M⋈�B�h�y�^n+�$�p��ݝ�� �t�_���)�7���_��Ռ�0x֦zC�6��2U�ס�D*��áD�D)�����
	�;�e\I.ntS��O^!�0~I�z=����'j2�9��5�zB��k
��j�1�
zJ��|ߐ,���X'�i��uA�����JY��
�����l�aed<�_��h��SխֵPD �@W\� U������^�USN�[�c	�e��#���{]N4'H�7���\h*�Za��x��Ӝ�o�ᰯe�j�+� ����%���:O�CL� �ƹr���GB�����i�`y],&���$=�nm�� Θ�B���E8.�aW���_�4�5W��a,J9��î���í�͡0?HP�Fإ�%Ȝ�Ҙk D�qE�6��������EO���7	c{h_�,9g����g�T����St}Y�j�N����*�Z���6sB*��w�SQYt�C	Hn��0�%�4:8�Z�
Bݖ�7��ŗ�������G�N��җ�{�^�1����L<�cMTE���=���n�>:�O�~. �F���S-���umf����$�UT��H�qnv�ٙ~	�.�UN
�f���'��k��6�&2�k�?��(P�y�gU8�`H驄n��X-�����؄��K�O\ku�L
h:X���EC�gS���WP�0⡿e��Od%���+LQr�$��%GeV�EQ�?/�wz��ؑ�q���"�0u��d<̉'��X3���LhL�U�k(��%yk�R1⤮�D���X����`N���#�^��J�e
��'��}�;�I�����\�~�TnyF��AK�;N}K-
���n��q!]�%i�C��� P�d�/����X��.�k�H��x�[�:�}L�	�W=�&�ɔJ�^MDuU�����ޖY�Y4^b��u4���� ��/N�|wx����G�n�hڀ��x풵Q���S�D��V�l2�D�GNE\ә�\5�ӝ3kr�k�:y�Ҭ"ŁݧV	����T�a z-�۹|Y��W-g�XJn��1+ʇc��yj�'t����d�~W`���}�����g��$��U|�d6t�w�.?���ݮ�N�y�#ϼS����8��|��N�\��p�fDm��,��8v��R�D<�f�"h�kt����<![#��WW�+؄4�Gp4����9�V���7Q��:��IC_�)gͶPr-J ڂ�����e�ޣ��-s���(�>�c�8N@���P7	 �'� '�o����7�y��^������M�Z1Ia���l��L����L.,��0��bʐҗW�!��}"��~,�������L_~WM��8	��/��|%W9��Z����}��7 ���� �#�^�lmszS1��X��sS{BL�J�H߲܆���Ȱ���i�3��KM�C2CV�+f�뻳'4݊�f�PK8t�H�ݳ��N����nj,�@$?O6����y\�gZ�Qќt醢��i�)A�h�Nj�B���ʸq_��;����`�Sm�'�1�.�h_�Is���{E_�)Oʱ�')�k/�U%��ǂL�TL(ꇘm$�l���&�k�s������f옸�$���.@�@�,�p>C���ԙ$c
WY>�*x"�׹B�F�~��Ɍ���&4��\��$~�x�df�m}!��0z�ؘ���$0�溳#DϛN�Y��F���l�)I�)����J��R��>��7�Xe��b��f��u@�;#��.����d�����i��K=�?�pG������Wޠ� ^�O�0�Wu;�TNgώ�#�I(����g���W�Κ�)�{8���1��1(۩��l��uE������M�L���'�Eh��5��G�G��2�nu&'�Vk���)]�-�2�8��+U�p74y:
W9ѿ~�L�C&d�0i�0R�ԑ>)�/&T}ř��y��v�k�)������#t.���w�_<�_�:�"H��ʰU1`G&`v9��7A��&vo2ό�/b��/��V[����`Ľ��Ʌ�7g�UC���ͦD�7Ԁ�(�5��C���C9�u�/�IA]��<���x���Xu>&�I+��^R��%5�3�M��5��(�B�������,NZ�^2�LSg�̧���,��C�W�����(�嘎�(�~?k�I46S���l#%��4�l�Aۧ>�z�2��l�8��F6�����N�Pw"za�!���26���Il�Qu�^X��udS<jt${Ѯ@9�E�������E�u���2���x3�
9�L�@�K=����k_A�\�Htj�����p~�yAyъ�!;��07m��f�L�G�+@S&K���u_	��_�/'T!��xSbˁ$M-��#6mT�Q��͉S�3,=�'���A�5l�������vR[�c�Iҧ��we�0�#�{|�����	����(y�n��z
[����M��qK�Ni��}q�#��[ӓ_\��bT��3��	���A��L-��������<�B��n%�Eu@��;ݒ�)�G �8�cO��4[�k���۾a�~�\�.�QTԛgbu��'g]�패����q�Ώ�vN����0$ᶐ���#dh+G����6|s��BT-��ף�ٟ�m�G���W7�O���pO
zX��-{=�j���QTw}�@���d_����j�H�H��+�0b)ANS��!�O	����\l����i��f ,��Id��B[u�2<���&J=�\Ÿ���$��)��v����{H��4m�h�v�:VvĄM,֏�.p6����ğ#��۞�+�����b[�]#U�eI�mc�����
��?E���j��'�oM� mON���6KIQ���փ��FV�����b<��M���]��A���2��N�l��jc��oFj�&�h-.��]"9	"3�
�'�Q�\�>��˺�1��`�-�"{���JX�9��3꺞�-tF� ����$����G��Z*^��Oh�B"�n*f���v���Z/楅u�/v���%��l&ı�	T@��!f7���E��
�j�Cr��":�헴������_����E�0"���
4��N�f��p�D�Lb�U�`]�]%�@��[&s��an*n,f���%��۰�6.0��� �@R}e=N) ��h��TW�V�ob��ٜ�iҢ���91��v�?�	�h�`�M�Y`,n{���{Qv��R��I"�/	�!j�|Ē_�䮀_�Lm��[@<N��<�`���	� X��0>�{�IՕM��X�����)�V͇b~��V!�#�n]�/F!n�9�O�����q�1S��Q�	H;\�V�kE���,j_��Ϡr
ǏH8}�R�8�p���--�aZ^m0�Iy�.�aZ!�+B�E���[�v�ّ���Q�Pf����hk׿���yє$��A;�S�IlPmSN�cH0+���e��X�d�����x�/'�r���+���x�۞q�K��*L"��v
���O�yA�r=�۰��ɮ!�^�sѼDǓ�pS�j��p���}�<=���j
n'7Y���ОF��.� F=@�K���~í����h�� #�"7�M^�o<M���ֱ�֞Q?���ڍ�i��$��։��B�"����a 8�o���k��k(>�`��1��$@u�MG�vL;t�hfw:��M���?|.D��}�U���	��Ep;o1�֎7�GW�M��Qt��x�T���	��+4)��J�����>�н݅�����T5ؚ�,�~\_4�g��s��"l}2l=��F D9V&QXǣ�#5�b��Z{���k��4.��:�u��JA���{�+@� �#��?~a� p/?�e�؇�r���ͫȩ��=��if-S�!s�:����߭ �F�8��G�oQ�j��TTJ��l��<�Y%_�T0;� ߿;��E�6
+��2jpU�!�Ci>h{��AZ(c��� ͍�tY��J8�mcHپ����[��q��=��+�|��/�k=�='Ħq7�^����"F3G�\�I�+�֫X�|�ઝ�+�d,H�B�%��0˹�`p�e6a�o:쟱��_���� ��3ƽ���z�d��&8���^Qz���~��8Ɋ�t�ͨ�`� ��2�9��R��$$3c�ɿZb�~*��W�.��,��vM������V��� Jj6��	U�N��7�K���n)<۸���3�XZ���x��9��'6� �E�k(s��ٚ���b����˵x�IVo�`�lJ`����y38KV�I��$�Bזu+��X�N� H��೔>8��m��	<�'�BN�Oj� �nE�fH��EԵ'�
]�A���ڞD��>a!�K��\��(,qD1g�tn['�5��ǩ�t�x�~�jC�5��냀3b� ��td���}뎕��k<�[C�B�<�~釱��U�?��H���N��Ģ�_# ��o�%�M�һ�~��'7ez'��]C#_PG��#ޥ���<~���Y��w����z��$q��ڱ�T6�p�C��"���,�o%kѲ���j�@1�w�d�è��mp@�,)��9Dr��5C�rS:����rH�l���He�����!�D�z|�I��]�L+�
�h ��Ηp1���6��=�O�v����)������|��n���
��/��LX���g���)ȓ���D7�\>H_DG��f�1��&{�6-��s��'Z�Ѝ.��uJ?�,B3�T�(������Fu�=��Q�F�rf����%YV�5�]�$.����}���5�"��P���G~/��y/���c�pR�s$;5����.���;w��`&x3�G�����+ϱ����rm��x�l9t�Ɍ?� ��3`�#K�04B�;���!K�w~��8��/���XsޯЎ����+��_��:��c���+��*�����J6��\$)~�84_��Tt��㠱���Zܻ�����6+���	M^U�ф�>Bp�,���p���+��.�'���1Y����&I�g|�u�=���qJ4��OR9(:]�Rnkd�l5,8�}P��#�u��c��+�Ks
=C����eFq!��sW[�"�!�0��@bˋ�.�eI�֐��j�i|��yXGϷfUww�"w��c���{��Twp����:�"�l��0I�TW,cxHz���5*J=��r�
����8�������KХ����q5�Fм*5q��w�X��m��z&�(R���87s5��B�henv��L�~�����#{n��rY�?i	�z.IN����@��:���z?3��ͧ��9$� sR2d��f�i`����MEE����H���?��2/A�[�����GF޷�jJ
Q��]Ep�/��7�x/�R��U�2Ӳ��rHL(ٸh��w�3Q�^rG�Z�Q7�F-��ޕSʯ.�y~S���<�|� �TWY��^�JjR8\��T�=���;!��ѽ�j��u�G��m"�~�iⰶ��Z��ؽ�۸!w�~ԗ�#�w�m�v5N��y������>�GS��Ia���<2B� �٢v�8/�if'��UN�π��hu��͌�(�O�?3��2=dS��G&����`��<%۹�1t&7sK˖�����\x^�5�����)&�'L~��k�O�&��WW��IZl�A��ڈ��Ζ�!���C�8�.w"f�*��,X}� xF�[�䛈�Κ�;Nəx8n�B"��/G��֐��L����ͤ}�W����V.?��˴[[�����&��ӧ� ��(���72��+�h���ur�E�PB� \>�x�	ػ6�ej~煌��
q���v�/�Wi�
n�����)�g�PKԖE|�(��"�e>eV�lO�\��EYkh7ŻO8�3��N��+���U����=jD��9#�WEU�6yFL&L}��h�Z��`0�9-����Fs��O#n�v���B���%\%�(�z���j[�Pl����c<z8U{akA`�����-��,P��Y\o��I��'1�u���[�
�E�2;Nm;�3�L��Gl(@ �4��t"�7�8��r_v9֢YCB�y[���)¢��-��\������B;�"�!x�v�W�.U_p^5�LG:]r-A�A�y�;J�x�>pUcY�� �1K�)�a�o�o����� �0���l�T)�]�?ՠBI��sEǍ���T�q[ИP�̳�YQ7�'�- b-�m�cx�
U��C9-O��D�WV�V���Bu4M�"����r7�B�T�O�p+�@�r ��f+�.����H����y���|�yū��<�G��(��ؒ^��rS-f�g��r�t���S6K7��:��IF}D��8='�)8w������"��F������@d���"Zr$��T1�lkMm���J����K�3<���ǡx<^�RP��M[蠘k�+��0'�P�g'ȼ53���1n�e����F�� {����g��'��AG��,�m�n�	��u���ǭ򓶫��v�AE_ߕf^VI_�.P!!�;�t�����+P���p�NAZ YA�_�,�vÛ.'khd���ll�E���csN�J�#Q2���LG���s�Nd۬��TL�^!��Ŋ����v���EyA�L1�������]��K2�M�:l�Y�ֱ���x ����.[!VLvBl�MM�S�)�O)l�b<�<��{�r�̆�9]uy�Fr�𔲳ov/�A-1�@�/z��D��G���wK��~������A4^�'+��[l3��6�cBҚU���-[ҕp}	\��$�ם����_� 	���jK�aR�*/�g�m��B��,���C��������2��d� ß�%��?�l�?�����8ﶷ�B�X�h��:�l����Qv���iθr��M���C����Z9�E9��y(0�b��*�{X��_;�h>��]�j�3��r��
]u��x�l&1�ɐ瓮�ș���ڵO0��y�<h�����ꃋ�{�����Ms��QS����dབc���-�1�ZX&藁�Ǡ܌���jr&�^n##/c���{��!��W�_$CC�u噜/��#&��)S:\�ֆ�����P�Z�Cl�]!]��jO R�����{��e���d���H�!z⣿<�&Gi=գip�a�d�>t�z��/�%孆��D���#/�������������]=�G���8<k۽Z0(�����4ۮL<����7'��u�|t���t}�s�'��s�h8O��k����Y��FM�#>�϶���rJ��U(M���]���C��Q���.�����=X*ќ`�ޞàr��CH.�Zk��f&�`=gE�a;��&=F���g��~`C��C &|�20n�X����R}"���_��'ay���s#��B!�I��+W!�EI& x���:�U<�[ILD�8:�qle-�_��#�z-�N�Mh��=��LUY�����f�EW�e�}����������=���_��潹�ݢq�ܡ?�O�H�A'�S�Us�jP%[t�����H�x0���z��"@��]��㵺}q��j���|5L�I�����⦇�L��k�Ж�C.$;Iafv=�\1�rWO���	��9Y��5?` �!G�Uu��-�y-�,xI��B{���h'��\�(2a� ���Q���ύ�)�h�����J�b@sj>�Ү|ne7ֱy�ID~����g̓.)І
��~��t�<ǣ�I����3�%+?�B���
�����'����'ӓ��i8���b1�]P	}�兎��ܒ�q{�2ː�4�Et��<!"�������oR~i}SC���O*Va��o�1�`��|����[d�_AP �TNzܽP��҄r<��6:�wt�O�w����(�,8��V�앨��i���Q�xE?�Hg5˥�� .G���${���h�!�p�����NB�{�����>�V�ZM����D$��d�襞}��j"�?T��22��dsZ)ذvJN�����^�֨���x��?�&��֯!G�ǳ��u0�B��F��$�?�{�4C��p�#=WW����d;O[у\
��\��W_Q��Nՙ��1�hJ �:F[�vW�/�&�u{b-bi/��}�����Z��*ba3�{oF��)������T{ӈ=#;�x��`��ƜP�t��s�
38�[�%��RJ&��� ����'�
���.��Tic��Z���LXgˤ\�EYᷱp���r���	Y�ȿ���Lv�v!l����@6�.�,*�؆��@Hn+X�^�C[��朚��C���� �[�%<�A��ĵ}-��>�"l�2�R������
��jU�do3G���h���ߚ���|u�4I[k"���	:��GW@:āpp$�x�{���5���&5���� uQ��u����ϡ�Ю#R���=,MHu��X
��r��h��?�m����� U�-|��	idҌe�ˊC��k������?�R��1���� ��y���7x�wVe�L�g�j�G<�^&ӹ�<[��_cp&������2�JIae��:�C奤���s2���<wn���l{HG����^�/f���6����{3��ؽ
��|0�m\ճP�н���-��G��7�L�iP������#�
]]��L` �*A��л*XVP'q��gÑt���n��fE��jK
�bd��nǝ�l�v��Q��h�9�����I�4�^7�C6s��9�HF?�<8+B?��;4Ne��:x�K%S��3��_\G@�.Ļ:�÷��='�/_?%���M2l��ޗ*8���F�H��u���[����:����06Lr1���Y�@D�(�:=1��D׽t1c\�q,�9��t��| V����o*N/�0뒦�iɣ"�DP�)(M�� m�/��\*;�S��UP'c��pŀ���얌��f�a4���Uu9�CQ�
��c�� js1��1�(��
u�[��xc=�y�ȧ����F�p�5�kj 2���LK-��0"]NDWPƺB�hP�|�99�R�������r{]#��b���ْO�&�"�g�M+P:sEҷ��g듻�L*fM֐��AH���-9B|�֍ճow{�U��s����Û�	�)�F?�z�B�_��P��xcˌ��؝�@������eMbb�bgP�	���s��Y�V���|(���W����*d�`$�����Լ�p�Һ� �56n�Q���4� `��p&��%S�!3��!���p�r:�N�s�m �)�0:07.�E��7��ĝ��Tx�qǆ�B�'�x����li�b���X �S���{� b:=#�`\�?�b3����9��˹:	K��V����*a	μ��o�QT1�W\~7��e��Ԁ-�gu���aJ?� �S0��B�_�F�}�w �qu_�"�$ g�J��j.*qۓ�IR�������Ѓ��
�x�c��6}H���y������n�pt֑O�f-�����D���(SmBt;��[�����ڽg�(�h�F �eN�l�� �a��Պr�ܺ��12����8��S��f�S�S�c��2}���\�$X_[k
�*�e�g�Щ#����FBd��ҙ��q`�ک�.I��`dB9�Jt�L����3f	��f��Mi�ƺ���!�W�.m���¨��S�ިغ�Qk�<}�J��D�� c�䲋|����RHUϙL�.=�ԏ�����1�~�d9�x�$d���_�� �\�:+�3֘��5��篏���-��5 v�f pD��)Y��7Q��o��
qm
1&�7�!���JA��P ��r2���7�����l�Ua��%D�p��4����`Uӿ�|Нb_�/��i����O/2�JzsA�]�@��)-(fu��d�P��d�2]��Hc���ox������Q:�4M'����ҷ_�cz�%("Y��Ƹ��uXY�s��Z�y�c�%��{_%��yᒒě-�h&/^o��� �ݪ .�+ӡ�D�շ!��E\���n[��g<����=ZHp�O�%`�\l��su�uK֝sk�w]����aOK���]�/��urG$���ч.�w����x質[���%��C���c�/q$d�~�]����D�pG����/��X�5��c,>���MA�]#ȲU��$-3E���U�DN=��������4��J���R�V�i{�_��9�l�P	�����C��Y��/��������{�����n(Ԟ6p��I�����52q"�� qh,.A	uuc���b�S��ݙ' ŖAs��q���g��=f|r���^�K��-��m/k��2���uF�������s�j	���sg�瀻^N�L�����y�KXӣ\ւ)�/W����=��s.b�R���_����8-��C̀k��b�VA�J|��@sqK����vEB�~�04ͪ��Y�`+i�k| �� ~y��{�������V��o��<�]��@���َ�ԉba<Љ��o��i�H�׎�Ĉ� 0��7��g�� z!�j�^�a�A�t���ھN��֪��?�>���Bf��V��
��������:���1%=>�#�e�����T�e��i1���)��&|r�*�E ��=I�Sס�8g]7�u��eT�_P�I2:�K� T4�P�
h�pÙ��p$I��������A��Hx�X+.�
)k�O�;NzF��{!�Ӟ��T�(�m����^ѵD��/{��rza(#Vͩ�(���R�yƐ/��B�A�	��@n9�ym����F6Y/w�36�R�a��!"���s|�� OzI��n��#�yv��?I�I=�>Ne��:�k���E+��6%�,��$��jM\^���@.@�So�~���?=c��z��tV�Y�ڨ &�y��Q��[�{p)`��Z�tm��〄B�nq��4�_�ք�ٞ�'����y!g�ᝲ���9-y�8�捐�I��V^�R���	��JO��(Xp^)?��޻�]2G����<Q
4�8����/�������-���&��!�Y�YV{h2f6TI~���#�Aa�Wl���������[��:G��G��҂���]�q\k��7+�V������5)h��6S���?q�j�ɧb��N����2�׮1]Xꩶ�
7b��F֭��cۺ���w�Kj��4�ѓ3��z��c�-J������e"P�����$g�"��_$��?��Ԕ�������'ce��vMܸ�ړ����r<��%���&�I?f��(�Ap�Y�&�)�@����g��e<�U��	�OX��x,l7Wi���;�G��&�+��ݲ�E��f�c�䋅?� �m���fC��ic�$:�u�s����2���4~7�%9�Gn�)z��?���'r!�nF�g'��z�i?jn�K#�{�-��ʴ�Y�!��zF������Zl:�m��Z����G��9�%![i^|;\�C�Ƿ���迬����'��[kR�(w@!&��Ƨӽ3���u:�W>��V 	YM� ��J*��M_j��+�h���O��ia���-����&�9�ʴӐ<Xk+�@l�6+e,&��/�Cʞ��:��ǧoy]��dt�R�A���������$3>��I;&k���i��i�[.޵Le�R{��ʋ��J�6(dY�A,&7��o�lZ7(�4�p� e?�7%��7r�+^�=��*}掁A�N��dr4�ܥ�}l����T�d���VR~}CY�#.��!�5=c���D����X����\��P�ݻۃn�O�� O�	���yRL�:4� 9;E��c<��ݱ6d���{p'<�Dj~��ׯ�Omh7<�A��.��i���9�p��{��4o�;��&�[(�~��٤O�n|ok؉���|���f�e���k�3���RC�`J���
�~�����F46>��zv����PG�f�6�6g,8/F�O�m����C��v�w���̻DKl!	�n��l�Q	�W_"Jŏ�RS7��N̶��di��/��t����X�h&ͣ�(ke$��Z<�"�j�Lw�n;��[���9�U����<?�ڢ@܏�9gj��$\m�Y� c��o�!Jφ;H�'�G����"ծW��.����B�E�>�����)��~�&���ca�(�,�k\*���7`�2.��Z4Q|j�SXl���0�L�*B{�6���ѳ��XO�޹�>V@��Ki<�9��"�$VWwF>�(l<P6�\*�&��k�^���X�*����g��lH͹�����u�x���S���=Th�ĝ�_{*6�����us)�&+�w���1��(ϩ�#�g�!�$y2�Ƨwx�x�/�O����c5<dRh�.yN;�,��B�%ZcU �[����ݐ�	iXb�N�C��Uˍ������D?TkB3�2#N����߷-�=�1�`7b��um;ϩ���wg��Ò� Ǎ��Z��>痥]S�k�h7��a�7����4�҂����!�e�[�=�j��N4��&N��\���c%�eߗ�@�d�7aс[)� �P^Y~�  Ä<�I�Q�k!�̷�?;Q�i5���/VJ�3	gbm.~�y ��\2,��=Vę��L�=!t2��o6k�+g!�f&�]�n��3��^w`��t0�������>Kjs�:�#k���3N<7���sy�/��L��b��:
���]���V�b�������`$~��/Kzǫז����i�e,*�%��,�ӓ��$A-�0�+��^W�R�#�f�ddR�wѐ���j�&Ⅳ0(q1b��a/�*���L���6���J��m�^�����ͤ>��7�6EO9��_5�?ǣ���@c�fl4����Z=�墳�VE��,�{<�U9X�-x؄b#�{;�n�:Q��	�X�;��bj�8�4��7\%�e.��o��8{�+�d���vޓ=�n�>v;�0ij�Eݞ�aS��9�a)�.��ᘊe�.��y+V����zT�f{GDA�Q�p�6x��H����k�w�U��i�n/WŃ�n��L�VD������~H�ͺp�f��օ������z�5���t�۔	+愭	@s���n09x"�$zʸ,K;}�`��!��55����GF��ZpeG;�=W{����zb:�U����� �.��s�f�c�V��`�����5;+��^eC2B�:�-R�K�,W
^3݌�f�uC/���B#b"y��^fE����\��2eF0#?'74	�s5�����*J����Yy�i��t�|ٔ�Z��ƶ�G��5/�k�ti/��`��K�1G��C=�S����{�(�,�>���m�����8tR�Oʝd���U�qt��/uvYM��bJ����qZ� �Y����P@���a�+����q
O
��X�Ǌ��R��c��12�t�CD�@
�+Dݠ�ܦ c�J���5[e7��Y䷉ŧ�C�F���c&Ɇ؁CK�����\{��#�e�; /��Y�N���ޗehW�a_T�'H�\M��E�����;��kt�8G~��RE�@@��ښ�^&�[?B���F����-���#��5~� ���Y�����E�N>1}����;��x$僠
�ߪ�AH�e���;�g�&��K����h�8K��~	WU���uB�z���״ [B��O4�e�cy*�?L�|�K֚�cX��~ߺ�m��w���s˻�@�7��j�]�>S(��������.+�m87���cR����] �(���F���c+)��p�0��96����P�R0B���r\���n���@ԴccZ�"u�BJ����nNi�F��Cgy�FkVF9�yW;>DdyMsA� ��cq?�u	�l˅]?`�Ռ=����]�ð���pP�ò0�Q��]�r<��-i�9.2�����K��l>S%H�cY�̙�i�D�g�	�ۄ��[�����i4�D�^�7��	�]���� u*����@��_���y�֏h�i(�@5LSr�Ïg��m���ɗ��KUvk���H�9�a�F�4�*8��y^�:P��rdh�i&N����9T�R, �{���X�)�ǖ
)���߃�K���C��_tec���j-�?�-�dya�%���Y�oj� �ou,��R�n����́=ޥ$�Y��ߔ$����Vt�m���B�N	3�pn��_�K����W�nS�!&�Q���2��)��B[Ԑ�-s�NQ9�ܠ��>�(�5"Ά˨����B9:�P_���LS�'T]�~�I>NJ涮���1ج󐔥�gY�A	�u	��2ꐫAf��L��88pQ,f�>����BGbx��m�L�I�)%&�dK��/)�L���F�N./�N?;���V������O� 1����q�!P�Mt��ش2����3Q�)h,p�0P��E�.��h�;!KQ�wB�Jyr��ᏺ�}8;�]�/���A6w�������tZ��SI���Ӻԫ�������~:֟�5�헁�M��Bɴ]�of��o�X��b5z�j{��k8�}�����ȯ��es��9*z�~��_����A�����lEk��Z��O�d�(&�¿��ǌ+aN��`&���"ϵD;�#H>@����sksS+�G�O�]�7��0\�b��c�����j�1�(�c��,.���+��	|N� b)jE"~{YC����������N�g7�YI�s(:�%������w�"!���ݠY��4q���?��2&��^3��5$ԇ�Ɋ�+�G�} �ԅ��BKV��ADB�Kd�B�↤?Ÿ0��[ODTz���-���lr��]�Q"�Z�b�w�������J��= ^��EH���K�7R��S��ȶ[��(@-����d���
~N?�X-T���H��[@ma��H9���蕋��L��!R'��WN�� ��~5msR���m�
�o!/���)�gHmZ�D߯Bq}���DzG:���*��������k��uѭ��IN��K\�"^=���w���TZ����o�WF���^���ګ`?�'H��w3�d�e����>,�>����o�� J��ya���f�}Mɤ������0����KJU��Y%{��"W�75<���7ꎈ;�o�8C��rѺ�O� �"�z��D�J�V�8�����Y����"5/�?z����&|9?0�!ѩ�+��s"O�b}n��c�x T���}s���?�#�	�$�����º����
��Z%.������ԕ̔N��۵�䀫�*����-F�؄������h������Q�^(�&dt��c����[�c{&F��w���^���7�m����ц�v!�z�V6z���P��Pߩh��`l����ec���m�Nwy[�j�i���O?K�AQe�+���y��c�����y�$�G�F���o�-g��(��D��F�)�2r���5��q�J��x�m�/j�1Z@�7�S��`�Dc	l�H�����Ц��R��y\��w���v�JЍ�v�K�P	�-o�"�i)��Up.��-��G���^�o��~˧�Yb�,�,��b%�+�_0[�53�Y�Z���8�w��"�i��%Ӫo����Y�����m=w��ՠK�1����;!|el�Pr��;�8Vll��_-k��f�%�;�ӄ#|��?d��q?qY-kK��V�d�;`5aې�8CZ��%J�ѿ��6[���5��ŝ'0a�)�����A��R�@�wf������튝pa5���N��,0�7����ļja9�Ʀu]�-m�.�۲}X\���@L3����6}�g���,�a�˭|�F�U�Y�F�2�kSG}͈�!:�@�5�Az�2�d�(�0�%]5�uD �u��JLK�o��r�0��,"�1�����ͱ^u���غc��.�H$y�}�dQRv���J���EG`��F���E~��!Zg5�ֵ��H]�P_ �TA��QL$�I���Q{e�pH��x3ڡE�)�~g�jK+v����Ll�{�����	�M��%���\���T^p��//i3�����&{!ѓ*�Α�Y�d�����FIWf�S�S��$�v�SNktX|yb�O)�++z:�Qj�8]���x���!ž��D/��]��ۦ0m&�������cR&;�?��~J[��:�|s+x�BA���YN�u�}Y���.7ε��5o'�~e��V�����-��^/��lN7"��rX<ӟ+��gV�w�����Ae�	ܢ��$^B��0��y�D�59�Z�	��&�^���U�ܬ��}r���ȭXs�H@XKxբ����o��o������l��c�D���J����3~�sJ���X8��.>�.�Zp�pz����QУ�#p1�{�g�
�c�`��o nMpU;���S#�ݶ���|t��/t+Ω��N�����q�>8^�S�~s�9�U��x�(�6<"�y�K�d|˓R�]�Pb�r���I��# �z�NRD`���N�	�5P��kK��1��J�w�
�۱I��8RP��!Md�i�1Z��< 0�oH������7	���͵-�7�tt�69e��^�8������W��$ &��x�a*��gG�cfb�0\8e)��s�+$��Fg!ΏU��r{���!�;�&R���m<Y$����-v��W��ǡJD��ꎠ�� G��5��yȚ���5<aO���ĳ�	�گ�r�xf�y�i��oW�%�fN~������1�o����8�������Vf�ZD�E�����X2t��v�ZJ�l�^qq,�C<��m�����t�zRS��
��H$�M�-���1�����L$���R�����[�6�ðae���-��`G0A��0����VA�N� ��D�o�l���Z�A����́pW ~�_�%r�z[�f�ymd�L�N2;�Aǰ�i�8.�RZ�#�`	�-Z{6����O��U�`������ю8U�0q��YT%���.^�Be���>��_lP. �g���9X��¡=�#?gxŭ�����������<a��X%�N��T�M��+u�q'�^/b�����.Fv�-.��>ʛ�/z\�gꀹ�����Fd�����{��KRx������Ra`0�BQ<Q�t
+�b^�E���"^ku򾋠n����2V_T���%�)�6�C5Ӎa�%3�SnRyB�nS�>�_Bǿ����5wɳ�t��tu)�$#���Vf#��i3�3Z�Z �b���?�����K�]b��I-��we���)B�R� � s0J�_��.�*��!����G"{�[��v�Ҵ����u��:KC������+S�m�١r��Ij��X,HG�`��N��T���ybMt�F�0a=��H���)�m�Gڼ�o��h�cS�{����i���cK�Y�'��!��A�%��RwO.M7����3�ˑ|x�����tt�~�(��_�����YYu�HD��G��C���YDC�gZU�J���ndQD�����k��̏HY�"f~o�(�Ϙ �'�Ja^�߲�k��rP`��N�3(Eo���6�Eo��'P�?�qP����tF����o ����d�?�k����D�MGA�������k�)L()߅�Ր�]
�W�=b�c��ۥ��v�S��2�y���b��8�ω�&��S��^��������0�3<_È�R���UI7�1�j�0��3� �]��a��S���z������٬���'��=�#�h�%��x�̳@�T{Q�i#fހ�Ց��d�o�ټY�3���aH�_�U�r�"^ո:E�X�����^����
�1�=��y_���=nQ@�#@&)��������;�s?s��:gW����GuSˠ�m�@��5RM�݇��؍|R/0�~7b��T�v���S������p`��AH����[5�IBm.5Rw��M��J8g��~�Z���P8ot$G��̺4^u�KR����R����@�|ۿn��%��|�pm@
����#�W8�s��ɂ���dϮ�$���Z-�>+�_[��ó����UP�Sҵ7e:{�r��s/�ôs4�m��G�nKAm��}t��O&GJL�1�� �����R�F�5�j��A�	�raI��S�x��b��]/n�0G-�6�C'�5���)jf悄#��@��x�[�$!P#���$�����n���3�����f�4v`�g,+Z�~�ƹ�En��� �ﱿ6vV�3�O�*���)x�Tp���ւ.Ḳ�ZQ��ѕ"�03�}l���s@@���ۏ�4#y~�7h߆"4��9c{ϷZQ�'{ZFgg��.��ݰ&��p�n�l�qȋ���7�R�l@]�b��:���/t�{�",��ʉĥ�'��6J��XЙ#�u'���>V�Í����#a�H�f���)��6��Q%oz�M�;\;2[ψ|DqG]d4o�y$�'��XA��� ��lV���s�=�nW��Ba՜	�~-?ڻ�c���0�IsY��&�P�Q>����(-&lĞ�5wƜ#�MWv�i��#Pyhg_����ԋjȬoy����5< dl3>���5k�K�D?'��VR�{�P�'Z�>�,-7 &�	S�J�@�	���	���K�RY��𵉷��7۽.U�R��N�DԢ%��#�I0-~{j��[��o��R����;�F}�����ӫ��U:�?b�
Q�r?��F���U���":���#s�|��qv�>M������xM-
vmK�]��ïE�G ��.F���uL�M�b� �����AW�F�忽����]����uB��vt�4����cr��T�g���ǂ��^����Q���Y����+��/т8��[d�pt��Ar����pjv�t\��X��+	P]s����>�T�D�v�-[>Ɉ$�<f��}OH? MW�������3��š ��;N}�*�#�õ�����%X;�g�,�Ժ�^^����+�y˗�W5O�c`�qDV���]���F K�cx��۞�B��G�r�ދsO��YKf�l����%�p!U��?�XÝУz~���Uы��`X&��F��VxV��j[B�k�r�UPZɹ�1:q�GZ��ּ�f�a&b��(�X�"~�6Oo<ӌ7>���>� �H�Z?OX� *{-?"�f�o5���}[��M��j~y�t%�	s#5���e���.���c�CJ��j�G�N��=VPUlwJ$��%66���j�"(���܅�d0A��T�L1v\�1G
 ��.�b.�wr��O�"�b3F@D���"g�W͏r�]�C ��m9�C4�st�X%�n�5�l�K7Ý]�N �j��mG����$#�V�0Z�bɬ����'.<{V�Rk
�T���;�o(�v�l�-čG6c�C}M)t`�?����փ .��n�(��?�F��,pD�<o5i{e�9�2�gH�z6l��Dhx��4����:�l�!�����)�ĸ/H!�W�~J�%�������п�ik��[��_���Ǧ.l"CV��v�=X1UӶ�$�9<�,��}�~U<,I�zRBS#�x�ro�R���7ҁ ��׀b`�G��M4��D��&��z�8��+���KM��P�|J�"3�M|��]g������ճ{��ٞo<O+4�+�I'�������x,9���i��M��nYb�Dg�ns6l0��/t>�Z�f�v'jIP*Ý@�?�G�kKByTFXUT�D�Dss���򑪁B�g����=,��� Lv�X��Qo�ì�u�p뺠�!���g�l��+�4��׎2k��N�^�4&X��
�~l@����N9H��-) "NQtX���K�A�]���r�ZiP.'Ϻ
� �G,��K����v�"�z8��{̧j}�>Z��U
�����%5VI�����|�Qg�<���A��/t9wi�|Ee�����]:n3�龆�2�&H�s�83:2���ˊ�+_'��+�^J��p�b��NB�$��"�B�^�!�'�F��{�u�!m
;{(�w��u�*��m��
4?|���ڲfVˁ�KZS��)�>�|L�AKěD	����y��$8N�2�rb���9��a�<���-��"_��&y�r���/_�mv0ym&F^T�A�1,�]�N�Y��/�rh��81��4lD��+2@�3�P�L9�����n�M��dTG*�!��iٖ���!�x���S��� ���g,�7 @k��Ȭ���dS�C�0e@U��-�֓�'e} ��M!�F��KZ�~W`(=�b��L?���v�;�]�V��w��:��ex�d�Q4��*?�L����P����]Zܕ�_Tu�D^Mx��..A���K��T��&����V����2,�ihz���I���w��_D0�NPX<�Ij�j�Xŀx|�]�_^��RM�Y���2o������c�gL;�L����-.��J�������`|i_�p+�~o8�$�0�ɢ��7���`�\?u(���$Lؘ9����d<�T��mNhs�h��C�(�4���*�"ɑvӜ+�����Xi�[KW�J �9�{1cήE�E)4� �F�U�77���>��N�)��[� f��iy�X��6æ�(ڻ�i�^�q��Pb:��vw��DB�%X}����r�?B�3���-���Y�%��迀'/fu7&���᠒�1�s�f$�'l=���6���~��^��,����C_vzx0&��̅�A�f2e ��]����ŧF���H��m�;�Tss��܃���釾k����{,���FF��k�q*��\+��ߓ�Dؓ�>�8��Ɔ��<��t���b�!�xI
���U˄RеNꡞ
*N��z��n��;�<1�2�v�,�;��zi$�Ȫ�%����X��)_�v�3��v�׵O����KK�Bj�3g	H\��Ǐ�܃��g��u2'��j��:��F<~G���E��2��܏�1y:�~_� q�;�.�O=��E��oj���E+En�����9���<2Nb;�@�@�g%��pw�-S�-/���G��f ����BC�׭
äF�.��2�AMIʉp]&��%���2������DH���3==u#��y}���ό)��h��7�5Ō|:����k��׮�p���f�1�Pꉙ�{ι�����7�BOs�*��)��a�Y#V�ءC8ۡz�6y����Χ���s���&���vj�$*O��pr,�[s�ܥfj��&=��(Ϸ����N�,�᛿.&���`^��L><�`Q�KK�[��D[���BQX邽��F��pu����GI��:��i�'t\zݼ����tA�,<�8Ճ�xˋ֛!�^{�7L��.}s0̝�?���\�!O�Dy��	�oΈ��)M��{:l���#tKn�m�;�ȉ��\V��:aAhڱ����f[�c��*LR�S#����#R}����`��x�SW�����X��:�v��4���M�K���+����&�2�&�!�m�N2[��.HVy�[t��٬H�Ȫ�T��^�H�m��L���bn:_U�k��K�_?u��F�������c%���W�?��ָ������E�B;1�/��Ş[����֥�0��1������:�Q�ȲS�,�<>l�Ε2�
��E���I�P�+'�7��E��yN��eK]�����a��9�
kץ�������j&+3ip�gN�����㫍y�T��LΪ��֭k��`'#1M�q����	����T>d�*D���Cwjk��(4�a���|��(=�$�~u��f�����K����ăI�C|�F
`������f�K�^��ӈ+ھS��-��Q?��L~�3�����TT!*�0�ꯊ���5�y�lu\i�$l��}W�ف�VT19��/�.���/b}L]�zM�,#�ċwi����t*|��1=��&��g������x������`���|'��7��j�w(5F����
����H����fC��Ԩ�ٔ�~ۦ���gPYzx��lo�-0��K���e.d�kYZ�]�[r0��A}���ʾ�פc$���ᮥ�~����}��P�V��X�5��U���C�Җ�ޙ:w�r�������s~�tL���7�">�t�^�z��>̾�A�g������>%A�$GB���ժ��[#��]�
ő��T���q%��B5����k���Z����FC�[h��V��jR/� t����vCs��]q�a�v�Z�݈UP�C��Rj	�aQ�?J�KYL3���g�"�iVFF)�b���e#����-���Y�v���+�z�P��s���3��a��Բ�JTL4�c�
�ǩ4�U$�NfF"'�a��0"���%��GlE��3/�j��4�]I�r�TYq�U	�kg $�>�Z�2��xI��0-��wf|@�Zx������Hs�w��s��e39�i4�+��!��9�ԩ����a�;�5~��j�������Ot����Jr+����&(��*���N�?EAGZ��;��c̗7�=�����ó&�8�Y�m~��"y�5��*�q̓� ����jɝ�'�4<�SAi��/�F���$�2֮
���/D����o��FA�,�7��׊q�e Ǜ�p�&7҇��C�{Î��Ž�L*�R���]��07]�l��DG����i
���*�g����ʽ4?%�Qh�9���lԻ��l\ʥ�v��!�2l���M>�R�*��槐����D��-���6�'��A��~?�W�Dښ9zX����h�M�	���|��>^7?�	+*�gb�zzߪ;������AcW95����8)�.����(����-W;E|C+8Vg��u=�6Ϫ$u��G�ϬS
+79����]�=~���$�
��]�(�Q�t3;w"���}_��b�ҍ�i�o�+�0(F:W�iy^��P
cw�dd�p�į:��+]^�a�Z�Z�O�
�@pQP|&|����s����@��/^��̹9"�����4BR���MI�7��r��!{�ە��刢��P+'�>r̨{�i�����Fےޥ��g�a4����.@��e`������3�o`S�j
D���2@�?���$t�Ӥ������ �����P���l��\�BԞ�T����u5�����p��b/�>��m�И����_��F�*{�^@������Z7�D�m�a�q�,���s��ZM�� b�\L�vn5���!�����bmM�����ńt6q�u�8��%Γ�1t�T�"�1/\��y<{y�/��!��Ri3����P���pW�,w{>�K��n����έχy5(��Ò9S>z�-��������^ՎBs��r0X��!!�i
��~����QD��sP2���� *���_]"�:,3�]��>������Ս��Xx�π�E⌍D��B�� �2k��ri���ƮlH�Q�?���9��U��͘%��lϚkɎ[��B��VUl/�EU� �&�W�(�Q`�?L��}(�QGv��|}"���n50��U�]14`�z��(2�|mB�ī���uz�@lM�O��ֲf~�������2���Y�����U6��y�:����w�^o�J���J����(�bO��@rl�m�q8���B�?�e:j0�����݁��jaf)}ѽVV�@��j���7I�?U���f?�*7�mqio#�QE�Z�a�\�l�*\ J��n�Uk6��Ջ=�O�k���h�1e7jǐ�@eZ�F<�|e�ا��@��^ڣ\#*=�Q<bڤy_�dV9%%Z��K0�W�3�'�o�X���m�	�u����h����0���ˁA��x�UNi��/�X+�������v��>k�O������(^�'�k�J�ܱ䴋����}���X���Ԙ���C���9�V:��Q\KbI�[��%�W;E�AA���)&�Dv.SM�?&��1aK������9^����*ӧ����s��6�J��_nk�M 8shX�b���a߅S�
���颎s�y� �k�?��(|ei�8&(0!zK��<2L&�6��|�f�����OQ�j��3���&ʦ�<αR^�/�ȵ�3pˣ�%�>�U�gc���p��1��UK�2Z0,�TR��L����S����r��ϣ��:n��E��aM2m��{[�����T��)�$-��%�9�i�ȥ��kj�T�8~B�_��S@A,��*���r�Y*�=*�6Gf���K�x���E�D&Fڈ'�y����8�� ��iD$� ��8�ϰ5i�3t����vaȭ�q&ͨY}+K�ܫ�vJ���A�� +wyy��V��T���H�k�Լ \��)cxuA=t(�yQr��z�H����Q2���7�3�P�īm#}�!a4��֩	����l�$�/Kբ�p��3���T�Iz
����o�鋣J�&C�"�o���
�W�P�oI��/)x�Q$͞I�Į����?�
�o��*oq+�+� {�rT�rU�j�t
������\��|����{�S�5&>I��E#�<��j�,�xPYT����B}����M��Ǚ��J�tI�����e2E�a���o��C+��H׆�~���w,��h��KX�Z��^(���eho���C�Ϗ|�O�,�����{2"�a�^�*?�����5�D�_�6#�;+�<!�za!�6q˄�\�$EX�rp�W g�gn����.��}�&��{����շzZ
�h��h�^�`���s���Kj������~�J|t>� ����W`�٫f�9�6NG ��*�{0)���2�!*�Toȵ�h���k5\lgg��������`�+Za�[�Y=��ǣ�xߪG���t��
�w:�bȤ?�O/p���8��o�W��W�2�/"�D����S��U�����)n��`DY=oh�`���ګ=�K��^X�h��<���^!��x0�3���	:k�6G��%U�<Y��������Kn|��˽[��~fz>���i�1!3֚�Ł6�	�X�������CeUjd��ō�G �$P�
h\������j��]f�,���ֶ����D�"���:$�Z��_��7�B{�8)���q���&;f���ҵ��L�a �Av��CS�^��2<�ik][M��A�B7��y�O��Ԇ�Zzh����=���ے��+ܭ� V2�����s,� �����BIH��*�#~��R&(KPM6��bX�AM�x^뛪��>}gt3�뿘1E(�ʧ4�`cUsM�V�l��'�y���]%�n�4�щ��+���0��@��6�OX�q}#l�#���`�J�	���Q3���i���"W��A�lz�;D��
�W�xS�����ʀ�Bxhz���K*�{$�h�\O�kS���&9�9V��ו����H%ԭ4�zr�&�CS2v����w�����쁀�R^�Q8�*&�cL� �*�'���V�>�<^0�L�v �������M!x����1��_Tۊ΢+�hX���̗L�0Aͺ�Ֆ�YM��&�)�D���  �B����[zD �:��c�eI�tϨ퍔x?$.f��TPFZ�L+j��H�/�Y�oQJr�y����hޑ��ls'���)�ܯ�6z��+��댉j����)h�Nz��3tf�|��%ÞZB�:�԰��A�˵ez7�<��N�À��+�3�n�,�%�s�^N)~f�g��g�d�h7(߀�v&Y0��{lS�@�:A�M;$�\��x�Υ�H��*R�*�X���sɴ�]Q#aB�u��B܈G�W�m�OҮ�T�Z���â��$���\צ/Y���D偧�yU(ڨ� ���39/�����&K�P�9�eP�]�W)��x*�9��3�<�ؖ	�K�v&���%=k����3�N~���i��"*��h�D�u�4ZPE�$?}���2��xKAW��$�z��R/ӑ�\���֭$Dʷ(�u���P�act\���?�
w&yE���w"TztB#����4���̇N��"�->��(ĵ�,	��P�A[]��U8g訉p���ƀ��:�#K�.f\��L'XǧBj(�s�T�\-���H;���k��{��������P�0
������f��q���2t��K0(���`���i�;�gc�|ǀ:	�	�YD���G���F�o�z�T�xc��l�!�S}X.�'�G�u$�E���<.gw�x�v�}!Э�8����VJ����#�=a�[& �<)�'�s�hTʥu�~Ƿ����_���#@ݾ�8�^\���^�_�bܱ�es���*G�������n��A�ҳ�6���r����4�L��hH {�&�?���񎕊L;jc
=���E{����=��3��T-��ZCܔE��A��ê��N8�������=���Ah���������HJ? �/1e�2��qC�]��ӊ�#I�W���|���;%�\H�I;v ��Z.�[�AAb8#蠆�_T�ir��=�[�.h2w=!��!��U�E���kx�3!dט�2��z-����T�a2�����p��2!މ�� Ͻ�����T�U7˙u���B�dW�d.��K4*�;Mc�����L�H�&~�7n!�c�PL��Dݜ2.>ׄ/�_���T���м�h;��aГ������Ơ��$�zy�-5
�#����oўm�G��%�_B�a�Bޗ!���*�����ޚA�`����hg#Kz���I���DMֱ�N�ؼ�U>W�l^�!���%���9����?��&��P"�#3R�}�kN�sQ+D�V�?��l�R��drg��T~5�9��L�V?��l�3����`nݔ�m�ZE؀��O��6Ҧ��P�/�5���<�	������։�bJ�d�艢��e�!�՚�_�I���o�˿P%	P.!������Ej�2�peƺѵ��E�3�'��,�����K*�$��d�\���^ǰ�ߍ�>�֧v�z�~�m���,.�
�E����m��(V���w�I:6�Q=u�3��w�|+�F�H�	,�&B-�ע��Z����h$�99/W׆��$7o�^f.��׼�@;��К尚QR�.רoQ��;�����d&�q�����7���(7!�+s~��O�-�X�)� Q�Yu\��gl� �lDi4#���;�W-*�J}�9�р���Y��)���(;���4�����`�@�C�=Dg���&�4x��#��%�|��7���A�<�U|tAL�Eˢ�4�:�ѻ����5B���]:����D��ݶ0Q{8�zmk�Za����_�z�ZZ�D�1������
gtx�;���aϾ�m�%��r�;I�6O�g����?-��d�W��Ȩ�G�D<V�">ԀeGPM/�c@�Ş1�+O;�H����`�T4�b'��X���GTX��@V'�8#G�g��U�9.�U�yd˕O�Q�K!"�T&�o�6�c����M�����RY��d���o'��Yا�yl�cW�w*N+��dD�3V�v���P0#�h�e=�i�f0�h"�J7���A�#^�n���]O|%�A�jMcF7�˥!��z���q[�(j��"̇;�)���Y0[!���&���o���i�c6iD�d\����OƘ�`��@�����D�.[���Pp���8�D6KE�!��٦��qj��]�����Ҭ�����=,��sA�����񛁜��	�l��W�ux���GP��pa�y��G���T����O/���:	�4�ڜ�a/��Nt	ې�N�8��8�`1h��bo����Tbf�w^�u:Y7��(�/`C��[��	��[WH��n�ơ!>�吙�xͱ��>�!zu�/���t�����=�c��K�=9/Fv��oK����cTqZ����*t
����d�.�����>tGQe�jU�D��=�6M�$�`ٗ��oM�y�4C@�٫փ�E��h�>��B9��u�r���X[�+�T�w�6��%ꉜ�gv����Q<VPŢ�Et��7Ә� ��R>����S�ny��aH��_m֨ �V�j��-�蜿諌D�:����ϫ��^����GB恨qzĢ*��%�������SM�ԋE�h�r$�J!�����t����������CaΕ*�]q�~z�����h�`k���ى���rG�P�RI�%KK����t?���l1|�n��zI�R�?�˯��z�*��8`����u����񮩮9�X�E����-_�ʄ�B�\I��o�E��mP�0�b�.Zc�VH�K�����8�&Z�?yɵ>Lb�g��/".~�㞨��-K��n�6�X�Tlr(�n���X�y����Q�/��~����ζM��Q��Uߞ"�*�U��P�sR��*���.0�@d�L��Q8���t}��f����q#ϰ��;)B�R��<(���9�%�U"�l8y�j�+i�o��2,Ax��+X�<;w�S���2�������P�N�O0�Q��c���8��^F���׎������_���Z{ok,0� ͸�����U]٪%�*}��ŧGΒ^�xo䘲W74�F����t�=6���M�-�:"���>�R\
g�"U�lk��4�7���"����Un�eb_���߬&� M�Ű�=]tߺ �|�����i�4̛C�t�h���5����%υ�"�:��UN�;o��F�p�����4�f*��Pj�E]���q"���꼀汙�_	yj=Tb�wi�(�GJ�{�"��U�!�Q4�|V��Þ���Cz���ٮA��ڎb/N��K�I&�v;qlk9��!���.W��~�k |̿F�,��0�|� F��ځ�|��6^�zTS쥵�L��Yo����9d<\A9�Re����$��N�\�	!�����L��/�V_�Q=��6��.��ŏ'5m�_<��`�4�h�*|+�O��0��;���a7�R����j��^/)�f�2�Bv)����WeAg8�w�h�$Ti|a%��hf �u�:D6�����|4f۱3bJ���G>���g��ށK^1��0��D<W�4ܣ��"������a�eG����`M�1�	�na�d��<�Q����y��J��mH��RB٠������2T0�98YH�\�"��3�SK�jn���N����[�P}��|��_d⭙,L���-$ɺ���8��ݟ.��_���'A�����TȠau;����*�G$�x��&2�M8�C�id5+/w�K�6�!�($��$��>�B��zd���9=� ʭ�;=�,�K���%a����=�"Q\ߨ�Ȅ<�\K���A��+��-ʷ`)X���5{�G�M�Z���W�"���3��mEݝ�fș��y#��s���7�/�M�w�p��R�ga�~��j�Ȝ�J;	Z(�Y$( ����S���d�f�(]�ѣ�q���8^�\d�;B��Vv��o�$�ȐЪ���U^����YN�F%b��g{r�`<an��dy��o���6\6���G����Ƿ�s�tw�dAYm��:!6��#��7��"���j��>+��w������q�*�W��E�P�L��S�F�.PQҠ��I�^<���c�;&ڻӁl_)ۋ��ZЫ��ų�["�'��,���ZV�����c��߳��� �f�^/�A�q�!�Z��kP��?�P@?�~@èA]���n��ڜB"t�<��������߭����sV�Z	��7��xECPA������F�� ��X�M%;�7rdL˕��||�e!U����x�[m�[`�����7�!d���(lp���OS��>D.����,��#$� ~�����P1��x����5|!�����X|1�A��f�i'�_� ��ӿ�\�`3�����H��㇩�ѯ=o��
��^C��Ab)�.��^x�m>��h:ru�K̸��DI0�ˢ�7L|Ţ�*����)��%k>��y0�z�%�] ��/�%�9�黶�X��s���tG����UډS�"���*3[�y]�-�o��&�f!f+y����ޯ�<��A�S��%����?w�&�]ə�spS�0Q�DR3�:n07���n]����A�8�J�5BK�B��w��7�P�����6@�x\��'4��3�Q�faB�a�ۄE���<>p�ƃ��1��iD�x,���U�E,�c@��L��g�|	��I{Z�}����w���d���{Fm��X?�9-p�K��H�+;�$�gf����nqpiE	vza.��Z���V�k��>��]�i�����!��9�+*8�u� ��!�Ch��$�	��ىZg��3�TE܄�2�g'�����X�0�I��=8Q�A��1@��:��p>�shƚ�X���$�n��	�H�y���_B]	]Q�A�lU��<f���
�,0�Z)O�O �	�޼Fh�B)�m��;���`�g:ư c��������K���u�4k��\�t�}�	r��eSNf����O���4
�J��W���*I��b��zaCFNg��l\�G;"d�)*�S��;�u�?����f�w ���~��y�b�mx�/ܮj;��Ė?v�c�m��MY�F���j�7��J�/�>��+ǖ��1���!Zq;��b��3���2i��
�S���ʢ'&U�p���Ź��x��t��P��c��rcʌo{ؔT�:�Y�N�U����^�NKjz�s�0�.�Y�c)Q=����M����7��JE�m&^�tw�	}ri}"LZ�jĩ�2'�]�j�V<�2x�Oks5�*1�'�D�ix}ź�������N2�9�E��u���	p��e�|�1<��<ʵR��N���d��&���|��Ġfv~P�A�s�K��'�0����;7�f������հ��{��PM9\�13�ˡx�����XTZ���tpC� ��Xh�2(����+93��ۮ�U�(�;O�NS���Q���l�h����'қ���b��_P�٭a���7*�*T	#�([L��6<��E��� �r��
�>�Gv֫ɓKC�v�@?�w����T�4Y;ˎm-�S6XA얿�Ff�gj�`c�XA3j�]j���\��������k�>���I��4�}2f��UY�/,��9��ԃO����ݞO��V�k��y�Fg�kmz���X)���ߗ{Z�r����/y�[�`@�Ls�`�?�f8_Sg��
���f�݁I��b��څ�����H��W$���c����$tO���攐ؖU��`{��ɍf��zt�V�i���<XNY[83c[:_d�  ق�EٕO!������=cmV�;���jj�ܵL/ 1�X"">!K�K[�	d��E~.��J�U]:�����>�����]�{��3|Z_SR����6�����6[�YYl"p���W/��W����x1q%ʺMrrD3̽鼩"!�yRXX�D�?<��ωe����+y��
�r���F0E�����!}s����8x�B`\H?Ѿ:�ށ��e��S���.�HϬz*�E�?v�[2 �u����|Y`�]'
�5�1�NJu�S=���O�&yÄfH� {R�����^���41�_nf3�2�����U����§ho��dE�ƹ<ϕ%�����7�� �4]k���ɘ^$�Vf>��wc	})-` l���B\4ej_F{��w�A��óestc۪ ��p�+���*�`�� ]�فÞ����L~z�$�	И�s�|�$�P�ڼ�\�%�;��&�#��YN�]K|����u�����D(���/^��#����`"ʐS�fě��5-��+U������`�~�-�E{�a���0��,� cF��w0�o]���I�.Q�t]��<��Z�(%����$.V��G:Y�饌���&wZ����Ҩ������Ņ����^�c��=H�B�AłϵleGY١�O�r��U���]xD;[X�A�=~��r��X2�"���k�R�TyZ��)�Ǵ=��D�3����:+^M�v��+	Q�����*����@�ڗY����bB)^@p�Ч�u����*ۨ�fW֪�QcPq0Y%��m" f[ֿ�52E'�]��Cp<�o����&��Qz6<"�+�zO��^�Ի9�&��11�\N�������=�Z;%�G�k� )��*���a�>�R\�p%�e����-9�Zo�\�x�q�T��'zr aZ�G�'Vo�ʹ�L����rD�llL�Y ��/���ʥ�G ��&H{��ŉ�6�-�rq�\BrN]>@��xgj�}vh�nͻL$VN�v ����R&�֍'���N����So�N.)]~(C9i�K��M�3)^�@3$����o9�c�|7�u�x\0w�5Q����~��I�n_�?t�EL�	�_��\�iB���}:%47;0Y�Y�4�!.��4�$۱�;��c�W���/ �ː:#����Xw�Ҝ���3��}�b0��21�B�Ѕ��ZH̸r3��Y�aE4�j��j�#�G<wZ�i��j�d�Aa��	�	|A"DVǤ��a⚚�֨�:5&�<�D���T�#G1��zC�z�>��l."�ӻ{��K�%Y���J�uK�K�/9�����t�4�i�L'Q4l��М�e�\�̇3��x;��{Mɳ3C��C�}}$�@-/�~:)�Ce�Q��H1��ܒD2K���f6&�~�öL3.�XO���z�@�J�A6��Q?"N��E}D.�k~�+��:��6�WxD������'�E��:%���)��lS���Up����������F���a�C��s�{m�o���y��Pb7l���_�Z?���U���r�剕+h���*�Q7�k�'��K.�	�f���FܙHj���G���]������QcԚ�*� �9HW�cw��=�\�����&z<��3�m͗��JU�zΩ��Zd�^�~5[�E�yǐ���Ɩ�(E�񬣔�`�o�gp�n�|b_zvD��/�}��y�5ն[�tK�'�6��J4����� ��݊�\[�\ҐJ����#��_��r���s ��,|/��P*|$7,x]w�x�u1T�J����uJz�_k�S�-���L�ń���5vB��x�&�SN��&hN�9 ���nH�Q��|C�%dI]��&"��w�	���������.��F�ǂ���f�� �kă-��R�^Rd`�nOV��v*����{\�<�co�����?0
�Z�"��k�!��
XZ����|�$A2���Z�^�? gm�u]�'��1w���!߀=����W�#�7���������N/�E����O��"�!����]i�h�qR@)z�����N��vh�d�������$�`!�8��~�V���l�i9�ـ�)~���>�,E9C�f�ݡ�%�|9��ksPo����Q�W���U���e�eea.S�J��ɔ%���M����<WR���v���8ߩv�v*:]"�g��-ʈ�;��R�:��I���q�Ogҙ&1_��0�M!8s$eJO�b1L��ة�l+8�}@OE5ը��v�Qm��`i�l�g�� ̞��> �r|=zUnUv�u� �fP����I�ׁ���������7���Ȥ�8�r���C'�. ����G�@޶Pw[?�W��s�n���9��Qp��t��ǣ�m�{"��:���8gNM�Sݰ#O=𑥖1`c����h�Lt`���5� o�*���"0��������[I~F� &ogt�\��:
�����!����5��	'�K0f�a���9�d܁�^�f��<pd�n�R�ȍPK������'b�V��%��<W
ewW��Z}=��������&�J>W$��m�[0?׈����ɜg�W�><�jb�z��^�EJ�*I��������U��\�k1�hAʼ.��'6�C�<�ÌY��T�V0H�#ý����b}E^9��*rS8�޸Ҧ��n�Xj�4����V,�-�é��wP2Ж{h��N��[�����|�.�0�d�s�KZI<���z�`��[���r� ��S��a�`:z%g��n�,�DY���>/Sk5U�RnR�9q
�ݮ���W-��'�-D$ٓS���=B�uG"�t��X��٦x-�J]'�V ÔsZ�HT�L�� �n���n��<'�!Rs��G���|Q��wP�,x��n�`�#��H���oH������^/"<����g�//��|��k0��T����2lBf60�����%��]��wI�@�.��eK* ��q��B�r�p�M�]]1ћ�a#^<��p�Oȸ�,،����jk[��f�Qb�՘�Pd��7�CdAg��8\-pʩ3����r�l�����J�[��>��0����O���z�����G�
�U#`�p><�ȩ����+��M��G$�m�AzȺ)"��Ѭ�5�*n�|��/���E��""%0�2}�xt���3Ђ��wY�ē�+s�N�_�S�y̤���)���a��9�Ƞd%�M�<�ew�G����"�I�w������W��sF��9xC2,:�R��,�ޛ_퉇V����hoc��Hʬ��DFOHK�vEu�&���buv�fv&��k�Gn��9� ,S��:
U({6���s���o�B�%����~��EkGN�! � tC�/`�B�9^�*O��ה��aY"�q3��R�����С ��\al����X��~l #�����C���-���b{��cz�/��w ��������fF��K�%{���+M8�N��^�q��U{ʶj��&8G�UZ��Y����Z�2c��c*��7�Á�%��*�NV(�4�϶8������}?�ET�K"��;��h0��R,YJC¹���`͚�j�(K�A��R��I� ��P������	���B�p]�.��G�B"�>Ý^�n�N(�<(_�-�����|�U�F�LigV:Ђ)��>Z'���,��mbcm�T�@��53��g.^����H�H<���؛�:�Y�c�(�.��C��BI 2dⶍ������r[��Xː4�����`5��B��A~��><Ą�J�{�����xV� �f�����7� �%J����"&MZ�Om��p��6�5�W�@1#�X���g�,�:�S����:e>��$u�Xz)l?��LM���^1��l�zl��G�0p��J�${�M䗞E�bJ���VL���u���<�H4~ ��L��k>������*�'���w�b�D���Ζx�v������o��A*=Ե���=��R2Zj(�W�7���u(��^hz�T�O�LC�<*Ddl`%�i7HL�3�v�SYg�-���_{��?�<#3[�V]�N?�I���f��`Ź� _N�8W/0�U|�����q��}^@y�Z�wyQ�H���{�|$w��5�H�az{����Rd�����p���t�MEݠXU�r���1����
Cإ
��}QCeJ�T���s8�Ap�ێi��ӿ����n�7옜(vA[��Kӡ�G���p���y1[zv�_���?��5\��U<X�ik��Tz�3h�-���4�~��׌��X�Ь��{.V%G�"�m��������h�}7�]MCX����v`����ؠ/ަ���ӹ�$��,�ݞ�3V���i�i��I���y�O��t?b�p|���$y��!���m��
ⵋ
&��������S%x��re�]��l:����G�,������˟�����`n�d-H��0��տ�k��V�F
�9�xdL��������[JD�������du�rӞ��.C�[kI���C3z��ږ�h	Z�]�?��?�F�~�ų��k>mZ�����vԗ�>Ɂ�+��{}*��o�P�6���y<��^(W^���S��|�&ډ%���4xd�t)�M�T�B���+��'�^ř`�"�Ɇʙ�X�6�3�Z�X���}��V��4NMŀ������E�v��x;bZ��������:h�AO���/�[ʡ�Fѧ8���,�q�!�be���T*����h3'v0���pV����]fy����߃�ڃ��#}@o���txi@޼!��ڿ4�\�����=f�]o'�Į�N׀�UT�w�CKhD���� b�c�ÓM��� eK���k�'�.���İ3�D+B�?��K�s�j���Pk��SZ<�kM���L��f�P)c���t���ϓ!s�N.��]�T8������x�1̎O�뮔�/{	g*��'Ix�v��d��N���$�����GW�n�[=0�b��Ƀv)��1�{��V��q�Q�~��}�'���&�8"x�O�&����Y���]�])����V%�t�>�`6pbe:�/xr��_��r����v����?peXX~,[OBf���\�>L_v,�/:��,�ϥ�8�?�+�\�ps�zb�(A!܌�֣̯��K魲��&#������8&��>�%�����G���������x+�����'�6O�P�~�A��Lh��.��/�������l���4a)2�x��F���6#�|z�b�!�'FA�B���Ғ�ۘɎ1��E���x=�D���%�
]~��Q��_{֟ח�
(���і!S1y@���1Y��@8���
����w��o���	�D,��je��ö́y�W���[�P���t<s��O	ɴ t�#NKȬ������^&�R������6���)���,_h�}�8�X�­����T\xd2��F+q�r�"���,�*fT��&�����j볫��Ǐ��>;���_Ttʿ�X�h��GD.��A"݌㚿� Do䮁������[#z@*T9QϠi[륾ZpWL\k��t���2�̳����Zn�ָZ�~�y;S )Xlh1�"]�g�bL�y���l�j�^�F�PRC�Z��:��cd�㼠S�:�F�/I;��m(���B��:� k�)�w�`�}�٬v+�!�t��IFP����R&t �*�J�&��bgÇ,$$D{�l�p�2΁b�n�C����K�HB��F��)�1@U�H2x�*'�����M�0q	.�4V�^W�o��7��1�6���q�/��Խ���Ď��|I�c�'c���Sn�ߡ�j��C��ڔs�6�W��%K�dS�"N�� ���+�݅�����ɲ���s�:B#�)��Md�׉�%|e�l���_���A�2z� �>�ط�%{�_;�{ְ�ا=�(����ᔊar�A��GǛ�%Jx(��aua?[.x�ǈ?ڭ�ځ�X�֙��6@݌�%-���Vŷn\[,�����w��z�K��G�f�]����ؼ�w����p�q��M5��?�?��I��FX�PW>@��v/"�[kS�%��"�xe�/+����jO�/�r(��7AGJ�
���!qJA�c|��p1<��N�(O!w�y̔T1󂣈:V^���UBw/��N����4�=�	]����˺��8�T#�SX�p����s	_�>�l�3[3R?�i���Q�b�kN���f-]�]� HK&��'B*���O����p��RcCs;w6η�z��?���c�p�o�ؘ,oKBL/��Ʌ�����UL^|��]T�/1���.�J"}�R��NŔ�Xu��,)���#��_,�WK>K�'�;o\�W��azC���	yD�l��~p�^���,E�9
W3$o�9*�Êz��9�]A���d�u7�հ(@��:�d;b��.3h/�x`���?QTk�)�k��!�h�
Ғ���@��
=�\�R:�;9�7��X��Z.�ݦ��v�`�@r���̏��{`E�5�K�V�M�6?~��'�d�1X|�_�r�%�x���^L���\�s��n�S��"n�n�:=��T�������W���L����}-3g͔�4�/�&(�{eU&e�"��K�ab���m����qt�p��v;&<�;)�1 c�Q؂ؽ���~)����XXd{�X�Y_sV�g���� "�P��C�ǎ�z�����i�72xO\q o���g豫��`dq��A7�dv��O��;��I�l[pd�Gy�6��1q�a$��ќ����i�l	�`$��%cꍿa��m6���`;G�^s�}U�����|�|0\�<�C�)(�;uO���"UGD�<K$�:t�M,W����1�7�z$��r�-`�!���K��2˸��&!�S�'��0��)"�ùY�	��S����L���E���K��� �y�<��Զ�z��4��"{���&"zK.l��A�ɥ0�J� ���(W��V�z�8��6�����3M��9������!���D3�`W{�!��q�N*��ҋ��x=߱���;̧h�?8jh�x�k����1e��s>F�}���{1 �D�l�S;�.�,���AfAk6Ka���`�7�e��H�j�_�P̔�p�՜�7�ƌ�ʒ�7�Fs%�;�%=0v0iM�
��%q��W�h������x�v����'��1+I�Cm�<2�����m7����8�r����m�\V�˛���܎E>ۑ�m�h�p�-��X������hKAv>��G��<)R��1�`�[s��Y�{��BVo�(�����g`�a�?R4��O�Qt><G�S=:�� ��\��p:m��%c�����8���>�(Jg92��,���=� �3��R&¶��[��#�z�6�^�z�I9��m�im�Ǌ���f\J�$t�B��\'�����C��w�>ײ�,��Tc��í�̌a�L����;�pe��W2�B���b1��/Ċ�`ѓ��=+����������0$�!��L�_�9]5t/�|���M��!�FG� @��%KUa3Dߗ�����΂�D��j���v,�H��)�4������CKA$75k�y���_^��"�ލ`+�U��s�m��w�������� a ����6�����A�
���+��R/߭Rzoڝ2��|�cz�g9�ؽ�y�X׈]@�0P�ǳo�뫑�̻�o�r��sPb:[J�g�"��w�:�KP�
0k��y����ۘ�c�%*}��uт����w��|V��R&�d�\#��oe �v�7��k���Y
��|p� ���(���t�;���xo@�ۛ�o�% � ��"��*����9�g&DI{�T�"9��K�+��F$�������I�3d��������/Iҙh�: ��y��P��qY���m��LiA�sb=�䯉��y3�4�� �n�>!i��9G.��vH��߇�v ͺ!��%py�b����rTXY���`��޻]����sE�o*\H;����ۿ�<��{E���#p7RNw�lC؊���>�����j�h�ϭ�ɚ���*�y���X��xD�k��V�D<���\I
��)�{�=[/��0":��*x�Tx{�d_��	e�����s�Gj0c] �Ľ��H��Q�w�]/Gc��8�G-�S�z��Y8�����շ���(׃�Ym*��<&{]����lj���FH��H!�k����O5���W:�a>��+�UF��I�v���X��y�x�¶�Bzg��|��Ƅ�!���Z��nm,,��U�{[�WQ�Y�=�W[W;X"^7�?]6�.�ςԾ�R�Լ�QX����iM�~T_������xz���{�S9��Tn�����I8?Ъ���:�6�L��q�����O��]�f]����FI���Eű��,�D^�"�Jr�
�*�L�l`q�q8޿�Q�/w�^���m���W��&.��;q�T1y�]M��;��kx!&�_fu���'�G����5�?�|rh��$�A沁g�<�r�;�M��6P.WHկs�+ ��+d���33
Xs�I�t�G������lR�jz�^]{"�S��Z �U���Є��t�9Go��;(�pt�#��^o��ި�xN�p/1��~?��p�����/b�+��K,s2�1�d/B�J�ǌQ��\PM��}&~���i"|v9�M�i�צhv�)�_5n<m��S�є������
�4 �H(���4LG僔"T�\W���xx2���2��% @>N%��{�\X� M�z4S�3:p����ـw��У|��3�L|�8w�.��l�./غ���*c���"��V��hg6�>$��gy�"����:`D���wHLs��&�gLGm�P+А�w�������5%�`	9<���2�r/H�S�`���DC*Z#��Dݠ�Iz��D�%3?�����U��X��҅��X+�^tϿy�����92� ��iR�vO-MSs~o��f��4ݛI��>�m {��Q(Y�l�|��1t,�o�ڦ{��d�3e�[�G�t3Ύ�,��P���}J1gG�r�jF%|^x���2�f�E��(�B\�M=�^'$����9�Ƨ�W4��V�����;�х�4"���6�a����z��U ����Ґ̨xt�ޘ�����bN��K�Wg>o��;��l��\*�5(?���U�H�0u?u�R�qذfT$98f�b��VQ������l���wc����i�l-�J�=L/;���;{�o 'nr-�!� �f	��⢪K��uYP.��X���/8F��v�CYe�#&9�";XV!5�����pL���HW*�ME/J)$���G5�]�RI6WNs�y�v������Ȏ��.�Y��sr�e4ώŝ&�����aD�xk�N�Z���g\D��k�^ ���	�;��_�fB=��L>�#���5h~����j��"��+W�d= ^�KmS�?�Mp�i�17׳�5���j�HG�"��E�����>�?�4�z_����-� =���!4�� .b Hx��&ѽ9W�lW��uSc�nR(	��蓛q�W����ï;0���ͫ�Q���6�n�b>��CN�-���J`HMj-n�ɗ���{;Vwn�:wcg�bȖ�9 �>�5v{��8�r+))��%����[=�;�&�z���2Qe�����T
Q�{��k�2���>>�� �y�Q����Og 沼���r"`���(��K��z^�S�@�s�vr!�uR�]#�^|��H�<f]&�)�+���*���:�O4�R_�?�_І��Ŭ����AD���L/S�WG��ao�����W���]��$�0�W���`��	�߷;��(�~���D�i~�K���N�����`9�������k�]��h�eRր@�J�2�fuH(���XN��_j�����a�i��'����Wb0�H\�q����sm��Op��Dv������|�t�LC�F��+ߖ�l�/�2�>߅��B�E�.}�oK
hsP�1�⑟1����%��븚Q�weثj,�ؽ������G>BG�#%f%�Y�}�Zn�^7���4:�.BjP6�+1�|���տ���m�#Vo�56���%�$"�Tx
�[��B��b���*t�e�F ��o�h�Z�q�L<�I����.��>�@�ܻ�ճ#�=�8m�oβ}�����Co����D� �q��*���1e�Hӗekt�j{��1��On e��a����s;>��	?a�x�]�JN�N��E���S�������7� �XY#gwS�'褭����@��E�7� J��l�w�ź�3�M[y��U'�U�U]"D����[�� XK4z�T�ҦK���4�g���:��6j���f�jy��j�q/�{���� �}.�����u ��w\�����BL7��o=F1قփ�F�I6�o��X�+ p�܁��
�yyhx�1u�^��ׁ���.'ߚ�p�>)���#Bۤ������S�x�veE`DU�!̈́Gj�j��B"�LlD�f$2��\�=ƗS5(��o���@�9�a�?�������铣%�Ѫ��6��r�.�5${�턔^��F9������̱O��^O�sS�� �1���6�"��EAΎ3�S��yJ��<�%���ο�}�����Eƞ��}���$�|He�Dt����~�/�����1�Mcq[�zn�`r 3h�'�"L��׊P�E���	q4���U�>���T�9 ~�ؔF�R�S<H���S?l�z}��,�#6�xux�k.�>B�ϫ�VB�
�ϩ���ya���3򁏧���q}���tï�g�)��S#��������]S�͍!A#�g騍Eg袱��CnVm2�/���4E��rZ�`"Հ�����:V��HS`@��_O�������ݬƤ�>�,�O5):�d�p���8���T��)ᴘ���I#�!��r�$m`Ekt�#�\=�<����A�Uʚ{X!�m��s��c]�nk	�rCR�#���N'4�����2�v�����d�AP�9ua�	0^�X%N �]�d���ַ�y��M-x�*
�xS���LMQ4b ��ɖ�4Ea���(�@���{[�cx��H�5xލs6(o��R�k�:x����:�X4��tf���{���>1�|�	�f�?��%�ڧ� s��&TA��A�M���� }g&�ɴ#9
���*[R&U^�N��d�-!}x't��?)�`��݆��o�>�-��@� �s���������x���	X?F�q=���v΍l�9��t���W��H�k国h�d|�=	2Z�/��8��{a�=SX��Ϥ�4���_	%�I���qҙ�F������{����ڒ
:?<A��߀�vԷ�ē=)ywu�s�8�{O�S�J+Я�	�]2���%�C���w�V�-DuO���Y������w	gW/"T�a����m^  ���*f��(��&�y���tȑV:@w�f
`=&�Rp�_$��M���HX�K0<�H|�i?�_����`�	�W� �w<���Fjp��B���6��Dz��o�vI�Ù��S,C��:�ܳ��^w��+��B�����E��g�8�vF�vb�7~!�{+etn�,?���=y�Ѵֱ����Ls�p�6���W=�s�����Һ�!���ޗ�:��O/%��ϐR��f{{���L!+�)l�������nJ��7@t�+�U�����3�rh|�`A���Қ���l8z:O�. tF����wg��'�q+�N��:W�l/ϟ���E[���1UN\a�2J�(�Zh�J�d/��0�D����b��ÿ��b�@st�b���dW�<L8En���dR8�	�FEw_^/�u���$���(g��=��5]�O�	&���[���l�&R�փ8��/��H��J�ۦ/��b�����i[u����.�֊&��%:Y���Ea��~�/���}�A�!�4g�XI��/CNb���\ηt����=�s����D�6<��e}MD��W��BK#���K�{�止�{��Q"����|���v��̔��`�T���i�����x��Yy�/waҪ�C��}��ԛ#<�,U%���&h��`�Ƭ0�V���t�3&�R��zZ�x�;�Ae�4t΃S�_�+ٌ�L�n�Mq�M�'d�1h{1�������V�B:K&��!F1�،��$f����O?W;'�H�Z]�ٙ� i���S嫞Ս�d=���.����� �QBJ�~�7s��鸋1�����b=��G��q)�`���?�yDP���R�����H�O��������J^�\;WH���8 �A�j!�􆷨�ki�_�F�BQ�z�\q�$�TΉ���6�?�j��)��V��g�$iw?L���1�BЋ�Fk��u@��;��?��,�'�ć���bܛ�$kr�?�s�Ǎ�
����٦���_6���9O�/=I�@����:��3H���O�
�wЁK�0�d�"�@}���<��1�^�0�*�����Ns�ն���`��路R�t�w����&`��5�4!$Z��8Vfi�l�ý��)	�"�q�� #�G!u��Mw�#��'�S�E�I�1s��QϞİIֶ%Cl�L$���?u~�,��Α�N�"ړ��S\��F`1�����?�#���G㪖Z����g�Zb�=]�~�1��C����l�y3W'X�m��[�)7�<�N�
�7�FG�f�v 5�����`u@�Ko��v��$	8D�����y���#�B��������)s$yC��Q2��sS�5���+0<���]T&�b?�ĄUwн�s�-<���h񚉲�E�l��jIw�W7ӦC7��ʃ&^E���Ff�J 
Z�!��O�#}GS���M���-�V����X�u�hˎ^����3��W[�㏬Eg6`��d_�ȰI<Ź)��G��N���=���Ŧޑf�i���ܙ�����)eܸ����ܺ�U�����Β �r���!=d"i)�a$�Y^c�;1��;����@�Q�M
d}��b)��<������-HS���"4m����g�K�U�����h�K����2‹ �h�&��OzJ��:�Gi�e��{nv����)�^f?��A�jL��0�����vl(A�\�)�W�~Ng�rJ�y�Z�7_�<6�j��_��Ԡt�����ߑv�
��6g��M�v�he�����G���#n��w>š��*!�/�;ن����f�U|�!X�oT�+y�v�����
I�QH�D���Ko��嵣�5�e�|���\��hG4�Y�$$���<�ۡU-mi�w,޳n���`��FcԷdҖF�6�o��#)[�,
��g��+0��1������|�R7)q$��n
��D5��QvQ�ǟ�0x�)��8��/n�5�7๠����T���p?�~/�NT���@t/�?-��'� 5�53���J��"�����!v��3�V?��{��\��M��V����If��y{��)A�r!��#k����]��$�m��U�b�i�_s��n��Xtۄ��D���0�}��Ч�1����&�̣Oa�R��O�<.f]��nu�u6I��;��u �@[�*�7�na�]#�`��X���ȳ��r�N���� [2k�*��EHi��ߤWSZ<�z���#�aQ;���A�s��z>~z΅͗����M�C�����!�xꦍyVx��꣊��D;`lc�����:y̸�Ĳ�c/7
��57ĬaƵ{	�ŹQ��dA�i!2B�6�]l��k�zQ�?D��1��G`�Q\�=<q��}�*&��cR~tn)�����`����4 X�ٗ�PP����wF[p4�A/71���O��	*ށ���t��J5PlA%�#��:a�:��*�;#Xs���0@�i�zb3�5��|1�Ŋ�5@w:K��2����
o�ڍ,ԇ@���.�dpl�����dC��Q����X�L���,ק��ҹ0�=�(�	�9;�>����uGk�xR�G�ՓflB	�Ws�hВ�� Ǐ��M��\�@���U�Q���wx"z��/��L��ū��b��hd���0�UL@!�� R,�a �R�i�W�D��g/�ͷ��{Iڨi�B�}?��9�����Ni�젛7>-�o�D��dݛ;c��9����Ԙ�3z��P^Eǚǚ���̡������a1�_�G� H� c�DO-�OƊ�ڡ~����UT��XO�H�#6�j���ʢt�����Т.�u������}��<�fT7D� �{���䤕���a�&�L�����iv���s�&|e;���ɢ������^��.���W[�y[� �њ���1����{q3"��h�����|c!��c�{�ov�5�갃���G��ܞ�M/x�xԾ�dSϳI�5��(�#$k4��&di-����BR	����XC�ъ�ޯ�{D#}��x���bD�a�n��<;d��\��A�(Y�����5��º.�שu-�ɤ����pB1�xe/wX�t����6�:�Cv(��_L��lN!C�� 2;W[&;}��]�`I�R�(]�æ��(�L{!����˥��q����d�p@9'ݾ��b>D�e���>��z�l+ٽQ����=QJ�A�SU�'0��*��1�}��u���h(�LH�ҝ��dğ ����&����,h���Ss���w&8���=w ��s3|Mp��V�D�H�~/�� k�v���7�W��a�] tՂ��#އ��V*�sI�J/�oߦ�����]밻�Z���ū���N�$B�PK�!�,�ù���X�ё9���1#��~L�P�>pk=q64�&��I��z����drh=*�T�\�Cw��&D�\{!�k����*����b�F�8_��)���5	y��lXo��r��`��@��+�@T�ܙ]L+�1�"2��lt� ���c�z�ճ@�EN*<�ܓ��3�m�۱�Y��&��y�)zۘ�#bD��j}��z���ʃ��@	�1N�hW��UR�]�M�DW��T�,�𶺨#q9�Ҳ�ew�%�1��R;��L��"�ot.R]�bΚz,�j�D�����j
(�<�P�d&u�Ȏ��is���S�&��s']����_�]]eϪ�'ZD�Y��e�dDo~��/d[��f�y��*Ix�����q��|v��5M>�M2Y�e����&�ag�j�39��{��U*ڐ���D�>.���}y/Z�Mi�M�'ev��m� ����j39s֭.[��mgMh�t�$Q�~T�&�o���!fT|/I�����n���C�����a�RC���#z�,�f��2���FMB�-(PC@�`�b;�Iy��6���)� �c��H�����Y(��`�Z��*_J�n>̦æ�["����)�. �#�\����\��y��T"��b�DűU�u��זXA�d�f���Z�?�<��f��H��ON����Z	����cv� ��^���A�R"<�q��/���(H�~��V�/RuIj��!�Ȉ�O¸��/���a�j������c���̅my��*�0�u~ZT�O��d����v�mV�=������謟����Ld���22�@DX�|!����#�7�l#j���ɰ���*:��g��{>��a�в��Q�	ťpa�֡�x�������@��g�l��!�����=���.���6rI(t�ٶ�pa�M"8��=�u,T�?��Q�l��,�r*��a$�0�DD��z�;@?���j��޶�u%��"䬇���8�&���=�����E�X���q��tQ�U��8������0�:�E�[Dr?��G_X��ٿ�8K��EtV&(�jvf��6�飘{�!Kn%��h�\�)3-DćM��㌡� �8����]�㌫�FY���A�yO���������_�O�(�j_#f��2W���p���j&�u��� �&���t�N�Nc��Xd�U�.�l��C�Cw�����vrIw�]�\�z%�}ԇq�B ��]�Ȭ i��+�՞,��$�B`TV��y�d��3am���s�:"�呱dZ���aEP8LMc5�,v��V�����;6�mn���sZ^�+)4|9���L��b�i�~ԹJ���2t/]�eb��A��:�<WK#��� �?�w�HI��	��o85R�iʟ��:��bŧu(�����j�MM�� �� \{�D,
�HH�1�&���B"��Y}|���צuuyОX�<��q��J����]����g"����hV�M6�dQ�n�}ǰ�[7�����Y\��nˠ?ȴXу����p��7&�@"?��YM�#g��������9�+j�'	���.϶Q&��D;���o��������Q"��W"{�{K}D� }&G4v��j5T����S� ��Ff�[� ��i�,�&㢍��?��C�[,������{�lg491em|�e��2�/�lh��U����q[) qw�9qő��E�y�ǐ=��Lt6x�a�r��Y����۶�]��IA�ƞ-�Q�w^{���Tg����z.[���t�H��f�c�/�yP3f9/I���Q��O2Ȝ�_�)��>�Z��(�lǷ1����*�hD'	���j6�脇�TI1A���F��ʛxt����/M!�B�͵����b��(�"Nތ
;♶?O������}�-@�H�V�2a��T�<��kw��jB�D!�'61�$�3�Û7��@t���2�%��n35��y�$�E��N|<���aѶ�4,�{�ܪ�<��劖�ž=��`tPj��� ��ɤ�Mk�B~�2�8j�������^7a��U��	6�����μW�lڰÒӚ+Q�N,?1���3:���'�\�A��Ͱ`ߴw��Y�,����7�{�*�o/��ˊ�f��E�=	*��:�F(��q91�xt`w����pꎀ��9���oG��J��^�MJ}�w\;��U�7E�ֶ�gb������!�Ƃ���e�:���R�1>�s��A�+��"�V-+?��`�(�"\�5����!A���hF��$^~b��N+�Dz�b���k`�[N1�	q���b<���S��F��#����W�a�n�� �8��W�or���
�!��<h|m�
hd�����D�uj8~aOAn�eV�Я����
����Rb�p�e"BN��+�i��AyV)̵I'���<�p�cn���[Mc��I9 7��2x�K1�U�W^�Wة��(;Ə�@�b�.��JZ��5�T=(ٽ__!%�j�x ��2��L}켹���_�����d�!U�-;�+1��$P6 �6�"?�ű�9��]��ߛ�h^$|�0�y�vy�W�멏����͌����E�8��m�o2l=����GV#�a�nz�����m�k5��M�Aͭ�X��ֵ�)y֞�C��í=��f|yg�?K�N^�ǐ�X`�13�m��F�Ǌg`\	��^w��>j�t�!Y�4�:ɲ������<꒠�9����݄�z���k�G��K��C�M��W1tl�Jϱw>�)�8�P!�c�L�i���	�D!ms��\p��b���݋nm�Xvw(���K/�|�si���c�����"���ʶ[��.֘a��lL^B2F�*��/`��45^�f�tk�ݖ,���<����83��$�P~���Q��h�<�X��&���3f��ԧ���A���`&A#�?��թ�H����]~C̼F�g��m��H�tB}/�Co���.hgI<��X/œ �˅/�������K{�O���t@��,���z����+5�Z5�����y����yF#�:�<d�X��j�\�Ʋe�]�\�"�����W��[�ñ��f�sy�GaGTb��h7�iQ�@�̈����L�}��~E{�+~%��J���I2,?�SqG�mɬD�\�ˡ��D��>)R��� ���3���q��_�a#�ȧ"�{&Q��"dV��1���L#'%g I�K� "��L�$$�yW]�J�n<GmY>ZQ���g����m��v:����F���%'@�*@ޣY g;��Bn$�<P�Nbl#Ĝ8j�T꓇v���ܜ`�L��'��Ct�}27Z��!���23C�S<��>3��� K���ѻO�O��~������Z�^���)`�݃�Jȸ��BmO��x��4���Fo�/��$"dC�]�Vu�ρ�>���XT�����)�M��6�T����Ж�9��e�'��띷'���I�k�"..H9��Ml�x�� 傃�q����%Qx�����3O���V�����@<ɻ&���m )�r�5��6�f��xsW~ҧ-���eL㛣�*m�L�m�̠k�Є�O�KZ��2�)_��K�Q�%�b���	�)�Eܪ\�{���b��)g�����D�F�c�]����~��٥����4�$c�f�&�BۉS�l�r�ڀ���9�-����:(�.���q٭kA�I�3���R2�m���:�͍�i�wH��_zp��9~aZg@�F}�5@l#sR�c<8��P-j���S�،	�1c,�"k$`"��+�,HU�
 �Ʊ_P��$��טQ@D hl�č�!�������dTZɵ����Y�Z��K�9��w��M�����Mjį󯜏��al���G�ҩ*a�U�Z�Q��X
�r�i��]>�S?�ʂ�,��L�R������O��;���	*#�~��a�0?H�����_�����a:eo1I��!��0���Lsn���[|t�`mw]��!�}�U����3��>�iH��r�|�g|��u�j�R��v�������vƎ��b�<k/�B{gn/z�g6D%Ko bI�M�L�#�	�3Ԣ�o�D{�R����hC�c��Dnu�[Cu�L�}4Uh3,��uCR�u}��u��~�-Ed��*�����Q:z�>���Ժ����Rk��y�4�E/o�}B+`��@�5�B�8\���D�gJ)f��1q�=���Kzx��3��M�l����_#�����5e��&����N��R�M�� [*|w_"�UcX����ĆsX~Sbdy��6k|+'_;-�ؗ��`�_zv7&j�N��{�*�0���E3��.���(VW��B��J�!2��F��.��/�R<f��Wr�a߃rsyԢ:��l�a���_����
�?�]8��]��W���3�W�=������M� gل��3͑S$��0
����T�[d!�:�#�-]C�0�q�)��]� ���k�y�6�2�@���N��[yAl!�4ʕxP��S���������q�X�zh��>^��&�.��L�䪹��b#�[��Y���.,���ߚo#�,u�-��8�j3MU�Orb}4�h��L}�e��zg2�Jɨw{#=�]��Rr})�P�Y�!Y�r���H!_��^y�Sj����y:ӭ��*^ȴ7��H}�σ�H�
E�VJ���"@9�:���N
���6������z���%2� �ҋ䰼��Ώ�C*-�'^.�MDc���m�6h�  ����V�pX�g�	�a2+U�R!�9~bG�3]6�S��_���a;c� �=�t|Y�����C�%�Df�fM��J�Z�R.�ɫx�60����lyO(*KX�$� u���h_�N&�k�R��Sm�Ւ=ZO9��`k�� [���t��=��_j����*��5�5�<��H�)��ƃ�mkw�����-���m�����$���GgG�5�����eK+���9,d/�m�������P�J�+����,v/-a/J�8v)l� <2�='���c��F��8L��J!(̊���_t��dˑts�ژ���cj3�0�H�-zՖ�P6`ci߻�����gO�|�ۓ�}����������3�$݀W3S=M/N���c�c��n4��L��� ��C��E�r���N�Q��e�8���F�B��Ƴ�6�S��
�x�^j��ͅ`H�k݀��U~T}ڗل��*�r�\OR�-�"0Ve��-�;s���K.�U�֕��˟�Bn�y�J3&�U�K��
��8���kn2O�e�EC-�L&���>���ir�.��:���>-�&9Ы՟�Y���ȕtD_�5I�N$&�v՜���uN��C�R�\�"���^"��`@E�x3�R��18�+�`_����ጉ�Y��/E�r>_C���50���H4���4e�$�ni\ҫ�_w:�5���A��j/�<
C�a!�.k�(�D{.�89W*R=�%9����fL*��E���G�K	_����Q+��(��8lH/�g��1˲;�R�Ӑ�5�_����vny[��Ӏ��pUr�
X�\%u	�(5%�S˪�Y��.����#�����YF7ȬhS*��Cgߏ�,�^�%���U��w����i5R]&*�v��׽|�$�~j��:*�x���X�I������=}+g���P�n�R_͢���$uOX��v���6���anT�<ٷ����mY���Et9[�q�<g@�|?�t���gP���H9>���� §y�v@0�it��B�q��(���4��k[���i��;��WNP<����|>	�V�X���v�%VY1�0�Zw����/o�ڴ��1<;��y܄vo*̐�C�'S��X���o���>����z
/��gH�CF�D��Ũ&���R��[x�E_6��R? �f���ǀBt�ٚ�=�W��f H��`M�D��9O�?Aef����A��%�ޅ��h��y�M%�� ���p�d��~Jݖ�V	B Ю��4�J#@�	��R6&���pV�g�F�K��C��i~kQ"@S�Ћ.A���e�C�dΘ�4t�yr�+cz��z'��R.���U�JDOjܨz�1�>�7,��"�r�mJ����	����_�݃_&C�=&�S�Q43�pTy���(M�d0����^���
��?4ָ̃��%IX�ⶋn���;9-?�%5D�*l�m�
�uP�LhK�=�b�!ti���yIP�1ֺB{~.E�΂�4g �4����8��/%�,�R�83������#�.!ۻ�4��^���6Ly����)[8�$m��I�u�YQ�D�i�Y�ez���j�C��C׏�3�#�`��4ӝ�X��%"�����˵1�s����G�k�����_�bR%<�nZ�a��*=
i�L]��u[�"��`�|�$��/�}y�y6��� �n_6x��1���u=�x[��jb��\\���;D��U?ΑU�5�������@�ǴF��J3��g۷>�,�ݨ���g1�P����4������_I�׽�[���4o`.��P���h~d�>�hN�r[/ܔ�&��AO�mU��ǵ-��ڨe޿���C���UQ���Oc0��q�
KG�mqe�K�N��R��Ҋ��DR�4E�	n�s�˛\^B��w�BO�*\�N��>b����x4��e�u�[�/H\Slr���U@�����	m%���dv�;�n9��7
ͪX_m�a��|���R%��:�ðr=�`Kxf�A����YG�������=�X�N/@�ڿ8"h��?Q!97���dM����\tq�҅�ǭ����B�XM6K�Fl_�E��L�qHui�h5459"�����X�y�p9�R���ɂ��R��a�޶�
"3�n<b+��{Q�B���X��%�C�gP�?27�[ܻ@kv��;�d�#�Z�<���q3��4$P�9�B�v֪� 1C^k9��/X>�־&�N=�[!Ǭx�x�����<��՗��?TÔ'1�2�uЇ�&2�k��C��U�/'.�* ��؟ԭ�����O�����P�'*�9�&b�>�H�	���^���M�2/�6�)g����-8�G!y/��dӕ�5׼/'[��]���sJ��i�,�I7S�QY�?(Y��*���?g4�������%:g���P�RDJ��������I���9\��ԯ~���g�T��^�fp&��͏�0��:��(��SNTm%�E��-�t���\x.iv�p�ϫ
pF�͠t�1����|m3*`�MZa��i�}��D��a�}����"���oy0~���'�!D�m��{��~��9�5no������d�P���&���@�
W����ky穻eӅ�І�7x�L�*<�����bY䴐��^����!��^�ݴ��U���m�Y!q�I	�N=����<z�N�����O	h����Mh�TyF�"���h��(O#�*��D���g���������&��m�'LB�cL͈�R�1�dbȈ�{��5�v(y�2�]��p�?T�0�[k���S�^1��E�;hD3쏷�m�n�����Tr)l8W.$ s�ڱ���2U��ѣXҳȃJ\"N�]N���5`�M�N[��D/�|J�����_k�Ċ��� �y�ХUC

�DY�&��!�$����;�6jYG�=��xl���hS�9�����m0�L�\|���]�&�O������x !z%��?����q~fV6����U�����X�-���xo��0AJN�L8����ݳB԰򀯧�Q��;�����0�kx���A�[�3s��H��]�B�C{�A�yZ�&Y@��7(E$��(	X���������Y��_IJ9��ؾ��?.���*�;�vw4P�>���٢��FÅB���0;=(�K��& �2�gj��
ߝO
[�c�<RW���Ю�D,<��nH���+���S�G�$��!H���"�v���D���u����gh,�uk��6���Ȋ�jW�6�.!;���]��T�]�Sy/�O�`���"k�on���z�q�I��{-�� [G������[�h����|�[~?x=��l�W�q �̄��Fe^�t�����&G!�E�� 	�����p�1�&�G���{�7���S)�p�Kc���/�i"|f�b� x�< �������`K	�uز�֖�-l`&)Z����A����M��L6_�)�-n$���4�)�D�d̬�\�MKu���"Z�+!k�bZE�"���X���*7:���D���4v�B�U��=�@&2��Ճ�ӊ
���I��+H��/��.�aRF�#�}�˧#�8�Ť�{�T�6�B�}$m�U�k��"p��ou��,�pq?F7&r�s
v���k3��e���D��.9י��f3��?��
S�<�`���Ѝ1������;�m�Lk�Z����v�M5mo�<�i:7ZWJ�m&��h�@X;��^^i9m��Ʊipk��?Q���qP�L������PKu}j��g�}�(�e�swa���0ف�aA~�&D��u�С���E(��n,CXY�d@�����J1^MVlǻ�H<�JkLP�r�?\B,	�5�+آ��5,U� ���(�����Y�8�9Po�sb^����9=��fF�H/���%o���%9��m(��_�i�3��N�=�I�ko�K�0-�&w~r���T��Z��V�� qc$���YT�����Um��bx[�Q��j蔴�$\���BUL>�?��e��Cz7�,�=����
W����M�E�*�&w�uLm���,v��?�TP�Db
�:��2�y=���^k���Vw}J�V	���-k���`5��:�0���� %3,��강5րd'�-���N�7�UHq�T��R��p.��g��mr�t`��	�F���1��bk�d'M�.�\v�5J����H+��}W��e��@ށCr�6O���XO�d!���猒�\fQ;�A�q��'��Ә���m�͠�s�s7@Z�ڎ����l�����Q���A�I�p��{NR�F%A(�.f���� ��0����M��`,R�����ڎq�.Y&�<�q����md���r��#�9��";��߂֪����K<B[�j�����_�rة,�L竜���Tw�p��۫�>����IP��0�A�P�y�p�!����YsR�o�1�gͷt�P5�7w�C�g@R�e )���$��ϒ�*GM��AޙG0�	���L6W ��� 0���yN�
��W��Mn��S(�uкĆ����5K�@"�����A�\��Cg��!%Z�sBيG1Dm���6/R�d������%��׏�ɡj��1H�x����!O5��}|C�f��'�'��n9��8e�i[~�D����p��J΃Md�O(e �6g�D6*g_�j�)%�*?0 ><�bKVt϶/���7E�/�'1�ݭtT�@1��G�hL�=��z�H�L���ښ�0�R�Z��ۃ�?�B��f�\��p��@�
���	\�\�a��8�x}U�BT�#`����m���B��Z�6�K=�0�^��w���
�!ģ�!Xn��b}��B�$�X�	����%�?���wL�f�c���yz"c��u%�s��;(�E�= `��r�8h�)%��/e�㥍!bڀ(�Ξ�;=qR2�Md%� F�W���7�e�4��X8ƒ����1Q�~���b�R�Kwa�CP�gD�S*�g�T�Ceg��D�l!P�~��&�1ag��8�6�����4y�(��Vγ`q�aY�#"_�B�Qpd��d(��V��m��w�O�)���5� -��#+lְ<1�}_�6�%�Q_3`���Ls~�q��8;SdK�A��&�FB6���Jq�FX�q��$�<<��� l>���A�}Ìe{�ދ��Ih�'�B�R�Q1�c~���s5�I	֑>��Ɗ�;"�R�A��j��KJ�Z�^�r &zLL����P��W	�l��nn�a������^�B>��96�+����kY ����2O*��z�W;Z�
��N�-���t���2Bj�&�]��4c�ʗi2f��aa�v�1��u�D�2zY׿�lk��SF��mUw�j43�p�)|��)
��'B��#�I ��,�+�7��#:�<N��k���|v{�wqM(,w�����J;&´����p���d��ӝ���$^�QxEy\�S��c�aN��;��J7�ϛ�
Ģs�/s�@�Y#�=�[5���JT=1$�%T<��LdZ�̵�A��^�@�\Js�3�$��H��׭�H�m�#�
@J��T����u�mgC���O�5�0�4y#�U���K8]�?���뮻z�޺���q��'�=��Z�{eڭh�?9���<�fo����#�3�Y��l
@��g�Tn@kS����)���F6�L}�����xK`�^k�G˒κ��a�DMߕ��Jf5�'�g)1�.����	����[?��	��M�O*t�V��.Y�m�g$RY�I:g]�)焘-���raj�G�'BV"hW~c5p7��sҟo��Ay�F�0��z0�j�++�|_�Ʒtr��i��P����g��i�T�D�$�@����xO ����n�;':l�L	7
t��U�@�!��*���'5��wju�3�=��[b���]^i3���S�{TrA���Ҡ�`��H���*z��@��"�a���c
W T����6�U�dɁS�#SA6���j����D�<|�U�)4tZ�*��>�D~�)>����3�1����uq���9u/�Lc�Y�ҿ��̘��_�Dd�
{C����PI�z�Qʶ�w ��&$u|�s�w��TEi0�9 �s�t�v��J_����p�#���yk��2(��5�~4�TAyQ�\T\�'�Ą���$���w�pV��p�/�3��`�~�&O����c��jR�??�|��w���`|�xs��>�<�c�ڴ#������@9rbt�y�̝�D)q�L��Gu���ƾ��c9�n���I�|Wp?3K�6�_��)S�*��հc�+�� $�����cP�;V@*kӆ(�?�6�L�R��R�V�T0*�s6�5S�5rW�^�����Lı�T�zǏ���dL�)��o�op�I	_]o{Ƀ����E�$��!W����<��۩yrI�[R*{��!0)�m*G�+d����K���*��u,��ݭ��nd�� d;D�*��L�D��c�^1�������O�P�4`�h���q�a���^ �s4������ ��ˢ��)��2�^!!��s��Z �ׁ������,���'ӦH%D&,(��1�9Q� GO}<��r{PT�l�@�H�a�"��p��>�<�<���tl�o�$��\�~}��@��~���;v���Lf�d�s�v�u���M\�RG+_+��8~�ZSA�}6���(4��ۊ�>��+C7���_Xg�{�e�w�	?'�~�*�bRO��6-<�ؕZh�UM�Y_���0U�ƕ%�Q
 ���A���_����E22_��'tn]S4q��1�Q4����iϋ�`?�چ�C�HYu�X��/E�t4`S��!������I��#��榔�Ɉ����+�1�~�Q8��Hy`�T
�z�RF��[$�����X�"6D�uc$�7��s|2�T>\AMt츘aŦ�情⼛1�R(���f�h�^����l�{�B8���������7M���ۗ����D:�iGVZ`K��Ŋ�t=Yg���v��cFvcVi^��M}P��N���l�t_W�Č:ܩ��J�9gH,��=��B�s1���7���氺,��(e2��?�W'�؊��V��T�� X���w.��d`���6�z$<jJ��0�U�;H��ZXt7͚"�\-cSPf�g<����1�oc�J�ѳZT6�����BLZr¾(�du�W��f@���r�]�2��'��(�R�c��M�u��U^YmuZ��~�^����{s67/��s �K����r��+]��E:��3(E�;A�V��b}iq&]nFǚШfg_�p8Q���Q��a��u?��ͤ�a@s��/RD |�<�x�C�~�ߋ���2_��K��텺�f>A�<�Ҹk�l��)��4Q�)����o��^��E��<��$���0ys}�]�薖U��!7�� �\i�&򤄆�1�KVZPc�6��ɪ.��~�HTo�<�ە��k��������Lo�v������I��yYS���Wɡk���&Wb&��L`Py���	������9�����%����xY�j~v�W̢KE��(���7��xԼf5����3�%�zNWMI{:�
tk��w,�)In�X�2�x�x%u�8�@&C��]x�H~���'���2���I�Z@ZbLdഈ��k�����sF��2�6�v�����w[�;<|�5�-�@2WQ#��Q���Xv�d��~ #7���˽kP���	��ϟ��+;��f�I�*7�f��W���*��v˙u*#� ѭ���) �ÈB�8�/�D����30�
m�}�9� �!�5�Z��˖P�6�^b|al�P(7������2�u3�jZ�ֻ2es���v2%���J��������^�C{���0O��S髤�������}����ET���C����,`!*�D�v&L���H	d�bJ��]fR�'mV�N��f�
j�-c	Hyd�v���l�`*c���� X���8L(�iQ'��KEc�)b���_�� 7#K��� mV�l��tH��6��
+�)y$m������R�'^ ���6t/��X��~��ޗ����+�4���L9�� ���+$�8�V���Pa�� �pC��^~��:[)<��;�
�L
��Zo5�5A�8�w�n��|�mf��prͧ+�)RW�E�	S\��-Gm�;�r�~������Z��=�j�m�`�R�-�k�����9���|u��F\��j{M�PCNv����Q�"��|/3%=m.4F��#4�+2�lq45!�*B�̽�ٞ�2$�	��d\���2�����>���H���O�ߎ����R������'��}�2�4�����I����-@R8 ˛�ME!Hu*�5��G�+�̷������<J���fR�X+~kAݻB���L�ˠ�Ei&�$����X�0���Pb������L� �My�M�ك��w0�����������1�G6�����`�ά����X��fL�&8A��0�:�$UqN��eB�@.�(l2�	V��O2E ��h+��:4�\X/ ����Y�w?xD��p֯
'��n�'_d�zg�Ђ	q��|��#��8n:f��� Y�fB��C�tN�k���2��h�%D���}�F�~�Q��K�d�;8=0~�!�M����}�[��72�_��E_���h��0d�SIQ^d�.Vwf<��~Y⚦�[���Cʂ=������&b)j�!E�m/S.�aa���	�#zu|��(d��66���yⅵV�|���?i�����!�U�7��^��C'#'>U����#3٥o{��cEލ���Cs�e��V�3�mxg*�~��A�Lt"rʧ��^Ʊ�1=��A��:���%�F�K��٠~:���/���m��Iԏ�)lң�0%�1im�2�0��<�����ܳE업�uQ�&t�ď���/����9��i,S��L݅.�1�.��nJ�v7�$&6�t{b�=w�PJh�Y�:!�u��u�Ŗ�k�ˠ�,Ŋ����2ߡO�Nd�_\R(U;G������2vw���a��gn���;�WH�17�_�� *�[���V�S���>��<��%c��Ŗѕ��1��VV=���{l'�b[z�{,�a.F���|)[��G������U O�y��mT��V�:����jf�s�O�Z���,�����W���%L������]w��)'~ ��-�as�'�$��F�uy{�~fN��|�>��C���$�a&z�H��8���Xy蒖na��b��%OT
��
�����xF��x���G3i�J�;����in��FKb�~���)[, ��,�ꇐ=�	�QQa��4&�Ś����)4�Y��_u9l�����@c�3L>����-����Y�HVݦ�(K��`��`�-�K�o��:sj ��h|AN��檄��r��-�$|hs�xz"��\_�r�X~�G�.}�(��EV̴�d��.ߨ�i�ǖ�ќ��a����e%�5��jװ�����Լ�6���P5M�E�G�|�T��_�������t��U]B�d?N&1�����;}*��R��2��+�k{���ɀI)����f���~kt�g ��Q�XZ����S2�zMz�C45%'�(�"l��3�r*ڥ��y3r� ��t�G"+���`f��j�$�Χ���Tc;��f9~4�g2��HF5�s<��6��d�)�{^��sM�S��U�y���@x�zl��z�$��``��c7#CE�Y9$#�ba�͡2��<2O��y�=���qX�K/c�����on%�f� Vw�O� l�)��( ������Z��
H�w��3� �>\�Wy�4W��Ewdz�=ڗ�Z:F����ci�)�J�j�ڌ��wBA����P8�S@c�3�ҷ�o�>hSI&�k� RE2���2�3�j�*\�<?�Ȕ�z��f�1۪�ȅ��ξ  2[pE�ttU��4�z����D�U�׺".�>�+BubNY����)��x��m���ΦYu�Á���)�@��@��$*h ����Dǝ�.�߬!0I@�����W*�Y�D��8}d>�^�{֝���4�� �6��J���6��9`Q��V�������´�E��#����׿���K��H�0���ߘ7;���ư�C�s�r� ��FEɼ����mFc�n���8Mڙ�m�tyU�l�)ݠ��J�,I�o�9�8#�#�_�8 ��U�}wݾ��z��eD9�[V-9F�H��_	_�����_�W�Ԕ��T�]��V� nZ\@e�>�]�W&�P�I+��X�i��Ps�F!*���_������gx�_@Sv��ݟ�:��� ��28�f����ӹu���j|�zf���Y�O����-� ���O�x���Y�N��W�\�� �Rg���B�U�R1�a��A�u����:[��V��άG��B�O�k���YK��߸I���ܶ�����;��`��6\�āT�2Q{�퀊F��9	��G\l�c���ߘ$s��\�Ndq_��L��,�	���#�X|v�w��� ������F�: �k�M@�0����h3WF����H�F���4?[I�N#HW��A�Vך.��¼��U�ZfG�f.�oFl�=tNj������C5�S5P�n��A�`���@�+���"�(d޵����e�"7[XMҳ{�#`�/��=�W� b�y��x��00��	���"N�U�<����(��R�'��rz���Eٶ��͐y�n$�<�(�T�=�����r�;�S�sL}e���q_k�dm�:`>��9�� (?h���)�0�*�0���j���&AK%:a��������WB�����9�?oü�1[�{�ݻ�1V��k���T��.���\�2H=k%F�����t����E7�|�2�Կ��&'��3��UQ�'H�Ƣ�� ��� *rH�0�s�$��d�����>��3hÊ�4���=)W�8���	0Ԡ�i��rAX#{�2��`�军���%�����zd�9�R9X�f����d�KIa
�zs��|��v��pk��bWQ}�� =]�������	7蝗.�"Q��#K�8g 9�RO���e�I�/�nn�rL��j�hb6Ѝ;0Qh�^��z�{&t���p��M�O@R��r�t�`�A�:}�Ƒ����j\e��)��*#�&����a7��ͯN�%��ؾ!��[b�����Μ��͡��/i@\V��|�3��f6� ��4�f��Jc����sgݬ�th^�FPv~��μ-����⽀�T�������>-��B[I�ن�KIQQ��U�n��&2B.�1�;�&���L]�vҁh
 �!��`���sI�vvW�M�9Ow�a�E)JO��\�(�ʵ��	_����1�e�f��a��qW�P;�^���.t?����W:Z��TC2���.���Q~�J��¦�LÙX�|USn�$D����8�{��b��x�}�?}���o��*�7r���H�T����u8af�����ӟ�K䢀F����Ts@WE陵��˯ZV0K��*�I��n��F�a3��b#U����i| e���\B �26��:9M�^����> �'��N���[G�@�\w�/8��b�1�ZB�yA<o�qPk���T��=SM����c>F�)�����pS0�����U�Lb
��M+r��J�ՖV�U���)�Z[YIr�M��"���8WJ�X�f;-~�:�Z]g�X�7g_d�a��*(�o ��א�D(?��s+Þ�й�O0�6�� �̈"�lH3�'`��c,K��0�Ԫ`v����P��b"%��ؿVq��m-y���e7z)G�u�=�3B,{��r��4��)ڋ�́�#S|�r3�?Jǆeg�iN��J�mrB�tOZ�c̈�
Z�[�7K���_ۏG(YZy֒��ī��~��)�Y�~�_O"�X��'�[���S��O�?a�-���QĞV�&t��߲N�7&ֆh���7h](�m��%�}��������LD�Ͼ�0y˯i�Ը��V���_�%$��T�~Ǡ���v�% U�I��k=�J���T�L �}�}Y'tCrA�3!��P��ƫ9/�d=v���
l�%LA9��,�a�!|��c�,0q��3��f� "d
Z��ה
��{Pq�mOD"%�*����̈́�e��+`�@�+w�j=��d�O��;�����r;-Tr�SR0��J�*g&pJ0p�~N�S��0B7Q,����?K��C��چ�5�ꚙ{<T�E��Hq[�H�Fw���dS RAjb��DZ�
�7��9�:V�5��/�B"�4��a?���@�w�]�MuQV����NR��K*I�B�A*:�b���]4���^��*�M?..=l��N"^�
���)�/>YW��1� ^�s�lU�926v��W�ʹT��tWO�Y_��тh�JTO�Dnם[t�T%[��Uӹ��Kb�lh�����*�������k��BNA� =J�� �D��:��a��+#���X�}ٲ���> +�1u�C�2���U7)��ܰ��sgc�g�P�<�3��ӷ�6�J�I/�!T��y����"<��Oag|'�Ha�.V�"ѣת�F�: �z��Y �C]6~p�i%
�)-R�L)��-: �9?�LsK�^��R��Z{�\����k,������5m��<��۬�?�c���>�7�c��u��DyQX���{��"x-���ACq�<cRs�:�W�zr��_�������t0y�m��ӽ��`���,�lo
�?-Ă�������l�a����
V{P��lW}ז?���P$��2��^7���l.^v�X�Q�4=A&]G��$�J���'.L�-�yfދ�?fλ����Y}h�j��f	�����ڌ��v�`"0h'�*Ҫ$��)���ۄ~o)���#��[M�x�:�q����b\��?�Zin����x�%~�?9N�+���WG��b���yw�b ͆�Uk��\��� ؅�ɪuT�9�&s��Ac�Ʈ;�v��Bx��|�><gy⣊2QxC	95��F�+�hP�u[��W���<�.m��P������C��e}����Or7Iu;���^�~���p̂烬�k�;<���#����h�oЋ�3�U=�E�.8Aq�ƾQuа:� ��)߉������i]m�S��|��GJ�z*��H
�4X�i7o8g7��>�-9mX�h�k�	�3�@��{ַ/\툂�~!̈�"�g~f6��v쉻^�@<Fs+]�۰;;Ɗ�XU�E���C�C�Y�~m><�n������ů�!b�j�1{�i�ו�mi�}�=�8]W�sG��r��.�'�� ����u𠏝���?&�q��j}N�T�G?�[n��(@,��J�.�G�y;�mH�.F@���FLU��̿%�|{������4�s�@_O����h�mC%�Ҋg���������h��m��6l����.w���7����TS���h� ��0�gO�����P�.]e��}'˂ Oj�KH��>	�fFJ�1/ A`D���b�d9ܫE�՘W-�HoxM�3	lj����G��@GiU���<�S�.�t)������m��BE�&�|�.݄����[FHdO�w �D�G�T�81��(�A��8E�a�E�d�D|,4�6������t���8\!(�ۇU9�z�����M��_�.N �إ��Bx@�����Qp�V[�w����XyFQڜv�#]�-~'��h �b������v䰥q�E�X^�ęTj
������gO�9� �7�"�uyP"#�[�����U�@�!�w�4!��3W���8� B�G�^��<���♲�h��`�f���ZC�SF�R�S��P�iMW���g#w�[��*�G=���=��x�f��*����UvY�a
N]�~�Nw�L (eŜgM�&�x(�pE�����ӄ�0=X�Q�a�;�`�\9��q�N=�|���������{J�����6�K�M��hu�Ӧ|ruc����9�&�VwЗ�/���U������g�T��[��&HkJб�����(�\�C 	J��\<��@���9j�Q��f1ւ���;,ع��9���+$+�M~�v���O�9>M|۰�f�(��_ޗ��J�Z�L�ص��/X:�[֍�q��_۔ �#�RމNJWr;kK���?^Eͨȳ&���B��S�=_�>�B���=2<hфo�럤A����#��x��>��y�}>�uQ���l��d0ә�h�Ï�J���� ��?�:jb p�Ts�����u����0P�(I������{�e:W\�tx��T��TAg���A�Cvʗ��96���6+j&f��X��#�)b95\�}n�9+$���ن_��ɋ�(�:���4 �Et�#���ܺ��뗈����^u�RaD�X��E���9;��>���n|�/�O;�NZ�M�)'��32{(#-�Fx�CRR ��~Ę݃.L�nk]�.$��rrp�t�j��}T�kL�+0�-4�.�_� ȅG�å#�����E�?��x�l�9�S��������o�E�t��[F���z����~8�t�qtd6Z���LR�$�/K:J�Ԃ��L .b�&t.���Gk�W~x_]	��P#�r�o��B�Dt�� 7�;|Zxc�mK����?��E��A�>���Ue>�[صͩ���0<���L **�����9 Ľ����C?��m�w)[$1B-�dl�?̝
�	�B��2���0h2��(�9�d+-gM���G����ʩ�_Z$)�8Z�N纇I���[��j�2*�}���	U����	yKN8M6!���iq���,f�N�+KA�%AX�k~�M�]Ԑ��i��gى��L�v��A���q���#�|D�
t�<9�W�ɘ�'�W����i�B*�����
N�:�t@�1#J䆝��ҙ�Lm덒-AJ�म ��s3���n�_���6Bl9Y��Q���ikEV;�X�)��I$��<����$R���k5��'�Y����]��	���5����!Q��(7y�����L>M!:!�y�Y">��H���v�����G㪧�\	gJ��MnW8���t�u�P}}Ϋ��_F��
�]I=ظ��ԇy���NA�����\me�;6����n\xbJ�����p&
ԑJd6��Fq������+M�����|��6���]���]���'���8��o���f��m��,�A�SAG�ZbR}��&�-]a���kt�Pu{�r�<�q���k9��X�E��7��h�gC�u(�!����g��p�?�)ܹE5^}�ᮣI?�&�^��GB���� �]��8������G�h��+d�X��T}p)S':�Z|��j�/q$��,'�O�NO�`Ie߮$��?-��0�|e��!N�AZ�UV����j��E|�K�?��i�u�y��p9<���M�Gpޟ����@��i���[I�.LoZ�9u)�#�V����^.P�!�K�t�Љf�>��e���}�h��Pe�*ϵ8V� ���n/FI��xc��@��l����6��rȲ�K�u��pׄ�����J���m�\�H�\|6E1�	�q!�1�Y=�+����>?>?��U[з�������>�tG}y����n���t�ȭ~U1�eѕ75�CF(|:���U��	����{�pr��ey��۶Gb�./d���K�>��g�)�Q���Kf�j�������R[J�/y���YEz�߄QO�A���B';��C���ĠY��_�<��K�պ~�v�H�]|�h:.�#��� F �.PX8��,%?g	�R�|~�����ks�O�؜X��>q��A[7��^'N���H����01�2�v\�`�;g�VrE�uYe�V \�'�ta��E�
�(��qB$�%'[㖶����5�����	����9��_90mВɕb�8���:�����u�f��3	�:�kS��\034N���11��- ����Ǿԉ�Q8M?yhu.�7����#d��zȑ��E׽�i��8�����{'er��q�)�2�f�
�w��`�Vb4�5���rl��ifsc�I��� �(b;�9�7f�i���H��n�x�{�n7/�K������fȵ�٤���ѷs��K�-I�/�<S�\=�����(l��&ϕ�G�u|sl)o���hս��`UL�2�l�`
��-rNV�ŕ�NX~|϶E?��D���#܃���!���@�x��j�=�^J���p����
+
�`�җ�[��DbҦ.(C^���B����ZhB��͝=��[�6�����+�VL,@�;����BSΫ���}8��IwA!��w���Ku�"���pS@��\j�P��r�넡��m�B�`7'���" �D��94��3񼑙�U�E)�`d�.�O�"�bjs�i�j�ZV���85��2B�0J�AYS��(�C�d9JE>�?�7�#_��0W���D�q���ͧ��y Bh�jr��^+XxL��-����t9��u���Hg7�U�k}�xd57V�"6��,O�Ѻ�:��A�gbIaXx�&g�;�qU�|�PF�$����ƶ��tz���.\+�Y�v�i�� 0>��\��y���K)B��j�!4;�6��&C���g�^E���<Y���G��;p*��Z��'�э�[xWy���ǂ�����B6�5�O�E���QYa�`e�ԗI< b�O����~��/�Ը\]�|U?��L�^9�6j�y$�?_��eo��5�H��m��u��-Ou��J.�����C����ak�:~0�^�.g��l�B�EoA��Y������4ـ�u<�rɪ=�D�%�OW�d��e���~(C���\���[�l4�r�U�@���9�yDJ�X�j���%3hQw�"�.*�����~�$�/�-��]ҁ�ψ^���M�%�3m>֪�{�8�y�\��˾��C�E'���&b]�;$�Q�b�!���A��t��&$����z����W�(���ޛ�l)n�8�h�纚�Ի���8;~�'�)������"��/%�l)e��})�~#�l���s��#�H`4�N�%܍XS�>�O[�%����,���B�O=T���B��e��,�����g
��<[	��uNVc�'Ѝ�·VEM��P��ۚe�k@�-����a��:�~b���>�����A�CB�F��d��¦/3~��5`���u���Z�޲����nڿ��]�"�������F qu �XE�^ :���7v�����o�q��-س'�h�t��69+�[��q���.���wN��`�u�+Կ}BA��D,_�JtP�K"jh����=��t�8��m�m�Е�ך���q ��D|��LϘ���p`G@�|ky	�ȴ��3���R���4�.G��J?{�o��l*���?#'F�˂\ON�p91�ә��%=c����Ǆ=�{@�>�k!�yD�􉵦�5��l��c�n`���<��J��`9pY^ϥހ_-%�|�b��q�i��*?����A"���,��˽�~�M���6�ߐ�F��d�l5/����#��U�o:�6��C����d`(��V�۲�����h�	V�7[R��9�22�J>włZ�M\S'ёū1���Tf��:>�N�&V���RȜaxN���q4�1T=Gp���f�s�0Âàl�e��8`9�O^�T�7�="�y������ �%����9^�p��}��:�t`tPu-b��'� �)�fB���$_g
�%q�5�� ��3�NƉJى��M������dSm&�˩���2o��z��BS�V㠔͂�^a�s%���O@�4QCA���2�Uˎo<6�x.�\��N|�S��=D�<gM-��PQaK�x��B�ז16�������(� f�L�Y[����1����n�(��>ź��o�N:�Wi���T�v�7�eZ��*�p;,�0%�!
#œ:j,䌃ۿkΣ^�"^Ӏ�"�H�-�tǾ*��L:}�9�1<m7WW	�ɦ��z���jt���������f�����������[Y�b���o�!������Q_�����t*������uΌk���2\5������D[* 8M�RѪ�k���,g&k����V��W��*��_x�8�{l�d�_ʎ�EeÌ��V�+��)ʎ1�����������sC��v�loܶ���b�v��j�PX���E"���O�X�h�$�QÙ���c71���Q���E�{"fF�MZ��)/��u�fԒz��:8����0�PZ2k����jy�i#�{^?{�Fܫ+�a*B	��9!oB*�����`)�{���er�ꔹW�m���Uf�m�jM�j o*om+�sYX;#l>%�#�/��W7Ji��C'S�,j�����ȭߔ�)�տ"�ƙ,x����B�o�h�]rJ�-:Ż��(�Dub|������V�&N�'WݘV����Ǎ��2X��B��q���љ����@�iQ1�|^�����B˺i7Z�t���'��li�U�	K3"8{���?cd�q���7d|ԝE	�������f�j�b{g`'��1���͡� w��B�'��aS(�ف����@�M����2���O)��0�OXDi���2�Z~]zNb@�|��<a�F��bTa������l4b��8��\����E��k�S��n�ja��a<DR���a"�,�Y����� m�����O��(-J�ӫ'�c�y�D�iY�_�����Z��������BB�;&�D��^1����~�@vYO!_���}	.�93�t����1�h��{�m�8�Z{���hs�����1`X�G萟��T�P�gFv�$,�Ł�4����|�)�r������e,���Nǩ��U�XH��b<X�X�-EٸH`J:6?�=S����y���d-�8�b֗����ޫ	�5�R:o����6�T�h�9F�� �/l����#8"�Uh�):��z��:!k(�u)#9�Q䈼́�ȁ��?���s�2�OG�[����~� �.����2�y���9��O��obފK<��/5꬯�z��܃���핁�γ��3�p1�V�H*���,8f��˨M�I�83h����aͩ��
Y�U~�f6�R�,��0��NⰬ�qo�3sP��E����5�6t����^EBKl���^zP�{��Y�J��6ؔ����?b$@myc�������Y`z�x�K��x��TBA��V�+.:��,�v��gC�,(R#u.&���z擧;���2n!k�t����W~/�sCfv7a�K"]���ƫ��i�ZS����%�e���7�j��=�s=��)zi�pQ���Z����wZ�>G2��Z���9A𴏵�P�b�)4({�*l��2���q��X�w����گ|�ǔ��n��fSdD��v?瞳���'��y �שa�:�y���#�b'���r8����u[�n�JzKM��B-���gZ�cq��h8�`ena�h��� 
^�{���
���M�M�$zOj)�{��O=��]��Nva�v4Pn3H��Gr�Q��y��O#���FN"B%���}�Hd!��5�j����c�̀�&��_�ؙ�P��&ֽbR&Ѐl����Ha�z��J�ƙ��@{[;���-	=!��E˵O�iW壷z�n'D���2��c�Ka���#��IVo��y,r�ml����CX6O����GزӖ�+?�r%�����Ƣ�������w���VǦ�X�-��:I� �s�J��#_��8Q���,lOOP,.��K������V�F���ip��	��p�[ij�!E<>�t�P�lN<��*e�R=�65&��x�9��}FǮ������]�9$��$�����Vbq�
�2VpY쉒m�??tFms�����[��f.U-��H� �
�+�Ii�0��/36��T�H�VI��晕͖���FxY���ϵ��Yȡ��J�LD4(�W�|g໘J�5��V��Y/�ϕ�OgR��oB���a�H�0�����w͸^մ�m�V5��%�c}�-L �Gqv@<�ٳ>E�Ą��`s	�"�eh�8
��Ҿ��|�����A�L>�Ѥ���I��`�a
Y���	���D�Σ�_��K����@Rm+\�s�Jb���-�����7zζK1��HXa$��-A�KO��]����h/��#<d�-������ c�s�ҥ,"��֙��ib��C$-�=�vKˬ�K �B��]���1���=f��1���g�!��oRMG&�O�kD�"��vQ��1�؋��H��[�<) ނ��=��2���p`�#)+�R$�SR����M��a0��c�7���=�,��4����8N9��ZqUU@Jv9:��Q����݈Cp,�pe *3+$�p`���k*�M7-.m���<O0�j#��)p�������e���`������0��[�Z�=�.��i[��J�&�I�K��������>"� ؀}�QÎ�G��	0u����s���4P>߄X���<n�]���f�S�u�?m���s�S���X]8T�]3�{���Y���c���<�rO�H҆�N_b�a��̬���;(��X���Q�&l�j�H5��|]�~������c�iL� Y48������n2���L~���g����t�pI�ԥ�6Ԑ�Z�qC���5c�2�I�3G�M���j8��k8G���6��X~�9*K�N`�ĊF��-����{m�|��C�{�G��Rs�g&��Md��@���O~��v,���Z\�po{��'M�	?�Ɔ<tmV-GV���!R����V��-ؑA�sF�YJΙC��*���:�ط3+`f2��MxDMWx�>�6�a���\����S4��ϋכ-�L�Ƙ�q�yx>��ok���e-�)��v�r�HhlS���=(-v
X����ݙ3o�k(cU� �R��?��e��	AX��\-g�0i���M-�b��k���lPQ۹2�7�ȢL�݂��(K��jl��
��?u��ٖ�6F#e���w�i��P ���6;�R_��v�28��[����El��&�DȰ�YR`#��?�0^�K,�=U��^aGکw�]?gE8Y+.�෨¤O㸦tk4����������*��q�_Ċ��d��"�PP8Dh�o �Ǯ*=粈�گ�^ 2�p����W-�v���#~5��x�@���ǱM	�<��Ʉ�U�_ι@�������>��L6!'Eo��N�ϷYNp�P��v��7*����b��<�]��b� �R��u���sT�@',����d,ݶA�k�ȶ����		a��'��V���I����ָ���o�+�4��y(�F��YDjklצR���(S\�W7!�#�#;��`�X_q<�}���H���2H`���(z��&3�V�b�[�8@nrM�Ղ�W�I*��Œ�:l�a�%����f/����ԤǦϖT@p#�/�;O�`����`��1�бe�b�˄����n���R<��C�7�t�ya�\����*��cX�N	X� ��E��
�;� G��qiL�tR"�h�u�DU�jI`8*yZ��9�Y��<-�>��� ���GEm�ս���z�@�ͷ@x� ��/�ߧ"C&�K�v`s"*&� �"���͠Sk��"m����#۪�a��"T�N;{��x>�W2���r֑��@ܧ,>�D*̻�x�w&5#��*_�G���(9�p$��������I>Ynyuc�$��»� `A����9�)�D&����v�w�|����p.��$۹��Z������A��fek�gs7ŀ9X�1-"���*�F�p�S�fI�����+Pb�A�U&*2�q�ױ�
��2��$ob2�S5���B�.߁t=�F��vh.b�Π�ܑ��[w��.�.�\oB��M⏏(�O���ygx���b%�]f���9���4q��T<��V�j�QZ1 c��/��f��+�3�?�G�y��n`
��_{V{���K�֛0���>T�m;h$۫�k=�~w�� �����1��{)�B���K��˿��_R얠.?@��>&*��\4�UP��R�Ph	h]E�ղ�E���2r�U2��&�n�1U�5/�	d�Bw>��Q�E��Ұ�jc:żR���D��`ten:��Ԗy6>�7�m��C�� "]�SS�׼��.�Q�_!� �����.��Q>S��7�@��󚉇g��N/�=@� U�:^#137w�b�u!J�~� % ?D���`��3!�|CH�=�F��r��`�dt}"n*�g5�4�gG64D �X���LKm(��ش@�k����-r�����Ӟ'�x�A�m�|���؆��v�W|�C!G*�|�4��Mk��Q#�"s��Wm��:��u�����s�����V���G�G��®��rٰ[F��vZZ�#�ea�o {����*�D&��ǂ=~��~-��7`��9Kb������$�h���n�Y�p��'�%,i@�L�	=�L/���K���t���\�`%S[������Q�x�Um��׳>����F�$rK_�����b@
��P���:YZ	L���x�=�	�#+qMX�*��/_��S��Z��-��l�x�i%S2R�I�b�g���9<��,�^���B���3|�l�Yd{����k"���C���N����.h��	ն7�s�P��1�a�_��{�O���"����P��ۚ#�:z.����,�b�b&�����$�;4=��`�`���Ic�T�M����|QO�`� s<황/�=�>��� �9���0M�ڞ�w�i���`���ww+�{WW��0C\� ��vFD�)�Xg�HN�����<x�=��z1�0y��&��T%�(`PR;s�A_��xqs��V�KZ�O
�Rȣ7󁲾�����O�����<rᳺ%�b�M�3��j@A{�e'a���nD�&�Pp+MqUٮ��9�e8Y�R�����r�I^ш��އ��E��\$M?]`Dp���^��8.2>5��v�x2�zț�l~��I�u�-��P U٣�Nc"������KGX�JVX��2����+"�rT�8a��s���?�c��y�����Fd��E�Y,̨�eZ�ZV�1�����N��hވ���*:W��n�M�G#� Y��ж�0�V̔�<,k�����*W��T��.��[�o����ؚC��˩n���;���8�`D�K�xS�8����9��ң�wp:[���0<��\�1[�OÙ	#��9;R�R���P !/lA18�k��D/����,�����^6{�K�Sy�bMA���g�yٳ���Y��H�^U(�LS ��k8L�J�~/NvHT����\��a�����^iY����2{�\N>�xw����!�v�X�;xɿ��Ŕ_H�t�L:u{�ձC�P����a�4�o�>�3��4YB��K��T�Fz�]�є�i����5H�4 {,��G�b��?]
��lnW׺j���;I)��
��j����P`�E�9�X-���6��ò�������Lv�C=�cc�X���h�&e/�F����1������2W8y��p:#�'�F!��?�PmЮ�:6����Bhq�qPR�R�s
�&|bH�����'R�\D�ͽR��9�tc����3���&*u��O�\����'�.�&����+��5���iM(U���"��߂�3�O�MZת�Zh�wW<G�~b9����eK)��um,k�B��sٷ�!�hi{㼺�u2)Ӑ�,C�7����g���aT���uP�(6�n?��+��-�x..�������po �v��R�p�����i��OF���˯K�Ŭ����%�����!���O��0�K�mh������N�i��ˆKd�����F�>9q;��
�b1Ԫzv��#���r{��k,��� ��e�����b`6��$��	������:�N�w1�Ie֕zRʮ�{{��=�8,��P��S�1E��?v��1r����C�'��ߵ�����^�$v�F��$	"Z0�/|�^=��t�u��7��@��;��T1�������h�u��
�U.?��7(���p��n�b��Ѱ�+
h�`(fF�3=��^Vp��/��k�l���Vz��oģ���#ܫ�%D �۞��-���5�N �ɴK��R�I PE�G��ZD�̝�#�%��4@�+Rm���,�ߣ�w���rJ<FN�1��Ԓ	t�K���j��9��tԫ� �p��,��k۵iu�`;G�����FQufan��s��:?A�_�Nl6C�+7����C��-αNk�xWX���zl��(л�^�r	�yHFԡ�������P�>����i��D�T�s���Ư���@+rT�|�K��#�$1�6��u,�6���G�F�[�V���K�pV�>�Sv��Iy�0z�c��"����`�]���/���� E1�^_�a����j���8��)㫓�N����V �J���f��$�i}�����g����P�eH���Ԇ_�8Ȇ5���~![Ye��Y�t�+����7wD��i1���FkH�������2�H������l֥8S�������=�ԙ� �PR����9�؛����ָb0 �wS��
���&JH���RM�\��W�2W�0[����[V�yʖ�W�I��ӊ��Uk4_)�V���z�}��,<8W�R������Җ,c�l~0���=L���TX���^���8e"߸�r��Mev������0%��^���o��v�+t�U+�"YͲ�vsr�1EqCp��E4ݝ%Kz7Ep�5��D�Ǯ'��M9�#(���!ynHťE����'�[ZE��h�������L�)�[�6KI�z�_JU��t��/PSj�p�S�'�&��m���;��K�zM�����m�"נ�g�����s��nJV�f3<�7ɯc���Ԙ$�=qb�A?�|�6�7�T?�Mwi�����e�i�'�6	��*D5�᫉��i�L�+-ܽn������E�v1�X�Q�������y�2@iš�,���q@w���1X̞"*|܍�͆P f^���e����fJr'!�F2e.���|�gG}~AԨ�㔪��43��7��yo��ֲ��Z��
�����>���L�u� �l`�r�嚮d�UiM! #WCV��6Rj�&t��C����x��;?g)�����:� Wm�����6����:�,��/�(�c���}<>��r�Midm���R�Q8�{ �K��|��^�SgX�Ҷ��p���etg�nG��e�PJ	o���D!O#��j)�r*���i�b?Q!�0e9kM�F�do��_��bOuPcM�|�s��6G
�B��t%�0�U�0�\ Z0�BN`"�P�?����)�������?Q���r�Q�`���a�q%�"}|T�d�0��̧]���i=h���$�8N��8���`/K�!z�Nö ����fƲGk=|�qL�T��8	����G�N����?ޚ}x�~�@G�!^�{���а�z�B���}�5��h6���Z���4f�+���1�L�[�*�1}b5�!ܗ�� 3�]<hB�J�ȫ�����%2 ���d�B���>m��Ҍb*��z�ci���B��$�nH��G�@����Y�W����J�w�������!��l�9�D���R�4��t�Q��A�~��e�1q^�&�&�U#o	5x��i�A�p8q��V&�wƓ�|z�l �W�L��@���Z�&H��x�R�5����cR��l�/�h��^��K���7��t<Y�����x�P`��,��/�б��p���lT�R]�`[�-.-À�Ȇ�8Q9��Q��U���d̂��qƛ.�u�WdF)���u:=RtN�xz#���H| �p���ݔ�~x���S�np�*��P0��dM������w�@�V�����O��r��)��+.hx����2���v������N,��l��#9���7��s��������4�6���!���h�W�8���a%�8�Ar��m��q�-�9�Vt�o ���Eg�{�}�`���2T�	�J���<�d#����`����{�-�em:����(�i� �卌�2���� x}t��{��D��q/��+f�� �Lt��E�R�Oy�x�DԾ.=�#:���OCb�P�~`�����z�A$��)����7��v�ΓJGʒ1�W�Q�{#7��3�G;���^42��Z�LxBU��?�"���E��RGg�G�YX^�o�@{K��b:hɘ�iĶNx��%������e5�p����G�i�SJH���r$Z|�����p/�mr���Z��I�9r,w����G��a|��[�u��x�k�c��9d-��u�h�Lg%d�F��Z���j�-�b�]��y���jq7^Y�o5��1-9noVx���Rl�0*,���r�b�$Ș��4�c� O�R*]Y�(���C�z��2H=��W=Å��3�΃���J�n@�����<��ܷN��fT⿊�P����oK���H���ǣP2�|8�*��v��$׊%1q��{� Y��px�1�� ��{c�y�O�!'r��Z
L�r�0+�m~��;�ߥ�NfM�����]��Ħ~�d��;[�YW��8)*�|㙨�^ ܅�Kz���g��2��,q�gIl���p˸��P�{+F�ŵ�/����ڈ�]ߙfr�������f�9� ~sc��1._��Pyհ��5����[�B�*v50����g[XZD��1z��K¼U����ڌ'k�W#6�u�K�~��[?qw����~ӓU��ñđo_����p�|ʭט�|�{����.�]g��IE��4	�z��K��4A���tg�J�#'�����u��8�m�Kˎ�v�n�q�΃��K:�k9|�$�=Ջ��8P;����ih���>= S�&�`!~�O��	�)xD������WY;����$`���9�y�a��B(�d�����,��_�'�����v%<�3۲�|�4[��=Ș���a�2��y�I#�/���_Q����c���r�{x�M>H�b�:�+.���K�����/?��\0�C<��Tu5�u���Wgv�����X����7iim{ ����1U6���SO�Gp�ɇ2p����5!����NQ��F�#��l-���$�Ѐ���Fu�z���@�|������6/��-z{�6?�O��:�	�ݴ�f�a�D̵w�c�w�5��I�m����(��K�� B���Sg��{�����B��}����F�8`�,� T&erK�ctSn�T/R�#���I�F9��@�A����m��I��"y�
馪�dы������\��3P�����s�d��jƜX^x���D�T��軔�A�%ס����Js��r���L9J������k9�d#*��71PM��mf�sE���4c /��e~n�#z��bï�Ox�|p�}�W�r��m*�t����������T����P��X���& �!oַBy�$�2������Z1��Ad2/�簿޿1����%�I�d�U�Z����E&�l��-�*��S�'�M,��eh�y��e��F�)���Qw�H\A>��I�@��U�l��������4!G�R��9��9�mfլ���@�hO��-�{l����-�)�O�p����}�|c��\��5���c5�s���Hf;��=��;Y��b��I<MM�ӉX*��ņ�vi�S�WVT�&h�F�o,�Tj����<�A��{��w;f�n5��C}z����Fb^K��H�Pt��}EV-!�W>+W1�m�4�"�|BՃ9�*cJ`"{ψG���X���넧!^M\������F�ݺ��Nz:���t[�,yp�G����	˷Q�������W6$)b�~��ȁ~u��`��Q��I���d7! Dk���b�x@Q#�>n�@���Ԣ����cr�>g�=���Y��q��|�i�s(�Vz
�ב�],�Y`�C�vo�[���C:f�p�L+�_ �����"k���Ӯ��O�����X�E�3���=�#�#�'͌u�޵y��Vp�%�"O����:ɘr���hx�l���v~�C���:��'���Ζ+#�Sw1s�c|�;?��7vǢ��Wn�!�"��|ç��ɖ(f��(|X6����ǒ��$`9F~�)�t	R�̵������]�_���+�jZ���ѠԄ���ҋ��7��g$߀z�Bw��F�!hub����<o_�J;�j�3=O*M"�i�v��U�C���Y
!0Y]�@�}�`_��'�C��J2���� ɸ#�A��a<��]J�鴷�s��qyo�2����q��sDꍬ=Id� q�#�,�G�aS*6p�2���J[]�
�/�C�Q�/�G>PS�j�UBS7;��N��J"yE���4{@��R/u,@u�K�욶�4�٭�P`�ޟ"ӳ۸A�O�������z'%��5N�$��X2��t��h�BRف��&��i'A;� �����K��(;�,���"�"V����!���2�%���of4E�mub:�$�FAg�kk\�:�>5N@�D��W�<69��.v��ފ��}�OF��2���?Z7[E�F���c4v/>��Z��@leI	:���� {j._/JӏR�CS2��q�#Ы�hMZ32�`r�H�Wܝ� S&i�,��Qn���4E���v����c�e�(��(���7��V���zV��;[��X���h�'��/��Q���&���cɨ��~S�s7��F ����{n�$n���qŀ'�]WΥ��TC0� Uh���wN:�ԝ�4��Wٔ5n�t��ϝ�������b@I�����\�8qt���9��k��#3�K�(("�k�qU��L	�b����+֛��#�)_�E�~Kn�y�n��>)��?�qx o ��3_J�m�qY��}�׃:CJ+�<�Zp����{5���� �dՀP~�%����a-"���es�VW�j������(C�JW�`	?�f�K,t��L�e{$�vl(&'�ɤ���O�$u���i��|����ʿ:8���|�X�9�M+�I-�R��"t�(J����?LH[�*V�̢����1��8I����`��od�Z�Y�@R��Mʰ�jC��ꚥ�"���͖��_Ҟ7�5F)*/L�(7Gt���%�b����ҕ�g�p#���d��Ux�y�[�g�I��;=
 @�����$����ۋ��"S �/����F��g�=��(]��:�f����_�q�Y�ѧ'�H�F9�sO�j�S]h(�u�|����l��*�n�oUH��t�e� d/Q��o�x�*��^�W�6K��O�%bQ�-V�� W���O�c]���7Etfծ�B���P�ٜ���-���Fi�ƈ�X�`F��V��$/+�O8(�IsJ� xA��zY�ԯ>�����ʌfɵ�q��Ɔ�E��5� �ǸŋE-k��N`M�,���Q`DqX��k�AJZj|�JVb�mWWbҨ�>�ak��6Z�	c��#�ֶl�T��JΛ-�5���^�������������^�k]�U'l�1�d��ɰ���{����� 2y����0=�8��L�L�nX+�nEk���⑈l��2#T'�m1�v���q����X� ��Ł:��o��<�g��@���lHQ�����^ 1Fr<�@����]l�
��O0�����+�K��k�>d�	&�a�P�k.�i�r�j�2�c���@��z ��KI��$���#�x�.Xb`�v���Z"�6�
�:�f� ����C�6�29S�mr[T�7P��H�/1�k��w:I7c�I�fJ���!����|���<�����&r@����y�H�&�8�H����F�(�3�Z��ϑ�<?��� {��,��,��Du6Sy����t������+~�h��]��\,���S۾n��yz�K5$��Ly�ց�����p$��������^)ވ�j���8o�	�\����}.������6��~�c�~8�g��尖UF�<x�O+I
	�ʀ҇�;��r�q�[����6:���Ikd"0̷P�h�t�?�I^����* �$��--��ϙ�bK�S��.���y_c�?��N�:�2^�� h�3��b��*PKB���9������.�E	s��\y#{�;p ۋ}SC�8{;i�8����i�S���:��^�.�u�0�# �)�t�y�"�����b���������%X;
~��	+D�/ s���6����ֱ���Tb�	_c �
u�������}S
�?K�e�g�n2 �UfY���Źz}K��	��	�U9��ɟ�?��@�Xbq��c�#!N-�c�@+o3�Upj�'uQL/�>L	�߰b���4L=K�ݐ�D�R��%�r]Ԝ	�X�	����?vv*	%��?�PK�H� f���>�Xo6Km�I�c�#��H���]2x�Q�Ҩ���+pG����L�a�{�T�IYP�n4̉ha��!�.��M���|�G5�L����\{ ,
�.����JQ�b�YL��L�R	�����k���_b�9�.����7���%,�����T�g�M��u�*�_I�]&j��
y�H�;��	&�CQ��`�%���vL�6߿8_?�Z^$����Uy��[k�ډ��;�T�`o�g�I��-�{�?r��)��|	O�jwZ�`KL�(�$4�[T'�r�5��po��6�u#�@
*Vu5o�A�]�����,��q�%�톧��쌈�Y��r��-��4�jl�:����(��얙wz�Ȋc���Y��~i��/�X�Y��SA�4bT�܌y��C�;��,w�mc�Z({������-� �X�t��sˢK��q��?��F�}��Aw��F�v��(��p��[���2��qJ�)/\ �#������T �����:{᪁2���X��Y�T�_S�3��m�:洠�XD��6\� )X: �"��yl��0��S���y�s4��o��ǈr�QI%����=?$�u��Hư`aC�K AX>qi1f��B����?�T�ܫ���L�MR�Q�v+An�_Mz-���'�i�vQ��P���p"�@�)B�; �H��ya��a���%6�Z�&kR�_g|��KK���2���$�hڤPXÂ�s4v�c�|�L���k?&a;)
A��GkI�$A����1:�4$��'
��f,���I<�y���D��;J���;^�%g{�>�(��3�N�A�_7��& Rc�>dP�ؼ��#�����z��Ϣ�P�e��ҙM1�'mL�P�����M�9m\`�%USn[�=H�_
�h�Pi�/��!��� ���7V�Zp��x�lLKhD0���o8h1�@(�76�[�+�do�oww2�e�ē�d!q�z��=V���A�W��R@R�)=�B���eRe��K��)��}p�F[L���Y��qL{���H<�P)2r����ûj	Z������%9�}u��t��k�nH�Y@�S��Uk��e@�.<��	���j�zϋ�g1r�e�Ŭ���z����b/	����ڰ�b��+~�t��w��ւ�t�/�3�ڪ(L��=����F8�\@�S'=��O�rߜ��Ղ�*�w�\�(&�S�~q1^�f����&�ޤn�
������S)�[�֮JH�.!&��(��aC�pl�ZB_�et����1=+W��C�~ıh%���@@u�]h,qZ�-���Lݟ�+�Re!�:㠐��k�eI��2B��MU>^"��[��.R({��Jϧ�o�oc��#��a@.�g��``aT�b�_���U���h5s���B:Yk5��tk��ep���-��h�R�ALͬb^ެO���V�����[���B��ZU��uZ�lEӤ_�]�70ʤ���%w�0��D�IQn��]cޫ�+��[��f�$S#��c���f����`Z%�5���!L�����T0o�^ן햗0�&ܐ���»tl�؜X��{g�sMou<�
n�v�yW���~�.����;��l�
3�oZv @z%:cxq�<HU]�]z�P���c����q�-�9]WK;�}��O�iz�Ey
÷�y���没J��&n^�x���j0:�ʒcƺ ����z��414~���������͕Ns�*�+膏��уLQ�O�#�Q�ߢ�_]�X�9&���E�O��ih�'�7S8m4b���%�k����I0_qR��ɡix��#��&w�pw��<�U����v,��X
�fgΚr�%����f��6b�\�W��{0&��+������;ʉ|�G]������ɸ^�?<HI,�^����dɳo�ԉ����;[��u�m�Z׬Ѫ�)���J�@�*�k#;Jg��~�9��'cH�y'�[�E�)����Fk�2�����j�U�&8`��ӛ�˥��\���-?�����Ω�#��;��=Q� �7f-�|/���I�/QY���Ok�lZ�f�֧D�~z�^�Ɣ����� (!I��e�T���kv�@$@q�&�V�����mJo��^@*��)�����L��	�oɮ�,�g�#���s]ϡ�G}�l���3q>��������<|�G�V	�h�;��7x��R�}�;���k���c�li=RQ�eN{�ddZ���rr"uh$���T�,9��nķ$iBJ���e�]դ(�^����9�$�ҺV��fŎ�W�.�ž�jv2͠vA�	����4�W/~�*��[~�du�GY���#ҽ�q��L�m��/r�<or0�Bovzܼ��0�Z��GG�^K�ێ8�+���,�S�g��e*�Ύ]|�<y,yv ��W�ζ����1ҮG�����MdP�2��Ԛ޾7r��
K�T��I��_���d����(�H���|kYQ
Cw~�0p��y#�Ђ�ף��S=�<MK���-�#��`KlS�80�[�����&���A`�*�'�:�J�	E1*�<.��	e<�k��'i�p�ⰾ�;vݵ
^�*C�'�T7���:�D_�ֹ�v~Z�ptd��(���w�Q�q�v�8�]�>lRe��O;�!�D���&UM��קL�{3�2i	��H�+�_�������YO����m�K�2s.���!�=K�8D�sB���ƻ�����=����ރ���n ?�=%_�q-������v�x9Of+����x�W&Ȕ}2�
&�Yu�W�:�[I�Q����˭����~P�u	�� 6��X�b�gux
A�/ԙ&c�_n��~<L��S�\�4���8�Eo���VzS;3�g\��ζ� �!FO�%ϋ#��v�ɁW�a�|@R��cq�Bݷd�X}_��-�
����/lk��Y����k�9��,2y}�z|e�F3�kNQ8�nā�>V!��оJi5�=��y�t����O��P����'��b�B������s�je��<a�$:¼L6d�*�DK�O��S�ѫegW�G��M�'QR�dL�a��#0�J7�&%=�S�3�Z��iiάҥ�z�҄v��t��ϻ�$w�,�"t��`�_��C�Ul�O��\�,���C�Zm�5QUډ�	���I��Q#��!�n(�T�t�Q��b%��$8��ڥڃ��J�/j|��P��[B n���y��*3~��&3AvOx�N��¡=��^�?'�b��o����^�dkYu�ð����o�K��� Ss��b\�*�\Y�ߥ-�}�N#�Ħ�7�~�����c�}������_�|�F��h�_I����
[&z`K���[K�(o4�!�В9�Y��W�r�S}ȥݶ��^$���T!a�.0�鰻m�o�y�J�Q�C��<�*u�s"[�-�>��KT�1��=᱈�k���=���H�c o����+���П ��z���ˋ�ĩ:Z��à����p���8)�WP�R�6sP$����*YT��pB�>l���f��m��%f�:D-1���X�m������K�׊���%e������)@'�YDU��}��z~VF�&W$&Ls��?��'H���hd;�Wu �y~<Jǆ��b>��$�T$D�틽8�8b�q�Z�f���Qkh��ERp��k�W�orZe�_JIR.XY�����o�d�*��T[ݕ.\��D�q
] б��;�T@4o�/�?�:9�n���#lך�At��|�4Dy��c��`�jRНK'bOg![��e��G��j!�jDN+���䛄��W�����{0�T��
��F�@��EQީy�������o.�N����ʓ/ބ~7�%��[H��]�J�������$�q��*����E��#��}t��C���k)ʱl��&']�n���s�7M��h��pR���� 0�h)�>�םF�U��SG�3�Rt�O��v /
lDHr_f���|��%������ �c����+��r���g2����.V�Y���'��b���� ��r��.���&�Q}��%���� ub���PX��Ns���5��\%j�(=(U � ����ʜg�j'�H�A�b������{�vYdHntu�?���؃�؉I���8�h��K&���[p�k��e���X�gH�X�P�g��x�N���Ҩ�R��!�@�O�bb?�m3LO�[f۱Tp��bz���|E����ϿM���p	dՕ��>�b���!�+�� ��<VZ��ڼ��l+N-7�[�y�DxD��<`��Q}���.��3�Ħ��?�k�:�����3�`�O���͢Q�De��[!gH/����	Q02�x-n��<v.b�F����v��T����d�K�ڃ]9�~�{�4���]��D��(�.1�N�[ݹ�ֽ�;$�$UB
[ͨ=��ܸ(!�Z6�C���!�l��7�`�$,xC�d'�(I��vP+4|e����
i|�;�'k�Cp ���SAZnu��5xRλ��T���{\���I�F�AJ�c~x�`P�Z�=?�1j71���j
�<5l�&%"�����ϨN����Z�H��A��TF�^F��Î��mdC�_@ko��v�K�eI+R���X��qH����Q���6*ҿD��H�Z|H�F�c|�;|�/+3%r�`$��Ӧ��_L-�VS�_ݥ c^w�H��+����R�-�W�*�4���ոl�����m���!��E���E��3}&<��k#���?T��-��ՏX$3��B��K�~Ug�# �C�\�uG��R��<V����jG,�U1�s,��	XGf2�ī�W����{�Ĝ��@�����I��@�	 �}�r���`�Ic;�ߌBVI��T����UC��o(��Q����3P�������������o��U0��Z���d����_x+��sePɪ��2R��#r�\���,�y"]���u�f��
���2 ��Z���%g#�%��jI0�d�^����s��&.+>���T�l�8T7K���_�]�r=rB��
��R	��u�1���	��JT�Fd$�- ���=��-����A\������n�[apj8H�uS�պK�;�Oα
�)S��-�
��0�Մ�D�,R��\�=;2�g|#�[�����v5�PQ��M�g��[��^xAH������̻��*te��^ �˛8���f�"�6$7꯿��y,�1�� ��g��R[ۆ:��Χ�������|��/^{���.����t͎�bU��~r��ʒv�&ɀ�����\T/&�C��H"2v:+��l\W�]�%y��R͜��C���C��'��j�[V��ה�=Q��4��7��ƒ��\�� �K��Рz���q����Q�g�h8Ѭ7$�
�7l<�h�y/7Z%w�������`R����^tʷ�M ��7<�˘1@�<0a���
b��dW=$(�s�QYQ�F���Yr~=���>Q1�������t���>�z�D2��C��\�>CjE_�R�X ~�o�k���Ɠ(�G�N*˿ԯl�O%ڑ�	��wG	"Ġb�S�p��Ĳ�z �5~�"%�K�҃5�\_*���_��������%�;f�w�\c�Dn]�:PԱ�1���T��ON�~�6cq1��T�	���]�9�R���'V�[��y�8��D����`s�	��V"�9S,���+�����:h����D�7��=hF$�!�պ������kP#*U�sB!1?c3i|����V�mP�z���3��C;l��gX^们Y��^�:o�l�F�w����e(CT�O����D��C���dv�N��$D��h�(ǚ�Q�π����_�A7�k�f�+�K�?�K��#��-�a�!D������ѡy�1�.jK���f��d�"qa}UF���_^�=1b�i��fb�ܓ����y��7�a�<:�>�=t�D���� i�QX����iPȜ��Åމ�P�.�x]�A��`hވ�(49]S*�T�Q[oT����-�f/�0?�xH��t��+��,&���z^܁�Ĵ�&o&��ۧ搜�o���mTc+�;\Q�絅#A0@��d�2���s��`
�ˤ�X1��h�F
��սFB���z[�}T�˻6~��M�؇=�Re@�$ߗ���H����j��ȕʦ����X���"��jڮX��ʣ8�(�A�xh��a?8o�N�f��w��S�g�C���bQ���.	��Ѧ�/֚|�MBl��	k�S��cnn�����M̱�u@��5��3�o	�l���)�}kҩUj	�wF�]+[�bέ����K��qR��� �i�$���|��.�͢���-J��V�ecD��حT��:(S$v�&T�v�Oe�T��%)�f�۴�^�h7��cv�I�
�P��Z*:��2U'���,����	�5������7�6��U�M�d�(��x�Uzچ]ކ)�dG1H���r�r��8eT�M�	��?O��i��i]�M��Khҵ�=W�������/ܙ L�\*��iRd�(��=���7�����4��"g�F�F6��s����iS� �N���jڧ�4��P@{CUȽ��8��"�܎O�>�'�ɤ���̱R�Y�ᰖ���v�=V�K<�Lc1�K\�{9�n�Y�Iu��f(��r~[��������<j ,Z�m�����|[�r	��f�+�}�8r�]v_��1*�v�е�9"��RA�����	x;��$Y���A7�U5i�(<ђ;Y�����C@�,}�E��sŪ����V�Ѭ3\����N��W������J�u��T$sɜ�[&�^��Icg�C���&3�`ס6v����/V���GRM�����<����1.&��C~��cwW��`�x!��7x/�,���?��~��P�Q8	�&M)*7���_�
���ӸQмz�sr!Rr�ʑ�~��2��R�w	���w&����YU	�aZ��|,��x�HoO����#�s�*vz3 �2��q`N% ]x�@QCi@�˼RJ8��篋������q,�*�y�KUL>�{{���\�z� ��?��$>E_�~hN�^"�ԅ��q�H�P�`��R��8ז��mǋ1��'����e��҉�'1!����hE�R���?�6�7ġT5���ե+�h��X���)Ieݤ��D�΀�E_��8C�_⿠���} V�WP���}�{���XfCe�ȥt�j���hܺ $H�5a�7�X8���ㇿJ�g�����w~ڽ�Ձ�i�Bvpc�c��Q�cc�C��-�7���]������s�hLægb��x����`�AtZ���z�e��	�$����T�ˑpn��4M�����Y�@�A|��Z0�R�Mz8����%
��f�F*�һ��m�?��(�P���jPڨ��c���mkl���r̈́�=�dB>J� ����H���VmX.��	=Vl��K� F2]�F�� ��\����(���h� ��!W0�WiuiV��i���{�<�� �ٰM���遲�AdVY�߷�Zm�����υ�����XѬ�I��Dص�{"&��F�s"�!�`so6)�<�,L�:�v�F�ݢ��-�ҸF�[2�zlT��~{����;�Q�ύy2����6F�t� ���w}�d�� Q����~��I>rw����T�1���uZ�=J2��9_q���8����r �K��������TN�����ܭRn��Ǜ�n$Xv(�_���ǔ�GW
p��|�x�Q�13�b�^�G���2s��F_;��rW��CM�j����Jܾ/.���{���<2���y1���5㔪Y�;�v��],�wܗ�춟�~X /ر��t�y�4���j��nhI�%l\���b'ĵ^O�%��:s�N/��i߀H���.`=�<sԉ���Z�n��KH��j�oL��=�~�NA}���,��5�k�mʉIy��2FCC3Fk���3�h����"�GXۭ�k��P��,���\��")Y�f���Gܯ�>1rl��&���k#�q�B��(��sl��1��/IBV�;y/����:�o��=k!ɻ}��k�Q 	�V[鞛7	�B�����|�6[�gPVz�T,�����Y���l�hL0�#��F`]Ur)��6Zda��
�4��s��$5{�ǰvU�����ЫT���i�8w���y�udb�O��}{wWLx������[�q���?���pپx��-+Tζ�4[�lu�̊��)�͓���ۄ1����d:k�v@:/��#J�>�z/`�<�u�8�r�O�Ki�>��+�@jD�t�lW������q���� $�
�Tf��@,�Ȣ��Z��!Q˿�yɚJ^S��[�cIFWV�U��������������	�
/)��� gW֫Z8ՕJ�	_���|g�d�(^0�+�b6S{k	 ھ����z����ͬ���ma�c6u�Zh�)r�|L\1ٻVGebq,H�����ntߎc�U}Wcy�2G�3F���,���!��i��h%WL��Qr��x�鞵�R���z��6i��[�z�Bz�B��`��D��S����xQ��ی]A� k~v�b9��糿�"�g{j�Y�uw����g�0����OZIr����ӆ��ݏva�������	�]�}�9z�=W��}���#��jS�WC��E(�*ɮ��?ݶ��0�^ڽYy����񤆃[��'�u2�z�*jK����ZA��Ͽ����q�.��Z���W�w���yq�h=5BQ�e���
��v�Rh�8�Q+<C��<5�dg�.�.-E�p�޺��z�q���p��ވ`c��u��M*7�6C3
Q�leA!�_�Z�Ի������]b47�W�%�J�m��0���6���o�����Hi:{m�?8�
D���jWq�roU9�n6	��Μ�Y8e���SK�V�'[��\4=K04�u�Y�U/�7��6%.�׼��IT������*�����"Yo��c	��� �nˈ�_`"�m�v8뒽q������F���l���!���9ox�E�s�����v��͇p�[�M{� ���7��0W�1D2a	a����QuT�bp�����k����\P�����g��9�4<�MA߽/n��o��8cD��/.?�䲙�_ɲ)�S��1��;�f�鈵�I�v��'�pb/�i���a�1�%�S�$�4��Cj>oN�4e�.Č �Z�8�jB���+%��ץΓڴ�-4���"R��0.���������	^�ϖ�륮� ��� �^@������2D�j��	�Ć^ ��Hb-�w\@6!�5�%�"�5F��\�#�ِ�;���̽t ��D�kE���lX:����`.G��K@�)�0�˦2į���e�!M�y"�#t9��},�.���t��\E� ��#q���8jc;�C����
7��-uu3��,�	B��@�����8�xe}줍��7�S�\�8��9�}<Q�A,�����⊓\V&����;Lރ��2A�B��wXq솎�L������9yik��ǰZum�3�P��G_E�H�hb��o��0�^�@��9�[W6Y��h@��?����	zu��@�	�V��6OC�uq��&9�����*��v6`�@9@v߁ �Cs�?
��XM(��R��@f1��oI����M��TR?��8F��?x>\}�|����<j������-ߦ�L��ŉ�Fr:y̻��)�X�n-�8�e@z�~���Wf+�;�vP�x�dU����	rlQ*�<�����ѷ��qP�(����a�-]�&A�ƙ��j�����@�E��� �H�A5%0Ppu��Q����e�6F۰��m���`���Y��?7�֫o�-�{���kKi-�;�nպ�XQ�?�3�V53�wK�"�p]�M��}ֱ�N�N'����SQJM�Aws��|���y��&΄�A|⧣9t���Ǡ�H&�S��玜���8;�1��IΈ>b�T��C'l�;_w7U��ڲ4~��1�W�����f��gO��o��K�!g��K�<���5/g(;�)<�0�m�3���D�~�=E��
�O[b�P��e��?eVd��K��/�c9�ͷ�~H�;�cH v�$P]��$��~��D����2�ɲx|�j��und���Yќ_�ᯮ���U�3#mÁW�w@��Z�,�����FՀ�����7�<�޿E�����%���&���@����mӫ���gw����)>ο�מɟx�>��/HS�[�:�/fg3@Dr�m@�����Nu�b���A�
�VU�I���]"�7�.������s�%s��F B�����+Q�p���S�C�d��\��$���!ʍ#
���
��3@�~u��v�ؐw��mA�փ�٩{�l�YW������!�w�W��M)�@�
�S�#]�ۙ�+���	:�ԉP���"�M�+c\/��ͮ؈�-�(.|QMdP�$��8�L�o����X9�Fnz�~UnN����Bf@-��&�*�_A�2B��X�#�u�O�Wem�I��%XO�"R|Y�Q`�VM3U��Bp��nF����U��G��l�r�K���u�, 프r
�!�։!]����QM��=-�_Y#�����4I�b���vc�'4�S��hLH���\�V����G�k�
�����D�G�s��m� ��|��
�b$sǲf�߷dc%�b?��C��[aWӈF	�1��f6r�D�CH�g/����u��Mbӏ�� !�$C_N���~e�Y�=T��\�����NSB�iY$4��+[e ���X����"s�:]��L}��t�%��/kw���4�E�(��~�h�4�s}w�h��ي�g.�0���kIO~0�%�Q��F�Bj��!%Z��hc�F���{!��Z��b���}!��?-����f�����
S�*����v�i'��h���>�����+$�6�����yx?��V������?�����G��벝�a�k�y4Cm��6���or5�.���I�����$���7�w��rݳP(O����,�2�#�n�0J�^�t�f�W+������J�>�!p���`*�fРL�T�͟����_��(5�y�1�IP����Dy��~H7�f�QG~�Ɯ-b�ڋ�5�)�L�)"�]�'v�����7���L߳�<���`Z�����|�H��d�a/l^��v�̓�N�8���$�UІ��4�.�����o�����C��c�t����QpM^�D�R����K�7�Q�)�S^N�	���f����������e��Oܡ����p\�'@���Vr���� �_�^}M�v�D�����_�ϧ�
Ȝ2Z�k0�g�����"�����!���D[C��5�];X)�3�g��}W�xC0��9tF�P��p�����އ���efs���	��P��6�<��h����]1V��(��?�{�G6$CKe���`�a=(dq�[�A*��iҶ@��ܑ��:�?�9r�.��xJ�4W͔�g���������b�Р�Ī]�'󈽐&	s7� �$����������6o?EΨ�Q����7���#�`�1j������]���x�8���T�Z�ߘ��Y(��7m��Y�%8DI&�`Y��q��3͌>�ʻ��5��Oղ&x
]gÊ}@��k�/ޥ�.b�3���������L����z�{��r9�.?J���Fz@�h��\w��G���)���r���k#��,��ިq�}k_L��] �K�^��8H7�ۘ�@�D�sp�C�1�|�k>�g"�ɸQG�TI��+swd�H7j����^%�c����EK�����zI�P��q�1�c߄��Kũn��^&c�^ͩ�,���U��pv
�{����#ohZH�S[W�����" \$}�0r�}@�$b��㜇��~�S���������		�I'	�!���F��)���$2�VQ\���T/G푌��?��;+�wuJ'���}����J����>�< �ɇ�jV��.��B}�,U�'��q�����ݑ̅���4�����&)0�;x�mZViT��JM����R�,�z@�z*�d�Ҝri��	�Mo@rķ�"_Rc���2��-X�`�|$6>�3v���FX�si�bAz�̤U��^F%�!�6��b���"�6La��Z�x�{�
�����ތ�c�S�}�&��U�E���6粯���gJ0��T<� R��8�3nU�@	�J��q?&��Ă�^�{�k(D�&㸻���1�yѿ�8w=�.ou
2�L�9��e�\�$=�������٪[�&0�?r^Y|�l�����q�ɪ����.}�a�^��]�&������uWv6�V�7Jr8=Z�Q�Kn��=�9).W���*;?�t$���`����*�P��x0�!���v��;6�R��8���N�|i8��׹���<'e�'H���V'�Ͱ۲�V.����&I+���q{2F'[�u�v~&Js?gh�~q�ؐ�
�ϡ��<)\^�p�X�����;!�=�1}%��.���.g_{��5}Ll� ��嚱$R߾9u.��D(�HBN���l��@l�E����+�M���D�g�����c�<�̾�hvc�W�"p��2���Ƣ��8�r�K����Y"#3��}.���)��+0��X�.�'F��-�9�8�vk��m���.�L�H��m�k�	�%��e��'�[ӥ�=/�e�� �lU�V1�V�B�9}Ɛժ0���D�'D�����bp,S��˪j)Ftcp8w����8�`X{I4��J=BT��`ɗ�ft{�V9�J�b%C���7t×8�i�� �^�cy�'��Ы�m�E,�k��U�j�d��&����c����&�thœr�,WL _�H�6���`�y���KP�aN��2���Jf�e�+�V�/���{;>pJ�Q�|�X�D�k��I(I�|ƙ\PI>�S�@\��p?T�B �4U�z$2���i�}�[\�K�M1�#X�z�E?`aq��i�SN�?�����F�h=J��{�.#B���f"�{�^R��8;jɘ���sh��6Vћ�ԓW�-]���	�1��8\�����w	~E� ~0��0�i�y�Z��G(���L�NUt����V�j�[HԖq�Z6eH�Pl�C�У�����oI��	�/������'�V�۩6��[�פO������q��xٲ�MN�]�`t�
J������}���5���|��l��&1;I�$���D�P��?������}�����9D�\����۵)ڂ����$0����w%���L\�(���B��B��l���d�½��vp��Qj�*��j��V��U��7@���lMo���w�w���zcImj�W�&���r�8�zG�҇;�G�kf�-_���K��>��,�����v>z����y����H���T"�T#"��O#L��/.b'ݪ�uJI�lcU#Z��T���x`2�-���9���9�1N��xHÏs���ďg��~��,.o8/����@��8^i?Ϸ4A��w��Tb	0��W�o��s�d�1��HJҍ��ɝ�E50���bꨀ�N���k��.��2�������;��U���=�?���& 4 ��� M�қȀ��ǧ�s��w�z��l�B�#�'���F|[�����
#,t��zs]C��q��=�V�/U��(L�V� I��ޅ3
e`���)4�:�[Դb+�0�f���g*8��=Q�5m����Mb�mݱ5d�"��F�!9o���V��99/�i٘�
&�RO������ |�K��İ���"'�U��&��ce.�jYNWg���/f�,T��l��#�[��XqX��{����@ N�=M�>���j��1+L�OUhR&]aO\�m��o"*sM��M
C��&���F��jʽ�{���6�ċ����n~�2G���j�Q �4z��G���ʅCt��hrR�M�.�JhB������r�{{p_����XH_�~m��R���<�vw�"D*yu{_� �V4�<��%��ȶ,plU�~=IdpȣSJ�)]��Q��ykmO��_�-?E�B�y�b\SA�I+;:�@7`��.�xZT3�� �9�M��:�_��A@AR'LuM�l��˂��z�dr��!jn��9�= {����|�#�$4���B�O��,;�ѣ4fD	�U���L��

�{�8CQeJ�y�IaY��;W�O��� �˖���C��
��������V�tM/��,��I��s������O*O8W�����f �7	���ɚ��$�TC^�%3>7����rZ�jl��(��J�Q؞�_�V��4d�8�Sq�Ǣ�;Cs�)U`M���c�B�9�;h�Y�Y_��ꆤ�IT��Ā�r��������fe.f~����pQj�0֦7�z��'|�g,��v)�Q�&�ˇ�cGl	�����
�p �Ԍ��З���ا���	�Z<�.h��t.Q*�
�u���������}w���@(�p~�B����N8-l���F�"����ۊCrya@ �P�U��I^R
�?���.�@�ȃ�p��CP͠�<�k<����N&�GNιA�5-�u[W��fM8Ҹ\�\�r�.�f��*�Ħ�,4�NqP>N�c�T%ѝV��&`/��1-���C�&XYQ ��|k�"{%˗~��Q�xn��ROT�7���,�+
���s��+��2%�{�8&(O�~&��:��$#�YS1#��~J�g�%<X�Oo07�dy�������F�~����$a�Rx���\؉��B%�u��MK�P0�L��-'���m2��J-xD����X���\P�0�*�오g��$���I�[qM6�1������$��臷���]W� ��/{�A*�\�op��&o
��1,�$��w�?�
����$#�O�}�����[L��h#�SQ���md�%�����ns���'��)�Ll�Wi+
�<�LO�M'@����+��Bަ706���1u�c"�in;�-�D������1|�B*��3E�Aq�O�8��ߪ�f�@��q�����Kc$���^P���:��E^b����.�X\�=��c�_�!uj4�R��q��^��Ō�T���6W��܄Ҕԧ[�
�d��L,u0��ŚS�� j���Sh?����|�yW�d�U��q0����zQ�+F�J�7��܁j���� e%fx\���@��#��7/�u�;�\ڴ/�'��bKfgB�u�%�G����}"F���=/,�����/\6��-�aЙ��
����]h����T%Ce�/�>��[�DN�LT�!��q��.�#,� ��vt�Ֆ����Q��P�m�y3����Z��m�Ը��>�u�ʚ���4��ư��L�7c<G٧��$�V���اh{?��"J�b�Tu"��!\��me�@`ʧ�Z+�n=�Z�Ye��<�b�&��1�aZi�XE��-��8G�f�#��CQ�R�W�)U �܋���Y����_bG�����ɕ����9��SG˛���5�9����r�r�w�>a��D���oN�T�v��E��Q��PͻJ�� P �,���Ӗ���2�H�y� ��$S�}��5��0��߃���*f�7�X/m2d����Z���CU8t����"�����_� S�cC�ɹ���4�!@�r��!A�"����i�������������`#�/�)'K�,>B�� �^�z���zM����ǧ4�)���/SҖivY' ��F-��Q��`&\���ٞ�	|����%q&�<1�N�Ҟrr�#��L��l�A��n�*���j(C�KC����՟�:m��
{��B�\#V��sc,0S�b�&�pHN �i�O��@�J������H�2�Rvވ���� ���$�;`:9��]�����$	�����+�d��$E�K���mF�l�0�i��qeK�7�w�$�f���--%�*������P<�T�{*�x8�h�#��Y�رREV�1�޲����R����!���o`��"g�ZY������/�d�:	Fsz5������(Q��l��5��扏T��e�)������ݙOt�IY� �{����%Y(K�j �k���M�ڈ����S�q��
�e���y���}8/i�>i�� c$�V�F�	���)���dy�xK�2���|2���6(��A�I5+�D�B��p�#V!�����%�v��O�P�N��*Ҥ�nE�se��  s ѫ����- 7^Hߌ���b�#�~[{���#
Z��*���E�n�?*�0�̮���|�jl9��pHn)	�1�������w�?�c6^n /�doF���	4�K��V��ӑ��0�u���l@��F��/wp��7�(?]vZ���euz���&�EN�!W=�(<�.&io�m�_����U����d�8���"%)��sTa��NڿEJ=�z�C��w�D?����!d:�#W�����Kf�|&�\ΐ`P`�}��yZ��E��]���| �11�6�۪��jy��v'�&�;`[i�T�*\ﳌqY��K	�Y?����!!6ą	�[FBtH��8��]= NJ��M�ҿe�������U׉�%�2���H X��A����B}÷��	mКw%WAg�y,�����9�
��������+Ah�� ~-��< ������L�W3-@���S���X���&`�"�tv�1 �6�ivRp��F��h���sH�T�L��:F�]������ ��������Uty��N�l���3��V��&�Iy]c��=xG#���x�����▦���`���l�W����Iy�٫���N���������P\Ađa.�t�0��3��.��|�08���ThB<Ү����K�_�^��&����;ږOd�^�~n��Ʀ��y�8�^�?P�T�����4{K���Z�Z�h$`ޠ�����IN��7��	�*W<�� �R)<�S�-��ݼkGmppw
�`�e��, �5����JE����qi$���c�3�; f=dJ�� ;���"?��^~�0W����N0�j�Y�Z��ݦ�*��.���a(h�"e2��v5�.`��Z��͓w��aI<	B�T0�_��)	�yR�䡩���y#AkΧZ�KV����+�T}dhA���˾BF('����H$�3'���$���G~V�h׹�p�
.�M��(�@���7Qw�G�0���,�����r�@w���=�4<�p�ca1^Ǌ��$%�;U�ͨ L6�}��{n�!��C�y�"{�@2Xɇ����K��3r� �`J�����\P4��N��X��oz�Q��>�?��J�-�j0pP����@��e>�:�l�G�:ɋh#_ls���﹨�Vj�\l�p\-Ľ�X�=����C3g �����!�S�+���C��2�~�ι�L�#OB[�h�f_y(���M2<����_�O�a��%�)9AΛ�[ș9�������*��xKS}���G��,4De9��=�c����c4W^)�հzM��j�&?��E�$�5��q��ܺ�x@А�Ю�#0�V����Z�!2 ��9+fe��8�����m'���$�,l�Y�~6���H��=����x��(qI2D�}^5����9��>�0j���X@�Nq~N�m���z�!����䪾�OeQ	� ,�e}���u�:���* D;����@��<����\	�{5�.Mk���⹉!�����A�o1ܩ��w:A�a��$Kd��RR�n�nU?`����rB?}O��]�V8~�*a��F�����k	;Aڡp�#� �mQ)"�����A�B �G�`�y�ѕ��ϸ���3��x�iJꋄ�U��{�;Ⱦ�1�����*<q�zl�Mg�)�A	Pf�6Ur�c���+���t�*xס[�==I�=c��=mU#=v4���,
��f�J����^�����.T:0�q�⭗��,�M����&��t�GsEꫧZ[���]Em�k.Fu����d�M��*����KW���f�Z#�M�ܗ������t;Ȼ^F��l_�G��	��\����q��;�9ts� .l�2N_�~�(1�3�B�2G**4�E�\�y�{I]I��uO�B��5 ���k��/3�8aՕ%	��/���{~j.��d�d�W�s!�O��A�f� ���CVj3v��� �!��.����GSZ��A!	�rRD���/$��wG#�n�lj�[ >��M`7�0��)���F'����P4 �#�Z$�;HN���
&����񧔻˚!����p8���+��0���m�,�h|oS������?�{Ț;
ZF�H��F�^�'�6κ�f�p9�[~q)����A��QL�j�M�����	5ұk�$"�N�P%ς�:9[���c�[�����w;��"�N�I.�Tb���(�o��՝(�ɤ����G�nZ*�>�#����^�詂���<�P�^ya��c��e��̔�H+��6���9���"�%��T�����I�1����/:Q�L�6�J��z�4-5�n�0T��W�#�٘�0+qZ>�J7����<��H���2�F#H�%�Yq�&2��^Z��g�Ҩ�˸�����)�uݒI��g!I��9l��d!z'���$*���>q��$���O�ͦ��j�2؆�ƫ�Ѡ�����נR����/����v
T���ޏ�(̒� G����_(|��-�iy�bhٵ�m(�(H'l���?߈%p#�l��ґط�~����9�;0Zl|9��aQW��	�o���'f�
�c
)�$�~Z�QG���p�"�.�5sVԅ�����ٚ�S�x���*� �V �'���(��L�nUz�ҿ�^]�*n:�B�̽(|bE���5Z�-�w36�k��8W�/'~�fԢ���T򔇠b�s2�K��>�gC�� �=}��&��+����1*��[�ެZu����w?���t��~��/;�a�q�LĴ�N��-���>s���R��Cڽ�TWJ䰏8z�Ң_�IokKf{3U!n����8'X��/�uW�O�`s�'2{`��o��{�U���^$�\���.����hH3-�,����|A0�V�����q�柍t�Y�j��|�
;t�g6����E�TFi��j����o}l1E"5��5�ǒ����J��$Eb��RI����TJJ���n�ϯ���YČ�2�ph�s����ǡ��8��\o�z��tU���0Z����� #�G�{Dێر{50�)��3o�g�:Ȑ�<Q<#���<�ܸ9��!����Qǁ-�Aj��Z�ط���$�$}�>ys��ޱ�]~x&��ם7
Vq&���0h����,�i���c�@]-���l)+����b�n��J����ҳUaO��|��g�n#�m�s�td"h̡�O��<B�������@�ɢu�+ʘ�h�̈�ChTq4���H�&H�OX�@E�
 �����@��g-\1sۻ�]���2��+��e��{��y��˩�SZ���B��t�욥��D�i����;b�U�['2���nM�6.� Z� � *%��$̛?��7�vce�4���YInÒ!����;7 �"礥O���?�ŷ���1N]:E��=̈�h��:<��0� ����R ib�U���<W��0�D{�?2��!�&�Fu|�"�A/��d��t��3���b�/;�[M�xl�v`O���w��
�מh������%����Nd��+@��ܖ����ID��D'q���N��%�����-ۤ�V���ɕ����1)���ݴ�n�
�G���ڝ=�S�.��⦖L�(נC�NS��Ooַd�m�.��+�s�6�O���)� � '���9�X<�d�8<_��c� �Sv��]�*���+c�YF�� N��ݻ�Nw���{٥��X�{�n5$@�%�W,=��ќ�ǩVh��o���bR�@#��5�MmkL'tŴi���VpZ�]1�V�)d�u2:����۽O9S`�[�U^ESA{u���C'��W&w�>��㯁;��L���(|nYРKZV倥��Y��s���U���b%L�j���
F�KY�89�_@��t�V��&@�B��Q4H��A��I�NR�Ff!:i�(�8ȊZT�g~�s��}�X�Ѐg�{��q@�D�Z�-������~��_G��
N'�c}�f�{�w�<Ƕo���:��9�=��ùGN ]��J�3�W�������ޣd��#��r�[iĕ#�ݯe.���Է����5p���ʌ/T�`BB��
�/�����6&��OG9���_�b?l�B�ʾ��T~7S}�^ł,�W[��0p�d1���7�Z�ÚlwXf-��4�����MO�z��x�̿f����t6hJNk� ���\��
^q4��7B�g.p-�NA�l���m�\H^����FW�VKo�F]Ȁ�t̕��Q�ß.9j�_�"��?eg�)ЪA$������n�޵	�)9��:��w����_jэ/�jB�y�C�@��dg�z*�{�^|֦��1b��h� ��"�Hb��N�0�X8��p��~�D��*g�}��ٕw�� _���l��*~���5���p@�2���8�H%��}�TŊ�;1�����%C��T�K��S���fl5Wv��5���B���4nb�̛&����k�:X�5��q����'��'��"=��(n���-��K��)չ�D\��?7�5f�L�H#Fg�^w:�&�ӕ #�Al��d�ei��WN�g�����_"���g��M1�Vʑ�˕���@�W���e2� ���׾����$�'S0�wIM`i���AJ�6�L��n�]V�2�8������<)���r_4��߶��x>s�;�>2�P�3r	���as\ԕ'9U�����)a�h"��Z>.��e�l���ʻPW=�q�eXɾ��W����UwH��3��:�<U|N߄��f}e�g�ZGwC��VןG$����!��C�����ka��v@�7ڽ�Aا�����m��P���|�ԓN��6��l����w���c{W�7A�=Nݎ�X�����B ��p���:J�4�hW������K���Ru"�P,@H'��o!hl�����PЄ9��\>���\��*��}�^Ֆ7�0Jv.m�Aת�>�����R� >B�1J~.��N���V6{tW�}�̃�5�x��nwO �'x����:��tS��8����3�ԩ�._��!���5�(������e������٪�/X-/������ʲ�M�Tڿ�Ӵ�]�Gy�︚L
��ӛ9
����v֨�����r)C�K�E�����Eڏ�	���\�)�F��.U�"-D��Ρ,�Ơ�p��N
ӣLE(�7S�|���y������ii��>� �ʶ��cW[��{���Sw�wY��0�ȸ|:�(P�k������ۺ���5;����E</uk����u�Yj3��<�����a�c�_G�֏��A�`�)PzJ�"3w���e�����V%%&��J�=� ���ý�lX6	��e����L|_^ޗ���$�-�h���Ľ��j���O� ڡ^�
A��m��Ii�d�/D��k �`'���K�gOF�q�ghF�gŢ�֚�0/=F���:�Ⱦ[�4`DBbl�T��4��MCyT�{"�ɓh�3g����h�1��'|�Q��ш��Z?Tmr<��.=}~]F\�y��̻[`Hy*D����/fm:�v��h��};h�j���*��َ��|ځB-uDm�x�y�;���Z�]�nb���%�U��싨m	���?׻���)��ԭ�YHx�c���%l�F9��Y����[OKɒ��r���.��W�L��h�;���W���Ȭ�ˮ,�$c�][�wL�<A��=��H��]����c��s����gS��A����wȴ�Mݥ�0�0&D|�k��	ָ�j6����-������@�˯�I
�W�~��&�)�\�ʗM�ie �a�}RJ7�!��֝�&y����UX��o^NGI6�1R0�c[r�>��cӏ��S�4g�RFfI���æ��r�?jP��NU3�v�`'(��C��N^�}�ԴLu�i9�@���*GN6���Y�`�'w��ɾEh�J
]=��O��N�C�˭�a�a�VN�4JJ&�o��r��A��]�ē��r)RE�Pi��v��kN��[8�P �
!U�՘ҥW����ր�O!�����hr��֧,�{��Wg}劥��M����	C~�+���&�1!�a��ŷ9PV'��Γ��|��CIzzW��Y�3V�)	��2� >����۳6�cf�E�������ͪwӆ���obMBK�2$�!���>^uf����C-o	�z�YC`:�.�l!Y�߱��kJt�d��N�O���!ĎOZ �K�n�|O����(�"FW�Q2��D�k��;g���[������C�j�\�i��ѿ�θF��D#ٔ}�ǖ3��.��LM�c�d�N��[hP(
7h\�ɦ�q,fv�u	������;��I��W�і����*��wh�[�	�I�"�4l��ѩ��~�jrG>�zx�H?�ΜM��K,Y�����p@�9慨�G������j���܆�2���X��8
Eb�S�\��%��b�P�A�qq��{t]����h垴Ķ�R�(U���@���|q� 3�᳣�\m��C�T�x���u:���e5�I/�<�e�1�a�T�U,'��H�fBn=x�E���ٱ��{b���t4@������?�"���(�q��ٜp[v7\��<��u �+.���-���fz���cr�Z��,���Pۯ�,v��'�#zQ�w�ޫk��cv�4,����gB���'!)Z��oc2��a1]H�YJ�z�� ��z����ۖXβ�0�����P�IH���S18�r��t�4�Ր�[0�d��v]?[��+c4\1u�3�#LN/&-n������q����E~�ej��<>Y�/Wo��;��!/|z��f�ҎVK@5KP��׼9��1ͱa];��\K�W���%����:����K'����lN�7���Y�Z�����^5*��^؂�ܒ��2�tI�3���m:�!�a=�K��K,aK�ޯ-xv�F�*��>�p�}!�QɽM�S&&�8+Lv�h��Ma�G����*Y<;�v����5�izoDYeZ^��
��挬�w���-t�x���o(��	A;�By�J���>f	}��`"�fKeqc��+:X�vr3������O�^��1�_�ю>�;'ޣ>I��>������͒/��Y�c�'��[�(8f�q��L�Q��Y1�+��.]�]4�B����n-I�f�XM�%D��`�,�
�Iν #Y�F�t��n��%F�ӭ����[c�(s�q�� v2OY�е&s��ȣ?��a9V�p�cQ1�Z���A���w;�C�[v;�'$XS��۴w�Ɣ��g�\cc�ȏ~���kXL��&[~."W=���� !v�q�F���2Q� Y��Y���grD�!�kɘ�s�6�s�w�N�ZET��Iej��8�R����1��O�������/1�F}�wId���i���@��͓źX��i�U &v���<b� /J�09�ݨ�X� �������ƪp�6�>o�̉��p��yF�<ʀ���yUx.>e�yI��Ct�F��"AVe�_n`�����q���˜o���P+7Ѣɾ'��ȡjr�c��>p�6��:`y�z�?݉Ν�H���P�lF5:�/${9�r�נ����X��t��?QR@vMP�1�<�'��ѣ�+��Z�`>�mf���l���W|��6�׿@�mX�)�z=IU%�iE&��ԙE׷�����*O����J�������V܀U�7�������{����IXO	�3����%/���~���L������u��1��%�	�<�`̦�B�u��N}��ӲX��<0$���TZM���u(7��?	��c&���s�,� ��ʄ��G���2R�F$Q�j�^]e����U�"����`�1
4b)EJb�!�+�|7��� OL�����WtM�	��b�R��?���l�ڥsē!;[�U��`:�|���8p�||��v��)�qk]��kg���� ���ABe����G=��8�C��U)*`/O�#_�Ő`t>��d_�O��g�`=��9ı�Zd���`="Uڥ�Js�#���q�����<�Pz������)U/ᤙHH8�c��Z��u��d����M~�Q���`��� RQg�&��/�6$!������I_fc�/�} ϥc�zk6�'��\i��HBg84���H��n-�-�ۓ������S�w��nGĐ)��J߰��։+��;Уr��q�G9�#K$�&�=)���mJ�w���5�D�b�+D�[����sE8�ŤK��ȝ�ځ4=	�E��c@5\voW��̓���V�����T�D`�ٔn�ǹ��X�D����`X#=��_k�)��4V��2 W�C-{�I
��O;�q?��\M5�����KߋW�f'/�Xȭ�7�i�A*���؏]�I�g���t�7���cy���L�-963���lL�£9%�����m�&' �@�U����oR�B%4�AU~��N��F��1�(U��Ľ�G�
o[�S|��� "��I�?�P��_���#={挣���H}+��9מ$��T�ֻ�	�8���
|�&��?��V��m��ׅ=�eG� V�L_�G�Թ<dÌ�ݣ��Mo��P�U"�wAyUHV2����}�x�ܘ�k��Cz��u�o��a�@��M#j�����U��)(����6�����}jNj�Иa�w��U���`U�A;��8Q��:��Bc��I^%�����<���4��v��N���*��4K��67�n�zb�dM�.� �~�}Lh�r� 6|��av�N�k�㎒�n�Q����5Ȇp�V#w�l^�=�����rx��j<fX��=$�G���Ϳ�A;�Y�1�s���Vž��$c��s[TZ��-s���S"/�o��Y''��i@�UE����[��9�W?�Nx�\{�3�����΄-��ѵM�}A8hh�$b�n����dF�z�TN��1^*�
�e�h��m�u�%���8���mh ��_�:�LY#����[ٛ�J�/��r�`���M+�̱j_��U���nj�(5Vh\��B%�Y���
�Zo>�����c�WE�c�ϧ,������t���:,��y��6��V9�����\��u<�Y��-�Z?�̒1D��v��f�1|��X�s�i\ �cM�E��bx�x`�s���W�����y8�-q�w�f,)h�ـ������\7A��pP�u�������z�,#F����dG㳥ɲ�u�\ŉ��5��=�e9)B�v�D��o%ͻ^�&"8���������+t�7��p��2���Xy*�6�Ō�]W@5g䙉嘇�p��o�]FmRk�q�V3t�����������?�!F�F ��X�,�P�.>
ؗ`�K�z��@��f�{�A�e` ,������͆�T,7��MA��[��0ֽ��wN�E�p�-_�Z;b�o],�{&<���.��w���(+������mr�� ����ȓ�f:�m�#U��UzO��F�3ޭ�U�����B�!���p�V����c|����6A���������(����[Dc�Y��l�Ó+nh�R�b��o�g�ZD�v^�b;�\>�nl��WGp�������|h�>Ȃ��#�>��ty�����w�$�@
���|[�.��D�:����h�,E$���z� ?���>i�R=�EC��U��g�9v7�=�����&ǉ�H����5عS([9����dP�2%͌�-Y	q��Y��*�
�#D�13{VO�i�,'��KTKq��#����,R�@Z�ǿ��ꩪ�UJP2�I���!+j6�8Mϋ�cT)Y�]�v��� d����(���+śh�Ydv�?*��
�e�!=�͗B|����|ñCA�;.�3� ����.2�����
Y��S~��0�>.���e?�2ą��18�l�M(R�R���!��Z�j��f�8 ��E���/9�]�bu֪DC<m?��U�ro��z��8�"0���u/�3����Ђ��ھ�l|
��6*7�{�����L��qЩ��W��MD)�Xh���\��Q��ePkL`*�(>�U1�^�+�@�D�վK�R�|B/�N`9�!��C�����	e���s�8��)t?�Y���-���POQ��������,��`?�o?XEmj�*H���ۣ�4w����m�>w�f-�� ,`�<�*0wщ+AP������p�F]2�w,e�N�[�x�!�9oy�Ft�P��Kҧ��{�wzUvH�k//�yc�V�Ki��᳧q.�k@mqe�V��Uv��cϟ��#�Sح�B1�R@�>ʛ�7�`ӌ�kƺ������t�@w
����9���|oّ�*xq�=�H��<7����n��(O#8�|�����0�W���Xq��x��>��Jn�8iK%Ѡ9�!��6�W�r�n�`"�b!gױIkH������82��;#䰟���*�O�G�"i6�y�� �p�q9qI+4��N���Vݱ�fQ`���>��z3�Ff��x�9��&�QZ�ڀ�����A��?u��%B�������Q�É<L��f`�����7[%��?#�o�p���3�APj��~��S�2����;〴�^�e��J~#O�M�iN����{|�Zɵ͌�fʍ24w-N~0/�.B����Χ;Y��O#��p�[��� �U�ժut�~�U*C<�P3i:,����Jgk:?�Q�(v���@=�
��d���mqp::�v���
~�z�C%��'�]������!ɼ��GG�G#��RKb'~H�~�Y�W�	46���\�v:w���S�����V3��-���\�Z��H���-Y��H�c_a�u�����Ns���@[�_Qϱ�2�X1'��#{��J���_z�$�HL�v�ݦc�Fw�T>�i����醻�s� �v� ��U9+���X�
�6$&�a����ʞ��`U�,eN�w������[��N��"��QGe���t�f�8ho8�bg�\�I�[-�~�G�H\��]}�Z--s�;@{\�2�1�\�	ۜ�,_7�$I��\,�	�5���Ⲇl��tU!�sk/E�u����J9�������:Eh8XQ�r^6v�����A�'�	Oh� ���~\w4}ݕpЉ��tu]��-�!�v��5.�di�����fJ�����~�~�o�$�ZL�d�P�-�N0y=�Kʥ�<�t�[9�J�SR�&6��b�s�L;Y O��_RTc��+��	Ar�*����'�g�G-�$���A���7��ׇ�T�CA䋅�b�ց�W�<u)�R�Qfp��5�v�SrI|��.@���oM#���'�هr�U���m]h!��vvz%qJ�pꐄ��'_���j���+1����1�rJ���jՙ
�e4n�ն��0�yN)Eg�Ϥ`D����]_��cF9�b��b&Ŀ��S�]��>�Y�������o�SB�
V���=����*�=�*]a�����3X��V�,=�T;�������}H��@�ie>b��B`#�m�Rί��~��g��2��S�
��t�j)�5���J�e��t;�~��EU�c�%��OcX�u�M�(����@�E�t��9�˞V����� )�F�zģ�n���v�ϗ�:�����#5�u��j��0�����/� �7NH@B��WC�r*v��%��͛��Ms;HQ��~ߨ.�{Y�����E�/[M_�"/���BU"�.��uðKsT*ՠ��1W��	�(L�F�W�8����8
�1�Ԃ�+��Rx��V����{�ݔҫ`�'�5��^J��"���E���[fNs!��D��e�1�$���lh��E�P:d�X�#�;�K���YO�8~�A���Z�x��Cq��x��Й��;��-3�s��!B�	ޚ�( ��_�E�Yq'se+�Wb�օ�x,������B�*H��"��ɩpA�ln�|g��[��9�1�0�6�7���xE��ץE��4NU$�#G\`#=uH��0�}�� O�N�tۤh����_�����ـn��мl�$��=ж��o�.)q5&����K�ֽ�X�y���t�b,he��0i���{Q��&B���5�50�vTd��Z|�Q�K೗%F��}�_� 팑`��]nS�G=��n'����s7s���b	�Ib/[B��sꭷkj�	ð\v԰s}\RLH\5__z.ϷȚ�q7�vS�M���Ҥ��(p�1���uHA�����^��v{�SxD���e��n>
}��}��= CG�=ɴ��-��G�E��F���4�=�	�L��(Sjil���{��T�80�0������<���Q�����#����gW�/fZ4�Ev�$��e��/O�Ǎ3�Zxx�� )t�	�M����:A4�B�x��$on�8,aT�¸�z�&��i�2[�]4^U+����+�[�r�T�,�J����1�M�	.��+�4�æ��	X[��|[1\Bt�H�����
*�vV멭�F"�}}��[���C�V\ v[| ��]�_�6.T�GNT����z�N����}A�7��J�L�@��9�3	.Ѐ��Cz>G�Ƶ���wJ��5����)T@z��Y�����l4LZXN�ŧv�H-:w1n�c�5��D�iA��x��Az�JMh��!�}`��!�&�M�\����7����V�R��U0	Y�.ѳ�8���8'6W��KPȿ67��-���\�x���]� �}}�%�������va$�lf��Z�4�h��u�-��(�f�O�|�Q@���#N{�i����v���� Z�뛊��Eoz�k�=���r�b��4��ֽD�7ͫ��5w�3����/�X^��H��A�h�],e�"�O}���ť���^�w^%̘렛h87���c��	4�r�T��O��}!!f��6��K|��z����q�;H�<�����B�C��I��V�~ψ�,��k)!+쯊���LCՠSL�1�&y#Y@��݈u� r1��-���HWO�ЋgeG��� >�'�͊�g]Ǎ�x/.�X��J����o�z�u�U�|��?4)��Զހ����!�����S�m�5h&�ik�q>�<�ؗ���S���#�Ֆ�󠟒��1�k�2�i�:-���1}����J�R}}�:�((���E�[�g�y�*�O���pmy�k�\�Mҳ�>��؍X�=�A��A�8�N|�K�&C4���ߧq��n呿�ۊ�K�\����=ޅ-�t���|� ����]��Z�|c���t@�c�w �Zo ^|���̥"�A�/u��������gC!�0v2�V!�*ꪌ�̸t8u����3O�> Ժ�{56���DJ��N�>>bJVJ�@���v���6�,Ԕ����S�a�C���~.�.ぎwGƾ���6���p^��e�@��Ml?�q���M���Ϥ���d`��LV�E�b���o60]�ŉ��6�T�z!n���ٳ�����U��aIP��ߨ�=x��m[��%�=�����ra��ŕ �
<8�z�=���c�/׾iDMA\�J>�Vs�Q�	�O���UE��5�	�wN��4�\���KRAlw=�*T���Fy�g���ڳ����j/�t#��X�T���:=���\�\{�(�D��5����蘉 _���?�8���>b5w��g�j�K��r�` �*����k������gzP�������� �cc����2�]�C�����Y�1!N��r�/�����͊�)?9����'[����bM��Ą	�p�v�����t��qΤ��p�*��$�@�^�!%0u�r��a�H��6����r�0�zP�,��:CK��%6a���򮁬H\q!�.�}ܽ�L��V���A��7�ʿ�d6�\��Wƌ[�K�.�Yo���}3�Y�XiL�er5g��McU��X��I��o=:4.t�r-9GWT�3��XC� !~��6������V0޴"Ǣ̶�A�!�ŕy�p5�)?������&`@1mo�%�RX�+�����*�-,��1��-/��O�(l�ƺa��wH�ɠ/�RR�%�(�3��1/̀9��4fl�8����.K6mƬs9��x�d�*�7�o#�r�y�����nN��&U���Kz5n<o�p �	HZ~�x�z�'#Q^r��m���_��O���=��-�'<�-�wT]����[��hn�����zJ�$F�Z���dYٿ0,G��ֹ*Q|7-�H������}�dצVռ�-�bE��w��nH-��Q�o�,\��q���eJ�1�v�Z�E� �7�Wl�\����&�
BaB~�'z�8�n֍C��Cg]6��E��v�p��'�gM�Y0�O7��Ξ�oN6	��A!�h�Ut����+��ɶƻ:�l7�p���~�)x�kD�;+�~Rg RQ=㫱�Ң'؟�^q��A��Wܣ����thB(�\7��KU+XBZ�+z"y"Ͻ{�;��~x;/��Kt������,�y��W7�V{.�C�ۏ)�O��e3}Ip|§5Sh$-TR�2I��D>P^s�����o1y�������h��W=ތ�7�9Hؼ�A��-�~�n�}�v�qz!�.�jN����j-Ͽ`�c0\+�0��:��7�}��
�2l��g-�E>P'4�#��Q�G��C*��(� Y���ĝ��֗E��~(�1��]1<�v��χ�����C���pt�w��:�K����_(3�!���Z�����Z=��v-���8H����z��w��之O(5�K�l�A�վ����s�=���L�S��*v���J��P�@�Dr{������j&�G/�"=m�(/�1z~ �˨h�[��	P�S(�q��0���\fU$����4�,�J�N�Џ�j��0hY����0�<ٮ�tL�J�S�"#�ff�����Q>�W'���᲋���j�ܰ��.���A]�Ḣ���>�*FT�{�7`Y��Ӆ-����?�}�Jݝ%�<s����G�:y�˨�8x>o9�3�̕*��t��sr��)ne��/#lWϸ�,��j�(!�}��R�l��qn�.v��([�ӣND
}<uݗ���4i这��h?H��^��*�l{ �F{�4��P���%Y���%��b��noӔ�G�M���1
è<��W9��h�+���AW�L��l��h��嫏�:���7C�r_}�M��7��V��4�����&��[�9�#������'s���&�i�>�l��������\ܠ��ztW>��i
/�;�e�	�ǩ��w1KN��bИ~��Y1�P:i+�g�&��@��R��V*m��l�uO��r�\B
b�^y؃Xm����D��h}��-Ip=��@?��j@�?۬��:�m�5\P�<��T���|rw�E'(��ӝ�gI�J�R���<��k �e~��K���li�2�Y=�ł+y����z.#K �=b�=�3#����V_:gY4Sj܊N�$��.�:7���A��s�������g�<{�cZ΅�\�(W����:3�zx�~%c����4'G���׬�^��>�I�Lw:@�(�F����i� ����l���R8����T�[���t4J���@�oBXYY5����q))�	텚ͼ/VCX���F��a�>�$ࢌ9B~��VS3?Lo��f����=5��=��o����S-��0L�o}���z0S��}����i$�VTgz6$%��b\R��M��f'?}��Ӳ�1nl�%�s��a��:MR���ѐ�6�I�#w���Z��i�s�4�8Sx:��ڢz��)��J�D�:�+�#����Gfˈ��'&��1ț��<C��ts�Y���s�����Gq���f%(M�.���$���ǖ>:�F����L �����F18<�3�����n���X�l ��n��G��,�*Ol��~��H�.��!�{\2��Bw�R�W:�#�T��?���u�ұ1����91y�K[ Q��Ab���)�K?�L��s�����sLoC����^"�Ԩ��rk�Gv��'[�`ʩ�n�mh�։s�P�4����������r[8�De�R%1�SҲ�x�V6�iCI�6�o�)������B��q�BC����{>����_o�=v|�� ��ux�_�X��J)�~4�i�a�v��7��9���u�,7� ��I�F��n��С��x������j���L\�I�tuC2� b;�R�y60�b_�US[�6��7�2�LCzх=�^
�C�e��Q6�U�����By1���D������j���L�[1P��4�Z^���=ۂٗ6��z_O����H�L�%��5�RD�b"(�<��J��n���36D��̜1/~X�p�����a?��o(qfyV������&�|�&���)�%����x���]��t���K"�{+�cRZRז���5v�n�Z	.b�p�?H����-�����	��ލ���߂,#t1��W��5�k@��#�)k��i�ե��_p�݁���g~��m!#����bR�S��rp�1�Af)�7�_t�L"X�O��	�{ܰ�����v��gP��p�t⛜ْ�dylp�e[5��j�+4��=���Ɠ@ϔ�Ŗ<�n!o��W�mmiI.�W/ȃ��s.>��K�HE�!R��3V�H]Y<��4�*�H������	�q�R�{E���J� �V8ߖ~�w5Cp���ܠ����*`�(7�#���׬�0?Q��#͜��bD�UԪaBH����RҬtk��JSL�iu?�:�t��A����[Ak'`��G{Y#Y������O�ȼ��i��;����q�"�(�� �LLR���Vf�Rw��\&=68��D`~�+�,��R�-|f!xVR��8��u��kY��RQwC2�5�j��� Q(5��6:)�}����L߁h���IF~LB.���=����yս}��`I-�NVsӵ�h.m�o/�JK
{A�J}`?ZE�ʽ��j�j�jCP��:�=�f�+�����]Ʊ��%�� �!���>G%=�vYC�אL1_-�/챔p#�������9�8��P��rxB�HooV\h�oF�Vx��� �H��@�V��:�t�eL��,���Rf旴4}��)�_T�ʺL�\H��f�~��<o�5"�=˲
��s�����5GT�Kvp')��kϱ��L���m����� <^я.�r�ӛb�@���"_�$LVE���L�#�QAk�GS)&q�S�����zt�'�$��[���YI �؋�G{i]β���毊R|HG��@<h���(#�\���t���%L����Su�XIc(�	�F�L�<�F@��u!sQ�2�<3��3�m>�<0����f\�5�7IMH��٩���L�
���zB��U�R�'��0hə_�	6�P���0��	���pͯӢ��s��Ȼ'�2���i�An���ӽ�~��MVG� �R����{w�U��	�V�q�T�Z�(M�j�E��e���A�<���$ J�-=	u}&Է�r�R�z��H�6 <E�z���b��\�.�Af���ԉ���"����C[f=
�����(���nP����G��O#�t�h�rm���:�{0���1�;[�~��Oʼ�T�^%Bev�|����gY���}��1z�|�r
W(�8�
�`�}�au�p���ޚ�oٴ�9[3�2���z�O4�1����cÙ�=��������[�@K3�m㬏ߜ4�K~��6a���%�,1�X�]�[q�Ɛ�3�1�0�%i�i��|}$R�]d�������i����Rl��>u�V� �<��ϛ_�J�'A��.K�0ò+�K<�R���h�������y#����WN����%��~�$�RW�`=s�k.�|��IV/���&�	�B�@q��yQF�Q%�&N��d~b�q�2)���&���o���*�d=N0��1*��.7c�~��N	�P��Wo�����[#�m5U�݆&>�I�A����fȔfܵ?2OFN%o��:�!ft��NRn��F�/J��J倲��93l�����7.4����b9w�J=P^$؜M��L��LFv�;=�D�H� �iB�5sK�ʔ�'����ݎ���S�K-���˼�IE���>���Kf�>�,2m�G�/ts�V� �� j,҆+��k!Q�k�Ć0�� TczR䛆�8���2�k��Nv�s��By�:Y�kuZ��k���䴽μ��������J5��>�z�w��aa��2f8m�V�VA��u�F��n^�V��lֳ�߫�e�_�R���m'�w3�?N��w�a���g�u[�H�i��>���$O#'���M_��vȣ��T7����Y�'^��ɪN�fn2Q�^y(b�]�b�斮sۉ�"���jpz'�s���b#N<���c:�����ݠ5ƇU�B��lg� �^?y@��N^�Ҡ��i�/A��Ar�<�e��U�%w�a$�9Y�؇��,�`�.%]Y��qxNy�ɑѵ�o(ր������K�[�I���z��JF���'WZ�w1�@s�%��G���۴ȵ7�/�x���C��6g&_�>��~�P��'cT��dmlWw:pA�}o@����d[ډpaO;�m8�ߙ/JIm{��}&��v�E�#��ɾo�>���&��ϡ�j*�O��i2G��\/�"��͔j:.5J�e����#G~]�D5&g��oG�e�CW�|N�?����M��ۦ�v�O� $�<����1��|k�x=�ȈaȄ-�{���[G%V����ol�倝�!f�h���-�L��M��.J��m���*�D[�C��l�\�|}!�D��M��*�e@�y$����!l�`�$�EѪ�;�=��>c��-1vf����۰���@s��z�5� ��܀�~��{J7�k�� .w7fAG���"�3oNKmD��c���J^o\\��g.��#�w?i�}������' r��\ìwI�f��00�v�@�4�����?��DK���%�����^����s�G)s��},]�9O:�Ĝ�I_��N��c���59.���=7^(!�-)�e�h��p��A���LKـ����-f}���Y.��H��� !��y���8Ă�<�!�n�؜��>���6䜴V���H��SY����!��Le�Շ�Ƣ�LҀZ��(0�X�����g{a�v���k_�����jbR�g������>iY;j~={��9�ՙ��^Ǐ� ��p���!��ӑO�67Y�/��P��=�W!f#�va�á���!�+�v�	K�,�>�߷Ӳŗ�����?{c*�3O���4�C�{���.6��7�	J�!�ҏ�y�Kl��)� /�J��}��
���29�DOA��W_WC#Ma�s� �1R����;�b]�M�
���E$���v��<-��F\R��݅:u�t��[����۟wQ���%r��8W�����1�,L��K���mZ�Opr�Ql��O�E>JJ�͌��N�L�~2~���ψ�o!�p�}�o��j��#�8�c��Iq�Y�$-7	�KM.�0���s��tC륑5��_�� O����&��"�ؿ�g͆�
�z���H��.�o͂kMv���dN����(W.�U3�8P��:�$ݱ�:�����Ej�wE�e�#U�.��d�*q�,����k�5���� |�@�c�c�?� ��ˁ��g��QV�T=@��R ��1���9���� �JF���験�l�Z��!8w��$A c�ߎ��x2|� ���IΘ���'��䂽�o�q��Cb^Z�����}ƻ�v���q�Xf� ���i�lO�+��=#�*��>$�[L��G�'�\a�û�Ѣ����(��1�#d�Zz�mi'HT�y"T�H�:ч)1�K�a|B]$�_��	��.++���Jm�P�x��-m���q�bt$�����<�/����d���)���e5GתcM�FYwd���O���u6׹�e���h�y&A����)	����#j��8�zBqFߤ�K*�xO�>���lf�������������$�?;��@�#�[C��J5@|L���q� �*R�M@�=�U��[�'y}x~�0�I����Ad-S���j����p������B���9��5h.aJg�8M?�4��Gm�	k��B"s�llS.,�\?�l�B����>U�ei��ô�{�܎��Z<!0���hs�2�3xv ���-�n6b
{?٭�K&�QÑ�+��CG��P��m�AT��6a8v�u�6�4�M��x�߾���2�����3�y(���������C�sa����k�,�0��r��(���C�u� �"4׷0��r��-�vr?�2�%R�U}�3�Q��G6�\tJ�x .��a�6ٙ��RS����Q��&��#����XR�r�iG�9�1-��<^�pP�w��'� cM�Y�X��еTRv����
���ʁ�FD	��j�3��g�4<��}��W�/�Q�S�g�MOe�1��ݐ��ix�6��1	b�6W��xo[�#e���Z98Ǆ�;�������Lj�x��/s�I��?:���j��y�.R�T��M�#*��1T ���i��N9��E�����hY���tM�R&�V�Ӫ胺�A�ay0�"Тc��iy7������'��Cr,bW����Z��mw���\��z�o?P���+<JZ����u����`�i ��������(�˞�*̸�Ϧ�t��r�L��м�j�&�oM�'-�Y�S���V6o��o�[(�����'�+��P M� 'b$�"H�?�[��#�pn�G��&��{6�P?�9�+맅�?�T����O��������R��� ��7t.�5����C=#*g����YmY�w��K��1[.L����}���5�W�7��'_��S��-Ǉ��3d��*#k٢��Vڱd��A��%�,��;7��]���WG�`�7V��G�'��0C��Ի6/��k��ڗ��&4��I�*�-z>�y ����H�,��dkb����V���O��Օ��KR����%�V�ĩ�IR�[>�õ�� ���Ju[�H�:E�R�q�Q �x�P���S��{a�
b���&o/qaJ޹�jO��6^9�t�4H�z��3Uq��,��g��콥��OZO�\�0�vF�&j�ŕ��i W�,�d���U��V2R4`��|�xt.�ǋ��X���T�"�Բ����6TDհ\�f�<rQ�vr̅)�>���_�s�Y�
�z��w4�k��5��
`��I�2��rǪ�K�X�WP��4W��v��w�i:	�7OL�w�-g6	��]�I�ʶ\�I�O~#4A���m`5O�*�߲0iHXG��|v��E�(`�{!_0.�{�I|1�}~��&�ǋ�ĪȬ��V�f�s@G���FB͒\�Q�㽍]4.��]v���}�	.�B.�"k���0�wH�o8â�ā�����F0z�ګ�E����M����^�ڎNr��(�jh�E�s'΀_��ӽ�GR�L�Z��~\�������?s��~��p���Y�!��h'��0� D��(�\��dd��1'|a���A(�w�0���69�b��SV�E�����7qv�w�@sCZh�K�UYW�-��/��&�}�na���*�.���|ڜ�֝�,%>O�5�C��-oV���U�~�^�KgϤ��������wg%Gf���zLE�w��\�x��$�k)�j���&ď$<���A�ژ���U��`:O�]�D��%�S]���֌�ɟ���2��`'��Q(t�U��am�]%��p����+\q<C	�"��-=�+���h#�8Z�_���p_������0�����=rO��vh�9�}o߫	n7pb��?F��:��<ي��/��|����5�&+Ues�{���6�t2
At�&-q���k��总��w��F>��.*x�>��憎�p-,&������&/��&H_��g�t�͈k,�>���<
'"�$��y�7o��.�#� ����"���L?Q���5� �aJg;dH[1��cE��T��D�NW���ퟰm]h"��$��qu��?EF�F%���6m�蓔OJ�ދv����$��J�|��Z䠜�U��9 ��pa�Y�����,������+���WY���?�д���Q����J���g�\R���Œt�m�͚�Ηr�3�[�����zY��ܳeY��?<���W�'P�ڛU �&����=L�zIeuk��;�ڏ}��2��(\�QSj�Է ]�p� ك�/n���J��j�;�a�{^9I��h&0�R�b!������h�D���{�0Q�8T��X!��(mYy�i �1����*����	�U�~{�rԦ?5S�)x�S;��@���C+WS�\�J'orHw�@)��ZO��壄H���i��y�o!���� ��!HM�'p�U���G��Ѯc��ٴj�窴
�Il���1>��h�m'T��PN�VC������Wg�@�P��{>4>��l#m�Z	�xPs@�"��q/٭� ��=T��ΛI���_�1�Zhz���R�`�k ���l��ҝ[ߴ��i�g�N��qc�k<(�s�����Y�/I*��+�[�7��y�ޓ,�=7@�{8�ф�<s�`��:+�hz���SĒ�Oۗ;ֽO*~�ͺ��@������݇I�S���ҧ��6�t�;�
(�� ���T��K�a`��!7������e2��_� A{8n.�ȾǹR]�C9�[�ANxxkhoG1rn�� ������2r�>�!NRv�9��%��g~VB�A�̀P��P<�0���kfq ޾���{�떉;[����>��H%t��U��;�U��ZD�.&l�X}O�N0��=�F�v�	�����[^��&2�N9c�g�!pwO��x�;u�	���9��"nzQ�O�M%KZ+o��}��{�+-�~^���S���?�Q|	�J�Cq�������.#J@h��VLl��_��B�zk'�mq�H��@��6IDy-�|��F�O����ڊ~v�dm<x�pa�&���?���Kr��˓"��Ds��#+�
�уqEEcJԟ�W��wo�F�˒��#<�~��H)���/F�l)$_�&׆7�-��cAZ�l5�{�����S��p���81Ͻ������.�L]J/���@8��t*����j0%1'�Â����Z�Py�Q��'���v�˶���.� *�fD�7�V�E�vr��/�+��K_����
�>�m5}u���=��F��[Y��څ�|ڶ!u�$���^���/p��Sk���Z���ڽ�%99\dx�zP��"�9�Kׂ��-��|���0.�/}{���tb����>�[ Ү�w҃��?�1 �T��M,"�Oܘ�E	��������:,�:l�'2$5��&���y-ꡁ�2��~���?�=|Zgz��5A�S�Y��z���������u6g�Fʐ����
N���� /��ޏ��dy�Į��)����.e>�,kb�z]Ѽ�&��V5�\Lt�̋��:c�R�hC�����m���M�������곮��yx?�ϰ^�gi�%�@��<	[�Gܐ��8�,�c�<~u�H�TaN ]��;,Ԁ��7\K~&��W�s����@��=������]m�f-�zq�Qfz�gR���Y��&(U�E�p��>��(�F<S�ԏy&{�' ��S<�� [�#R��}�5k���O�
�
沑C�3�;OE Z-�}�+5��H��)1Čz-8K�E�6ds#��h/+�u�nT�Я��-ٝ��7Qs��U�"��T�]]��m�ͩ� p�AJ��;(c��v+�S��u#�Gm<2%����\[:��Ŋ�a�Hn�ڷ��Xzp7U>�q��0򀒨��{�"��� �=ү��7n�N\��]l8���[jY'����ۛʾ����u�<��P����H��*�ύ�*�ر1,�w��שU*��k�s�dG/�j!{�e�ؽf�1?�59����[r	(�aϐwcU}�(-��V�T������]�"}2>�XiĞ�w��ݩ�p���(�Y�k�r�������t��ì"X���.��d�����M���� �t��ȶ�g�9��e��Y��ӏw���֐��o,���t���)����~y�|ǰ�'�`��=L�����e�HxU��sw0aF	�)o�
( �JU�����=�\�D��o=���,�;�Tu�Ns�nv���Q&�z7}�;�	u�=�5�����~|}���=�u����i�\֔�6.�3;�'i�����_��c��B�׺h��+��Nx�z��� ~���xD�{^>�Y�!��3����Xbҍe�Y��y��P+��`a����I��S@���\$���<zA�`ɰ@i0!�
L����ؚ�)��x�xa5�hg�M��ȗ�U���$�;dN̈�.��f�HpDGb^"��sȲ��wF��ދ�:i�g
�)�m0>ebj퀋h�  _��g������%]1y�`��.��I�5LbN�V��v^����ޝ+�"]@��P��i�|���-�)���t�S�|x��I[�"�ϖ�Ć�J[ޣ��o	X��O0Ǜ���z>5^v��i��خ���#���%�*�c��9��pع���-Yy�-x�'��ԣf�t�I�4O�K2Kv�0]&�Є�Z6�X�~����q�×�(��K����+���n08"����r��9$�jXl`f�3-)��Ec ��'�>2$}l�Il��*� ZӅBK��#	g]�%��̀����G�R��1�4˓xm�%��^�'�B��T)�.��F�Ơ	ڜ��+�ɲ>),�dV.��N6lW#��j��U�B<Bb���W��Cʆ0w��*�]� �)N��&�U�]��Q	�a�X���%=�h͜�K$����������x5�<���AǼ�Ŝs�U3J�`� >����WU�[R�2 �. ; 0��\h"��V�I���)��^&��B��۟��q�t�+�����Pe:s+���DXEl�Y���r+�%c�5���ە����h-*�?I���O�{��<V���@�:4�Y]��B
.C��S7������q0��3k_�"���ΐ�G��tۉK�%��:Q�����=����K�\�s0WǛM��m�(T��&��T��*ZI�|O�(�v+�Bk��qS�V'We������0�H����}ם`u��hdX�x�L-���X�$C���kY�#uW-��8�S1�[�0~L���8
|0�wr}�6'��J�6E*��~���%;"3�tve�ܝ����!R��t �C��;�<؊���(a/�Ț7��aZ��z�}��F�rF���A�}�Vd*����Lk�A�ܩ��!��c��F���t?�w���nTL����Z��P�I�<�I!{v/I�<����zg����\�b"?���^9p�M��z�����=��A��2k���Qq��v��QV�%uHӶ�X�	��;3�h�<�c�H兰eI�u��/�(7�?��-�ᦡ��$ɹ��x  �p���� |�,bW#�6�_�A�j����w�?l�@�\�d�A�d��ާ�pyř`���J��%q_4�*-�P��KF�?C��ټ `�Ԡ�HGp�)]N��v &���Z�����ڙ��+��y$�^PK$�Pm}��cS�1'��V�}��g������Q0���*����\R,(G��ȺĮRS		��>km��q��[/Olh��8>�1� �ٴ6Ǝ,���H)�� ���R��ͯ@�}���%������t���S:B�ݼU��!��	����Fĝ��X�Qʣ@6��t��l��W�:2����n�z��b2[&���:��״e���.��fJH���(Wų��
���t��������oX�E����n�p���ҟ���Ē)6���2)���|ײ�:	P�.3�nC����J;�ubCN@�+yz���?�Y�����,����|��4�C�6�dj����}=y4����*��>�3�-o"��C��eYD������#��:�Su�TpVZ���/(�[�������,<��,b�q���]F�(BF��꺊��֐/�i%�.4�T&:�<�r+39q#�g�I�x�O_[ �tϘ#zR\��{�-�)r�׏�ȱ?��I���!#xF��}pVr�.�X�6��-�*��_�r��:H���rA�D
��	=�=6���	�°aM�V7�k��Y`p޳{���z�����g�y5�9�iĢ:�~�?���<ڼ�ɣ�x��/X�}-؂Gdr�2��^�� V�K���sf�SCC�T?�u�7�KR��b��N�z tMq��qW�;���n�9r�s����ޓ���ſ�2�p�W)Z�U��_+�`}m���H_=��a�ۇ�EU���!p�}}�� C���0�+��ag�g����݅H�{�՛
l���;��=;���[3����os� B��x���F2�����ؿ]��O؄���[�	vQL ���w�Bk`N}��:r�(��>vc�P�g��=|����B��iR�O�t̡��p����U�|���-K	���V*oJwʈ{Ue`�qj=���l��n[�|��Z}��S�c2J��@$r;����S�O�>y��D! �U!�����VgkS:��c�� ��'���6c%+vX��o;U�*�s��|$���v�n���f�|�W���c�R�d�(�יICg����O'ђJq��C�]dA ���3�P�������o�6����OI�ogKT�_�O����v��<.�Xn�x PRb���-�r�Xb��Ԍ�z�)�v�0no�z�?#]�����uS������TS�����l6�	��?���tĪA$D�"X<:��D*�-.����͊�b�������`����^tl�y0�s�7��h�C_�E5�Fr����"�	znQ!�{p)�I~��'�=*�d����½"��,�=S;�3f��f�2)OFk�"�V�Ӝ�ڶX	`]������"�ҕ���y
F�/�������NY({��דO-`��v^�m盏Ggw�ez��
,K=����4��lRµh��3��xug�3�*mXr;R?ؘ�׵�w�Z����SŌ�;e�s�9�Y�!&�i7=� ��u�C���heM��u��SN�Y�Q��<����lH�����#�Mz12�(F<���'M;�u�{�l��B��D��u��1���Q��2��k*��0�Y��m���Sre���ÆN�6q��lYR,�(��v�qD�1ה�w��6d	�L�F۔<�!P+}�K���T��p\H�� ��y�aM<ٹy6�K��*��x��.S�P=������%탭ϒ��h��DɊw.��!�/ ��F8)�;Uȶ�7Q��ċ|�8r��B���(��/�X�^O�1���VK��〭U���m���(�>W�ej����o��O%p�OSeuqS�U5I?��o���虊G���e�/+�,9As���&���x5�@f߱��7�o���ٗ�������(i$#>{�;�\9?P�!�fʈ����ޜfc�N���e� �)G{3��̨״�#�?˭m�ͭ?(�"���t���lMU����������F���嫲.-E�Y��<����}�Z�:���1x� �0RT�=C8Lt�כ�6u+Z���qv�F�k|�ՙ�3�@3`{^v�F-�� ��)�᥋Ip�&W���C��������1~�z���9�e��5��~?��F�3q�4�L��1��o�ը�:�v6VEn�5��.�>�*s��_�S����7F����- �/ �T�Ar.aO������1O+��/ke�Qɽ��HS�A,�4�(sT�ᮖB��vVvD�T�ѤcF��"[�����r�;�~X�o�@b�������0#�}�5�EAmc_"o�y`6���kj	S����ػK~,y�f�ҭۢ��{��nq��$OL����DTX3�Kǐ��)���-�����/T��E����t]~�R��-��������<���>d� ���|��FPB��E�Rױ�䰛���gz!� pÝ��n�1x�
L��c��#V����P<W����Wx�7���S�	H��..��.=fH�����V�`[ŊO��`ؘ����]9^Vڳ�C���f�w ���VO)!�����A�8]�0�B��={�$MF��jC�A�^��G���|y���C�E�q�� ����"��W�6-�1ok���|�h�pLU�[	���~5��O�6��X�Q!h3F���c�Q�:u£�����xMu+�s:�5��q�s{�Ni�T{*BtF��d7�Zh�����
i��d"������c��E��rP
Ns=�]#��|iS�
1��.�7�hrO��[\���Huң�ސ��$�݆"���=�А$��c ^�u���  d6��{Qg��t��4�/�r��L��^��2>��ƙo���_�����h'����� �]y~*D	�G���Ѥ�R�^�OQ�>�/�3��%������.���}n1�K�	�&��<�r��3-;X��\�)��Įq%�a���q����0�T��#�fy2U�h3{�P�0� g�0��:�*�F*:������	uÅ�R�NcV-8��D8Z_<���!�.�]B�j+�7-л�}?T�4�/2����o8!�6��R�e����� ��t�Rhu���v�c���� �����>��L��	�9{U��ת�.�rD�*�)9Q�S-�`�X�*��B
��.$x�rN�}U�g���P!�M?V���n�%Yoq�_�QPM�؇L��g��}�w�O*z�c��&>^ڞ�E�6Ќm�g��e�|���V߈�9�C�ga�)j��Zx�)�
��u�f"��W�qGx�~�(�͠���1A��8Vb!�e���b�f̽�M�R��C�7�:����~h��e�.�n�e��X^K�H$-7�o�z_sU��T�p�l��K�jR2����v�b䣝z�?Y��%.9��2x˦�eW��Z:�`��$���s��'*�e��EL�_�U��š��T��!W��'�TRT�#�[~��J�kS�n�Jq�^&�YM��݈�#��V9���V���O�v[Ff��:��%2�"+ew&�&V`:@!A���];�Y�zWu����-0Nw�Pm�)��t����&ɴ�����*]x��q欓����[φ�����x$��
�L�a�-_	�ZW�8?������ENY�u3%!�1�@��t
^d��nEt�>%�i?��Q/z	�7^\��i�m�6�ہ&�Sȷzo�����t�L����X����w謢S�o���b>��;�XB~!����af\���k�=K:�fh����%���� f9��&9��R��p.c(�ns�k��5�����f�$:R����ô9���o�؈�����S���̹����Y��xs���M��v��-�t��~�p��Yg低S�&\9u��M�Q7 ͆業�|�l����)E��~�ь�?o|K;�`��Q�I���������| :����?7w��4H��6���
�u���9/��#P����?��▫xƼo��� ��vLs��0�p�0��1��^4�&�]�,8y·���$�4$TU@�"⏛��gT�5��~��.���*	a�j�S`| �I���_�̓���&�K��k�h/p�x.��ú��D|�>fz�`�.��� I�ƵG�x������K���}���Ǣ�%Q��5���Q�|�(�Wq��T��oQ� �ؙ*X˷E2�TN��'f"��W���dr2���EX�8�R�avu1­��(swK��#��!��o/�k۫�\20ٱ	%��^���&�]�z �eFUL��ӂD�jl�a���6�$����<��S��s���X'aR��j�٭x�� }��+E$��SN�\�n�4~�����L��\A%�Z�l�bp�W��ZU�\rkP�9�`j�Z�e\�ĝ�itW�
i3���c����>��	�s��53%�"��(�2]���a�߃U�f�n'R0Tb��S��Q�{sIWש����k��x^�Q��#�]l��$0f����fw�t�ӛ�c��F/�B,�����u�7�~�=�b�֓�>�ћ�s@6�-��O�gDp�}s��-�N�����NG��$��Phϼ-~��#�P�ܸC��۳GE�����R�5�z�TCZB�uH|� ��\�����q�.7�܅A�ӹ�<��|��,���?�<R����C^v�E5�oq��y��?��H���,�|�J(�sC<%��� w>1��#�ײ�p�
I��HVM2J7��:n���tB]��կ��H����8/�^[K�����t���p�Cd����fZ�@t�u���"��ɷsz�Ƥ�Smߊ�T/���#��)8�ŜX�UDk��ҙfw']��\�y{gk6`��1����W�âۿw�27mW@�,��*\JӍl��`gX�>���Ȏ-��i�Y
zB#x�Q��PIp�����d�K��į2-)�7P��R�| H��[8]�d7�{���*S�A\{{�>ĥ��Q���B�q<�.�ޔ4ߝs�~_�-2x)V��m�xʷ�,T���mB8j%�͇ �%��(`�`�8'
5�!b��4�2ɑ����,�2!�iH���I�1�T��q�݀�Pl��D��9�ɛiE,��ט��<��h8�I+��3��<|���S�Cxm���z�`�K�����>���=�
*B������9��&���d(
��ҙ�ϡ�B
�� �M��5i� 0EGYV�tZ�d�w�{O?+��O(���9��C\
b��6K},����-�����k�4PNy��6>�X'CFKk�#�e�rw�����	� �X��� W�l�`h��YL�sa��A@��}��i������n� ��Yc܄�c�"R�[vtZ��n=���\�7�.Mu�KEbݐS���k�E��ҝ2UGD��j���T������Lh�M�ՏP|�D��D�	�w��c�zB����4w��޹8��@l���X�<�w�̲İ�.4���*|A�h��WN�9mD�٭û�G�'�R��(�|b��(K@�/�r�/�M#��8�z��X۷�[��}�0?57��C� A��-
�x�$,Vq�o	����dY1�FԪS�����:ix˅R���&l�E��xȈ���>�L��E)�%�� F��?�L��I��,�%K�\ァٮL7m����;��![�O�f�A��M7м0uI)���H!*��jB�ҫ�#�J���m��.ա<����[ص��(�c��NV�;�����&��VT��p�}[Ow"�tS��������s!X�%ab�0�ؠ_��k$�z84`����v���D��μ���ğ\���e�R��[� ̥ -�]�[[�ZzbA{�����L���z��z�G��#�Fk@l5��0�:�M�bc����8�����Q�P8�H����H�BBr��d����X:'W
��dg�L���j��$�-���x�r#��S�@���%[�|)���ԺȾF�x,��8�%��_�&���K��e|�������l�>�c�QME����X1!-k��sR9BU����YTQ���)��5{���[h��|5N[�9~X�2�c�~>j�e�#�aX�$#�T���t
�����o��&Q���*�J�11Aȳ1f覷x)K}I� 2.o��Q�����H�9�.�ͼ��j�<���e�w@�m;���Q�{��A��\�ٔg�Tz�[JC�H�A�f��"'�#{�Tg�����pn�Z�kt�ȶ���I�]����H�朼��D_&���Y��{�����$Ò���1�4�\�e�i����?�6
�@Oc@1u|ߨx�[�I�x8T��@DL 5�[ u|�ϊtw$�_�H
�=^�����0O��1���C�)1|��*�dF(�5�卭�4��N�*�z�;}]�� �	�[�W��n�p1�A)�����vvF�7]ۦ!&6���u�6	b�Q�h�{ݍN
���_�4m�<׏��ؗ�Vj�y3qjZ&�k8�>6�">�+l��c����Ť����B@�cЧ|U�8A�i2���+�C-�Ö�708͋��l4n�h��z���m���~�I���^��F����+�u�}�Ux� ��T�u='����H�˞�PD��%�%u	�a���|Vj�(�`�Ol~ǳ]�<�~��w\�^����1�tw`�A���}�b#���/�D��v�Յ�;YÍD����ǥ��םT�8WVn��H�ׂ��qIE�J2@0B�b(nd�ʀ��;��XO��vm�!���3_�Y��qn�\�Y������\���1��F\dM���Xx+ԛ�2AhƁ�!i�E ���������/�G��|v<���r�&�W�Е��}��j-8ﮫ��Z�B����A�먙qwg�ŪN�Hu7+�#��w@�O��oh.Cbu��� :t�(.̀Z+�ZLtWEW Eմ/��&?�-W\��uh׼>�)�׵Z��i��J�����Qq�N�]����̂�Q���Dy����u�e��T_Hq�ٕ��d�* �L�~�c=��R�TQ!���xv;/�	�F��\���h��<�Vt����,�i����KUm��?D��S��E�l���|�e*G[ �����(ҫ�Zt�H5�DAZ��QS(z�Zf�Nع		�n�Y���=����6Cvןo;��ۇ��jTa.(&Biȋ��`��������3w�y��8�N���P:�����a`�j�WS�EE��U�8����C��t4�3p�?���.|~�>l<D����ʗ1o8�e[��:�����):jΑ8�dVۃ�@���f�i��Qb��q�F�Xb��Vǒ0��hvP�g���c���%M#b{PvY_����4�]���j^PG�Aݰ����ȴ�7)�`{[l��M�2��f�F�!��
u�ON�<(j��r~�ۀ��acG*�U0�$��fu`}�db=��L2�������E��Ns�UU�w%�p�ؓ��v��y�� ��d]��6����y}`E���}�6H�m�w�o�b�o>h���z�8뗸/N,�*ܴf�=�	�6�ԫ���ݝ>�qK�U��|z��J[A�.t|5u�/�IZl�.��B8�f�~��m�{+l��C��$þ��ʃ��A���g5�c����;�b��r�)�@}��~��}rHH5b�P�۸o�Wt� �V���w��!�~\}B|���ǎ�(���vW���/���+�o&x�PD`Z��xY��P�oGUkXY�i\�T�mF$w��?'�����|s�4� �1��b�6�E�OK�h�c�D�{D�fy��754e4#N���v����:9�m���V�i����� � [\K�(���۞�|E.�ĕ]��s�����O[`��b���K����=��n�8�#1� k~�>����f5�s24|t�r�ƻ���Я	�}��?ϡ��J�L�\}*�ި�I�j�� ]:&�X���f�Jw�y�SH8^-�.�r���5ͧ��`���ةX�v�$y�딸{�P�6�aX��t,\�f��
$+���^�U�G'���Ћq���}�6^���B��h�֞��@�[����m,�StX���zrF�fe#3c�ST���&�ۇt/b�:�`��u��z1(S	_��HI�Ź���nn���+~��/�W����r ���h�R��*bsMG��R�#��Â*�ʮT��3�M�@J�^�I;C�v���"C��Vd�'�Zs_��4��Y(��}�ON��j��y���kL��Պ��>���D��P˕����5�]߃E5n<y�xҞJ2s�y���Dő�p�F��6\�U1�o��֛:��BZ�#�؍�aq�+5D'19�An���e�Up�xl~�`�A8��C�q$���L��[˭]��Z���~�����|�\�fEz�1��s�'�<x���@p�����7>+���X�X����n��R�1Y��k���?+���o'�t�b+0K5�i�1	/oryܕ"8V�(� p3Z��x�H�y>����(6b��H�� ��[X;}K�jؑ-��H�)*�l8�h���a���>`pb4D?�����\�Q.��2l,О9&�H��`j���(�[D���^���S���F�4,@�Is���U���c�9(J>���Wl�U�������Á����S� I�y���5�`�cD)������n��Z����t4E/>x�A����'��
�����`�)��RԳ�P~��Ə��st����l�lݪ`�n[�]�a�4���9�Z3��iN�J�>y!Dɽ����J�]̕��8`�����/]!�ћpai5�M=���S�)�D��]gB��|���It�{<���_���U�i�		�~E�b�[l�8z���T��Yj�����FL���zZY�컙����$���|/1���7����o�ɞ�s	*"V��\�ڪ��=��V�  �xK�lM���U�B]�Foܑ���R����z̶�ޯ��YǛC�XN�Z��d`�q)��u[�>+1Kt��NG=��m�m�H�LEmײ�$ �������}>���r%y3�:i��
<~	���-�GC��4m��������0m��Ҕ���i��v���Q��l� ���wq.�]h��eH������_��-H2s,(׾��B#؞�tRKM�~R�FSD�6�L*��Z��|3�?��2Ù��c�;��S`�hQ�z�ʅf��<b��Ԁ���Fi�:,W�K�ܣ�Д����$/iA�u��Eo����[4ͮq7ؘ��Y�3J�F�}��TeJ��C~�
3�H�����7.~�=ҽ!1��G~0ML��a��l|���Ň��_"�HR����^�����h�k�!�7 8 �P/s۝�@�Dָ�1sٶ�ޗs�z�I��l��e�ܢS�`���F5d�=/�����h���CY�[GOE`��j3�'�]����X����)��
�\)�߅"h�����nx O{�c��hY���͒��}��ݣ#}�p�C����f�q�:�ؓN�{���E�y�du�'��m�63��'2M�HV�w���k.��"	��5�aqp�t��ǋƺbE�P<b&9<?m����FoY]�1g��
��1�}�B��i����)��0Tc5!���]�d�`b��*ecG֎�0Y��nk4�ms����z¹���zx�`vۍ ��bE
%p��9�7R����0�0ZO�]b�F �kƹS8o�[���p�#��U3��g~��2����G�Ad"�K�^ޠ��1_�4��i��|��w-K����$��
�J��5W�}�	�y��ۥ<Vc<X�����	��T��:���۠��8c1�fS��������(i���<�'z�į���!"�n۷�"Z�;Dm~��V4>���[*��{(�r��j���h5�]��[�f���Em�^��:.�ҏ	?�B�q��2�􈄒A���*>����ظ�����Ar)*�9a�&�_��-��6�A� e���Nf��8���Wt������m�� Z�M^��5�)?l7��G�Cj�D�B��{������*k�.-	�Ui�����kklӼo9���ԣ��5��H0��Cu�>��~�`�>Rw�A�)֭�_)�fy��p{�@�&@�gmD� ����1Z�^+�m�`J��ڔ��i-r'/�eǯ@�7�)+dL�{@���<�<��ts"wT
x�5+Ӛ��%���� �H�0�U~ԉ].|�\�ϗ�v�<u+J�#���"��)�h��+�!��X�t#Ȅ��7�;J�=ZZ��}����^��k�U�,�#�D�>�m/����GdO��SR��C����(rw��N�H5�x�z<�X��$�!�+*�h�������J��6@�DF���T��J��;�)Y�����"��!��j�]���s�s��M�H^f	\M^ ���3r��Y���7�'��3�=}����ғ�F�%,ٮE>Lf�`V ����=��EL!?�@0�HR�R���o�h8F=Xw�����b�o_��5F�[ӝ&2�g����`X��N�!�Y�է4B#ϷE���%KJ���>������m���uh�g�mJ�ᶏ��e9���?�R2*��*?[f?�s��6-����F}y�!�'��s�|�=�e?O�m�R�0f"�liZ�r��LG�N/��5�[a4�ɤLҊ=c�~��m#��^�4���9���_���0��z�Y?5�c���q�򽙵�'l��r�6����T�$,�4O����v�CS��Շ6ÂK钛�����aٌ��'H�oq�ek���P�#]e�Qr��O,�˼U��xU�\v�x?��&�C�|�G��#}@�=�M#`�_(%�{�b�����a�46����s�h�~�k�[>��$�MDPd��e��iΰ���D���j�>r@��|M[��v��oOc$��	b�(v�3�6'IM�<�Is�u,�Om�l\t�VK����/��ޱ\ߎ򧀀��4��~|@E��1J��g���aG���=�O�g$�����֮Hɷ ��Ի��>k=��ޞ\r�FQ��`j�{9���S\Z³�+�S�9�N�;zi	�����ZNt�����G�s��CN���U���/�D�>��-(>���]
h�{��l#4!�>��kK���tf��G���K���=e$�f���^A�q��jx����(�!>��FpI���O��u��w�p�GY�& K�j��=�^Pl����Cfh�idD��bJ;�5Y"��1_��q�z˹Rψ��TsLa�J�(��>�ĉ��d�7�R��-���J^ͧ��ǃ�)?O�SOk4���1�����)����p�me��xW����w?J>�2LBy�Х)�.�Q\Wל��a*�c~I!��g
*7yK�D���"{z�,<V4<@ܬ�
��)h]��vݙ_x�ex4��j�N�PI�8��eF��F�'w���u=���E�6%bE��?�����S�=�<�*�'�-�����@ӣ�T���Ds��� ��[=#���ocf�p;�c��� �x��d�����&�������3.ܰ��,<��Vz-GO�7RI��ڥ���x�y�a��G�̞�^tk��o>�2����f��zo�ׂ��T֎��e:���ʝQJ����.|��WR㥲��l��#]�ob}�]%p��b˵-�&�3w��kKpqE��c�k�<� c�(m?�{"���wԥ ьr���2cy<,���:TŘ�T���P(@��pE�!�1�����K�iƣTa�=Rv�H!����C��&��~Zˠ!�=�.|���濞��4gJt�����d
��$�<���ފMlW*˝F�<(���5��0�t����c�1R!͓B:{�"���@q���kZ��B.A�Ъ3e�UJ�9��T�bW0������e3!�fi��҅�5����>N<�uG}�����[[��d�mS���k��1�|���oW[�.9v��<ՑV3����\9��$����<��6�϶�>�����
-IY�j��)�#�듇/�\�bm�?��p�*�NG���Yp}Z�	a�pfݱ[ nZ�{=��j�n
z[Ɉ�I�l����8U:�E,����Ϝ9mȐt��"�G��d-B#j�>���S�i�I��N{�< ��:�WxT]m-��pj��������Uǋ��g���NK̰c��Et��t݀�ó�#�_�عyv�(tyC��@�l�KE��5���/5�ŀt���W~&-�=$Ɩ�{t�3�a#�N2P��!�<�|ka��٥�8��0��	)N�I]����\ac4=B�N��E�ͮN���[J���Q�.��e����6�
_��ť.���_V�����5l��dus�q9�ILڑCN��M�0���>X����ϭ_�!8�c�Tob������ˍ�J,�HM����Ać^��M �����{:@|@i7�n��q��P�/5�����l%4�5�̄5�[�W�'�u\��@q��	R�K���Q-����掄�
Rx\�sԪ/���		���������[( 7\3���0z���K�#���aA��1�̗�z�����r~v�)���?O��f#�I&�+C�Ȳ���@$���qd�V���b"�\�|���^B?&���d�H{.��T���YD�2��)�\MW����P�3�j��~� ���??ΧV:���x" �fd���Q'5���8����$/�qb��u�ܭ��Z�1�r��TI���8l��Y�ŕ��(h�r�(x�����7n�ɮ�Os^�j�%� _�h�Qt�%A���u-���lˀ���K[>V���L���0%_70L����kE��z�,�˭��
�����Mއ�,]43��L���c ��'y`�L���'l�a@�C+��xF�C�%!�T��ľ�ZA?�v��b��`�b3"�m��#.�]Գ��g�����t'����U ����ʹ��;�q$G�����\ ��u�ڦ%t꤉r_7N�eIu_�-�Ω�!���<e����h�S��8�����2}�*N�&�5���1 ����S�m��:{�G|ׁ1��ǘ�=�����u�2̦�zͫ�j��q�%�KD��P�@S.�߰��CU��Mu�,��(r��V��Ԓ0u-l�^�f�N��m�3 aW���''��c�����"�����X��1�-��Ϻr���_�L%	ۉ/�K�H����h��o��:�W�h�C�I{�L�8�Br��Oy.}����� CDb�W�����f���\�Op7ҝE]�BLՅV�\�I.�/�ʜ��o�w��W~���l<�|���A���/ȍ��|�$����c@�;�w�W�gkC������L�٧��'�
�%�l��Z�,��F���֥��׈�:�sV+(
M�t�D7P$QOcoP��'��T@�SQ��w�#��h]��s����1)_xK-Lp�)�T�1��{j�v�7O�6[����ɶ�f5g(NN΀Pd�p|έ��cJ6�j�,��`�E����Cﲤ #��U���:ɫ��q�ċHt�gg�ZѰa_����}�u���Q�����쯃�+yw[m���І�����G �$}G'hز�
�fw치̂h�<k:oC)�@���Y;a&�ܴǉ���(?�s����zWK��=����lA�r*�q���&�FB����9[F�}�.=�4�p�%��y��
�>y�%��2^�TϺ�����ȱ��^��b���q���,�����[��2��{M��䗅q>|�S�&��D��l���v ��ͅ�-�F�|����2|F��܎�?��+Ɂ�!��y�<�`�)ƹqy~i�Sͱ`}�B�M��?�����,�з�]q�����( S��џ�|lJ�����<J��Ὡ~���e�Њ(6P�L�(��VVF���o�וzq��N��v��a�Μ�ţ��i~���d�h��6�/�(�*f|�k5�!6_�.F��r���4/�R-��\pa{��� ���9��D�ž#ͪ�����C`=���g��Bh�w�@��<����f8�}�\�*�Gl+��	fJ���4R��R^u��s�_�7B�Ml�d�O�%�+tJ#�Ѧwv��=\���� (J�{S��89,�Gl���u�L_��_���y;Q$M)ie�y���?��CZ�k��9�C��hm���h^�I��x}���q�>a�0?WG�8�4�l�M�.�k�etauS"H�P6{�\�~�}�p���lz�5�����?�S�������f�C�7�d]&G�K����1���v��15Y��N�2{��h5HFBT�T`TzT;k�M%Ǘ�`�%k�6"j�z�ݭRZ�b�̰,3�����>�-4Pmx�D�`�m���ݾS�-��t|M��8��b���O�V��QYt�@�te9��E�[�9굤<⪂��I6��7��<�������Pa���x��؀v:�]T�-pq�]$���3`l���a� fۿJb��ڌ%h3����zM'9ī�+�����gi����n��4�_��� }��J���o�21�q�Q�^~�����?́����M����H��8��="�x$м����~���ě�bBh�!'8X���;<�ķ}N�E�*	�]��Q��~h#;RW2�Z���8?�0�YK�fGh��kH^���(h;%<���{��c?%�LZd��
�?�m5�[3�5=��_���Y�:�ƛ7ى$�@A0vM�%�'	K�wd+�=�e(Btt='���7L�s�(�n:����Gi��|�@W�rj� <X<�Y)4��R�ų�gX�7�j����cxٖ�X)M=I1���}Ab��G�LkZ��� |ۋ��T���C45p�hQV������c��@���lA��\�(��2��o�ɰ��H����E���lʠۨ��Rv�!҆r9;�{�E./�(�^7���G�*���i����J�R<�����r��I���W�+_�b��>o���+3��k��.W �*������pP
�u<�����vQ��~E���E��:j~m�\�sZ�-Eг�$��Z,U��U��b;ͭ���d eBR[]j�� -���@����_��4͠OS��l�؟��Y�I�SYU�Ҡ�t�ŏ7d=���+�/�z����Z���n�g.ۑ���|1�oؕ��Z6+�_��V�������L@��� �] ��_����9�>����憔�hS������k,�:��E��_gj3�����,H4��
��v$7�L��X�OL�0/Y,�<����2P6ϯ��K��|���fZ�����?�qN���قc��VHG�r���^z���Y/f*��3dQW�_��(���
�r|��įh����t���5b�#�һ�`ͣ-j/�0��:�R=���C�����X5E2#(�{���8��ȁ	�>��y��C��G��xS���)����(�5�j.��h-w�9�/�� :3;V�2{�P�oG�m��C$J�
&]]�Z
b����>�~}��	P����Dh&����N��A��-Z�t��֛����v(f�&�x*�&�����a��'�>ZE�K��}茂�����\��ݡ��o���|���6��oqa,�C �x3�/j�>�55�M(�-�agL���p7�h|�&�� ʁ�|=�¡mLi%e�
�˸Sԧd����<:WB�ʵW`�D8�.
q}���0)�����-¨���B�;���2��w8�e;��p�tov�� �9�XxS����쓨:~aC�)N@�� ��}���� ����;��b����.���Ue��;'�����/��wN�f1��>�Z�-�|"�V��Xݩ. �[�Z���z4���b0e[z�bUm�#�IN��+���{8���.[F�����picj��@����̘���Č� 	���l��3��1<x ��#�ґ
`������YrFl��,���/++��u�#���7�11i$�z�)��	/Jy�W_0WK� ����~������H�*Ňp���,�lu��e�fJ��\ ӫ��}$����"%QxH���6�~����3L�mn[oK�ttO��B%�"����ث��=+fP�Y�����QW�Eb(ZgI��~Ǯ�t�{)�jf��^����4�tz�jݡB��t&c�$�\�*{�!
+�/�,��_`��������Y�1�:�ͷ�1D� я	�4w*�`d�e��m�����,=I����~!�Z_��g(<�C}&-/~�B��� �i�*����	��r���`���Išϫ���������$%�����h������>��Wd�f+��F=����8�a��̟��ׄ���z�Ѡ)[&ȨV�͊TE���21��%!R��Jy@����kl�E�s���H�[(ĥu���B ��D������V��z���I���y���#����yt��E��d��J�}x�B�?�
���
����H0v�;96����k��z��z���Ц�7f�sG�Z���1H3J�f����'r�DF�������X|A�y�x-��0�ˊ������v��
�'�*��K��W-����I�K��x�m�}���L�Eu�Ҧ��N_���x�q����9?߂�2b|Պ`J�l�^G�]�ʚ���{We�� ���Co�0���)|����zutS��Z�x�|�$�9��<)�%�L��4�?X�g��5J���&!�K��꿱��T��C��b�U���O��f�G���T�X5�����*���;x�dE���
C�(�o��Q��'e����إa�vC?f��h��y��Ӓc����nG5$�e��e�����\��67Q���/V��|g]u1�k�s�K@�j��>�Ʈ�����]�9���dhF׺�N����������1�p����k�TD(h�V����2|������؏���r�(�2�!+�'�����ɐ���#D$��hr�^�7�J�).�������u�����7:��C�4���{����Vt�(S�,
��6���� ����}O|r�0�Z���X��'V�������^�|�1�pH+�J��g~��CB1t6���
ئL*g<�_��V��%�IiJ�����������w6�
"`�����/8�P?a�j�{q!]k�k_<6���#�*p�7���x*�#��5}����?'$�i�}
!�%19ḽ�Ue�\L Y�SP��ܞ�d3݊������~�	F$ǧ��%����7��p���b�a�؃ý�r9�]����|��/����޲��ml��o�`�� o�;�Jffn�����A}�k�������
Oo�fk��	��d���t��*�)�=��/"
d��uXey�W��ݣ����6/5��Tꊨ��m�#~�8�%|g�z�D�H2�jPr)d�da�Y��q!������5��S�r� �/�2�+�L]����wB�����n�:�������\���/-&@}w�ɱF���ȑ2P�e�Ǿ��9���Ʌ	`k���� XFOl-��f�z�w
L ��E��Ygg�W�sS��IW9�G��>���3�R������������^^�Ǭ:� �F6�ܶ��ORR&�(�A��c��K�4�\,���ag�P���3Ѕ�T��Ь�6m�%Y���� ���Q�n�*�-���+��ɵ"�Gϙ�4��!	7�T�x�#Q�r92"���9�2�A�J:�5�9��"=`��.��"�\vM�*K5����"�Qs��#<�U����ƌ.3m�rJ1d�v������Y��T������x"���i\���T�E=���ߤ-�4�����8�>s�ĵ:��_�IB����d����'��πat�K����BԎ�5;Rz�������U�lqu�+�Q���1_Җ�2�.w����5�����K;����YqjH��|0����o���-�*h�m�n�%X:;�a鵰���Ԋʹ���I4��-��6T��-'�#��yA\�~IA�U��G�C� Ϟ�,�z���.���.�tr�S𣈅V[��X9|��}��%UED����͜�Q�X���:NZ1��o���B� l�9��b�ծb��Z���9�h�x��������G��U2�����S�!G�G�z{�哏��@��� =6��m�+l��$�`���6�c-���[�g�M瘺��wz��@1�`�g3����j�l]+�C���a*�X��D���Ul�s���ഋ[t����~�sk�Q�wp�7,ǣ:�R��?p]�,c��E���/�Fw�j�E�?�S
C�!GT���te65v۔�'�\����$�l@BPLI��t��=,�.��3�YF��9����ak�c���ޓ�%�Y�lpqq�B� �I��[�qVî�ۡ��C��d�^���i��1��T�ǧ�!�7�dۄC(�b@�*��g��$;#_��1m����܆��ӷ�a��;s\����b���U�����ݪ�,�ʹ+�G_D��;�7�}�c���p�Y;��*tӣ�X����:��\t�%��=���X�#Xp}�$v+i;Y���K=��MIW�M�P��� @�T���ҋ��G����2ۃF6k?H�ꈋ��OJ�_��%�m��K�xc�\RD&A%k4�(*�X���<M!
��H\t)�lF�{}H���M���Ew�~�T%��d�@�����6��s�J<p�x���`3c����,4u�Q��,b�l�|`�^��ц5�	��n�uX��e[��s�wC޽��c,w!&��J�^J�j$�A�H�K^0o'8��(�1�H�l���97�����Q6\�V�2D��d��0	AP��::� V�Z'��yP��(JUb�׺�[�r��L
��6��(~ZgC2� h��H*7�n�_I�5�B|	����P�N͋�}�M����E��YHt��z|���g�"0<�ൺ}!(��9��Tv=��(��]˪����&{+�.���w��O?@��x[��%�*[�020o�����n�#0�Ҧ�F��+�Zʞ��|"�:�L��2Ѫ��_p���ʻ��,�`] ۑ6�$0����P�����S���ƃ՚��4�Q4F*_Ί�3��!���6���b˭&!�bC���.�p��v�z�f0?n�B�k)��ԗ��R�.��7z+ ���'[���9�^ғV�*��} �hQ�����Iz��kJ?Or��a�|�^�	r���ĩ�Y-�F�a�CΘI�K�L��az�΂IJZx�G�&b��E�1�ϳ\Q.�->�2Z��0l/w�s�8�/�L��$e�K����٠�a�5la⪹��B��K��3�xZ�TU���m_7���{յ�k��N�N��/��m�M��5�)���Ds��;��g��3+�{>���Wi�+��(�����U/��#=��IZ�8e_��jy@/�n�w�ǲP�Y��V��k�,Z����"���z�(`[����7�\ᆳő�"�)�K_vaDB�V$ʸ��G3�$h �k�	��M,7K;|D�0��3H����vS)�߃B¿����"��C ���pvS?�@.�E�@�#�J.� ���V>B��x}�&$�-��V1�1V01�[��[�bAl��if&M��e3Z,y�a��*�]���[��B���F��b�������w��
;[��i'B�`s6~��ٖ"y'�CQ���e�7�d���%b�',7	��	�`;��d�:�z�zD��$�۵˻eI*%�8���9����B�3}�K%����T�suh�<o��a���6P�����^"����r����i?����g���iK"�h���s�DVP�
={���}��ӧ�(])w�
�����]��A'�C/�����x��Ex7����%;ش�٣��&���{�+bdQ��q�>@̥A{7n�)��eȜ�?��٘:��[�?F�gj�F�o�d���Zӆ��>�Q�v��@![�2��'m;�.��Յ��%�PT��ioJ��,:~f��hhKy�[Ga�2� U�i%��B��v@���"8>�%ѫ夏��\h,�	<�����@��qWK=��PNa�IJ�F���v�g��b'�A����]��`b�x�ޢ��}���i"Ë&�;���Âb��8���֗GڴF�m�}��E?�I���l�M3���>��%��4�+�g��Q�=:�ݙ5�Hv\�M�a||)�������\C�R�k��$�]C�>��(�ʞ��3������=5��R��*��&;��������G��įo�A�H�,���@�(~�R�l*�0�vcS˚���A�G��~[��v�^���� ��ʛ�$�yyԃw�}��{4���0l�Y�g�۾Ny���y�r��g����ӊ������H�Ց��<�I@~���Q�]���X_�)��@F�*v߹K�����ȫ8�HƘ]Cr������-��r;!�A\����0JD �A�~@T���-��z\[�ѯ��e|ʭ�f�b�r������8L܈3���X�z���}�bQWў�q1v,���f)�X#.s���PUW4A7	�|�{�Đ�&V��2�.����J�Sx�a���L[6��3����ø�5$��e�lY��C֌:���-7�ZǱ>�������N1ҭ&����2����i���_y�T����$�k��}�I=�VJE��o�*2�*]�u`��D�:�E�,Hi�R�/z�5�!s�Uşx@�?�q��sB�P����%8���G�+o��a������p��O����]��� �B
;�5WPz�L��W&��#A��U�8]wѓ�1[��ح����.��-VK�&��m����Z�ԡ+U�y8��v�N��w��
2�P�P�(yx�l/�L���I��2B��ǚQT�q �N�U"x8ZY��)����M0#�D�5��'χ�ts��XUTF�3�5�v[Fy�h���\䰪g�de�Z�$ϯ%�|�3:��!�N"W�t����urV�(�4L�G`d�\�� �����c:[��Q���l_�!�:x���2�;�Յ�e
�f�v���)�	��<:��[�a��&�Ȱ8�O��7`Ns�^� /Q=���fw:Y�:�K�f�N:��<�KD0�"F �����LW��`՛���;��-o-�hc���G�W��iУ͆H8$�&�-@�}�*��4?e�^��� tև518�4(�L�-��e9�c�jrA�&x���Ǳ߰�>���P�n1$Z�46��1xq��#%�uK�%�������.*P�^7��N�c,w�e��SHqq�ї(Zx�J�,�w^�Ν�CƇ�%�Zn51� ̙��<� cnkrXuS�*�1��I�X�1lZaކ�U&��wUk��ƌ)zZ R*	���ۿ2
�2H;�ɐ�c,ϲ4�l:2R�pg<�@�t�b��Y��jH����J���i��Ng3�gP9����q��d�]�k�_���H�ӆ�e��̍H
�e�$�r�Vۧ}.)������7.��f��w��uS�����1��G���F�.�ޏ��-W�E<@|���x���)¦.ˢ��;��?����r��;-�� ��Z鼴Ì8dq�6�]�����1 :^��!n0��o?������7�4ķ��:K�/��doϚ���Θ���aPWt�Om��17B
<V2o
�]J�B�iYf��#&?�B$r	�O��*m�=��u�+�����I��aR!Oj �!�Y�B
��{8C��lj)�ju�e�6,�/�����}���r|z��Y�E�U�C�C������Is�uU�y�����UO,o���k���R�>CJ��pچ��1X;���
ɒ��!_�HN�t��V`H�&#O$�_|G��%�����\�v;�,j:��Õ=�t�"�qY��э�!��C�,!{�키��JK����1���?�2/:8�n����5�f5�eU�hw�)ie4H̱�ϟ�� W��P�?ٜz�d��O��R7ZX�ֺ�������>�$��7�"&�[��iB�3y�e�*x2��h 2~J,%�`�\�Ji�G�xP]!��
����+�m��AI/c\�/�@�冎����K��$��{%�.�q��)�=Ꭽy�s���&?���-���^4�*����D�8@`Zc���lP�B�f�k�(�[���������݂"~��p���S�.
������0=^�Jx0s|t-m�i�\����+Of�S%?g���@$*����MCƊ&@��Ԧ�����ZWXA9x��(-�
Ā�]5֗ހ ՀD�(��$zfK�pٰ���2�t�\�Ȩ8P-+ـ����9"VQ-מ2�>
oI��,�R�\���#RG�.�X˂��!�>��O����z?:�7ꚙ:���2�q��4�e>��l���FO����d����NYhK�״i ��$�ҒI��p���W��t�<_�[R-�Yv\�!$e��7��k�8X�`�E7�J:P�Ŋ�hz+YWpֿ;K�.�`R���=B�>�PJ��H���:�T$X����>&P��0�~'<����`oh<�.���r����������3t3�k��Zw��#��)��'{D��)˴���+=�҇H��
XdZz��X��ʟ�?g[`�}�YV%V�ˬ5���[f�Ű�&�uV�]���<31m	�`�m+�#���G��=!���47O����pxټ���v�}a&�����}}o���F�]PT�M�ӣ�~d�,L��/�1�# \�<����1ig��c{��W�e�']���ͪW�axs߼su8?x���h�jvv��͵�㩋��xTV�����@=�I��d��j�����4	4�06�P�)ZZ� �PW�:����w0؜�`j3;ڣU�*3.V��E��V���~i���F4|#�_�t�{1��ֆl
C�O��A���Yu�߁�쫴t�1������W)vu4��
v�Y+b�l��u�*�(�|^��|b=r��u��%%��8��3���("�U�1�g�	l ��{R �j+��@��A�I�Β@�s�l�wN�}�Z��yiT�Q�P��5�XJ��~��_l��H�
��>*n�� оQ�':�z5����p�)=l�ڎ(�m��w��.�!�}�`G����i]��A�E1��*�n�pa��)�/b�8�/�ᠦ��%*L�$s�ApNؔ���Z�ej��u����h����h\��	��A3��fף�d�}�8��vj\�yl��9\��sl��w��Aā���.��d��y�m���[�j�7�����9�{��`�t��/<=��ޝ$�Ξ�8��!��C��L8�� �zhま0�@�g�^���q|�2i��|e����̭�C��m��)��AԖ�W�|���X~2g˳y�N�Cɠ�Wa�`U��w��^���AOԍ{:@����ڸ������&��;Ҳ�g�SIbKjD�\�I�$��u�%���*A�u���\��}��7��T��ឩ���M+ѽ����]���7�u�5�.��y�Z�ܞ��~Ot+���A��%�}��䋻���ѧ��D��p�ƬD-aC�EX�]�'_]c �|G�~@��J��m/�~z'=�H��˾�ht� 9����jVߍ�	ܔH^H�+��y���:+��=J��-Zu�"4?��d����^�����^>o��8�g'�^�i� 6K�?4e�)7�	ca{U&cc�G�9{5��QH� ��yY���d3}�o�:3������V�,̛:(�a�>��u9��BLx�J��3�A��2��K���PA�3��!F���3��	i����0����tc$�QV��K#�h�s��!��?A�x!o�G�u�/�I6�"V��rnξ�O$#g��C]uq3���މ��iK(�t/&�q�Lם2�r�Dо���d��n�kт@�^�١��jG)�#�8��=-1�A�e�գ8F�{�/ٷsBu�{�d�Ѯ��H�Ca�أ�-�Q6s����J��|HN��1F@�B�X�:~9b�jf�'�G�.K������d{�����)ᘖ߶�J?V)؛c��j�|���� �����w�����$6P'�婙g��L�0?�}��IK�݈�
����ޣ��z�Ri�F�(ѱN�x�����V��1~�M�Qh��@&�A�(x3n�֞}���ֽBEN|(�X���狨�����h���ŕ���$�_���z���<��\��ݴV�"1D��ɥ�P����K��@�`�Φ�(�5���J$i��������-+s��Hu�t�`I��^��gj8�+��ϔ����4��u�泅L�>1��o�ݰ�j��*�'�B��+�����
���s~�Y�5�`�zc��;�l�ä�(�
�_�}�X
���K/��%�O?����r�ƘR��]��5��vt�-u���Lw_\I�����~O7���I�W���B��:jF�?�����/�n��TYб�Q��e�q|(�x��������X8���A�P%�F+v�ם�L���-T�e�p��<�jG�k���,�5I�k�O� {Uh��1n�'��1&��eo�݂�V�J�}�o4w�iv�-��v$t�k[�)bE>�TW��1t��u1+�jE���Bo�����_��&���% �vBn�僴�N���i��R��ʪ�2 S��1���$F����ʴ���ԇ��D���0����f����&�p�'�C �z���积���c`��G�"��}���3�r\�Ww�->�.zD��bp�u:q�7(HsgL���i����H�N��<�1.���8���"�\����
�4�l�Y���l��"��Bah��H>4EM�f\"�{n���p����{���ݞh�.��K�X8��������H��ILTp���[�qc��ffX��Y��s�y������qe��'�d����ӛ�*\qI�����_[O(b}c5ǒXv"��s��d��)��{���
�c#T��-�a�Z�ʘ̠�K�=��ɵ���~�r"N,*6�׮#ד�X�4��l2�q�@j�����m���i닇���Ibvq���rը�w�{��Qjb��87���R��y|���f��ը��ɤ*�2/���͑�J܈��o� �PV�K��MKa��ѹ \����_�Q"EҌ,ߋ�P�%+{�Kb���h��L��
��Yp�����)��:?�V9��;��t�#q���n��(o�1�z���8�^��b�F���r_��]�ݳ��}6���1��CO��dsf΢�їC��<��ĥ���X*�����[],����[: �9����A���Y'�)AR8�f|S���s�˸��wK��q��@JL�IZ����6\���u��b���I�R!�֬��; D��@t]O���(*��ICf���1o����M��t���߫�2�&���D�T[&	)���*��z���� ����M����M�����m��C�W�jם�����q�;7��
�_Y��~+C�i|>�m�)�('$������b�u���{q@"c Jq��/���f2�����,ǩ���Y����l�E��Ʃ��q>����G��w+TD�Uh�e�8ub����ٜ��7�	E��|�["ܕ�62����L�t��_�3y6�:��� 0lòZ��ۂAA���%s����ގ�{�l�K��r�`rk;�h�qɵŨ粌Th�����&�ˀ섐�Am�|�<����>xA��nƼ��Zx�쑜�g��>��������x��|ٿ�*c��vޤ����B��?�>)��KL����dIz�5Hʱ���~,�D�q����xu�<��y��$�f+�">�xun-e�g��9]!}�m:<��	v��($Ǫh(��Ȁ<g�,6��e:�NY�>/p$8W��mW�l ���+�>b�N�Hs��G���l����k�j^`<%�&����t~�+�Df�1��,ol�\�j.�O�y.�v�CNu���r����U'����B^��*g�.0g}��m��cH9�9p��ӈ�W�׻lQa�з��"���F$Oi�V����?AR������:a��19$��E����?6�#0n�?�#_U���H����D�V�#�M�@R�}�Io7��P�n�q�yW$��_BE�I��`�a2�����N�z���4�Qm�Ǿ��~���/"��թ�ې��#ԂQ@^od���R�V�dW[����P�z.{�,�5z-;����^��<�M@;�6���^��i�`�X@�&JE'O�;a�^5Cf�6�#�&��M�mK�28lCx~���Trn�o�B�D+��aF�b���l�,�*y#�%z�Ԙ#����!��M�nJ(����<�x��-�L���y $Z������:�努����T�-�)Y!���Q�"���$5��X�l����k�h˙}PL�+����	z�'"�|l��� �n(I��Sk��4B�-��9\S�c�������Y��Ǭe�E�![��+O%V1���@?���̺�rQO�х��^�/*�h����m��h�@_*�����D�'j�˰#Z��切&Y]��P��=h��"	�n;�Z�x�x��g�%J�����<{@�kKd�-ea��~����A���.��s��8-�fJf��p���Ӫ����}	�4Uog$�P;S���ߣ˸��o�P�BYI_���Q�9�=�(�*���Mm�8%�7�~�Y���ه��Q��C[��|e� i^�o��1���G�祥�	�霈�����$�H�^F��O�����=�@fGE\�C":��'��0ӡ��T�2���z�$�갌����ˊ`�S�H�C,�����?ԥ�%��Nb�8���מ�f��@�6i�?�;���cD����O�.�����
�zy� ���3�D!o��\Mh�ј�m]����V�pb�b���1۩vDv��-�n�SH��%X<c���� ]�;T�o[�&�䙝��6���ln	��w�iǤ '6�Å��/�uu������j�*S��#��jҁ���$	j�4݄מk�����m�y[�|�2(�����W�&P�̷�I��Q6�v+_���@Cd;��3�����jB�ۭohx��/�ݔB��ld��"^��H��g0R���AY�� �����5�3p0�髏	}��R���]���}����C#�:j���mA ���̛��=�Y�d�5`fy�v��;|��\Xa��u��%[h�	���;�?���4�5��l�]w�+�,X*���ɧ��?Dے
�����������H�Ҏ�0�kP���e|�.��f�Q&��?4@�A�[a��|����_�W� �l��z�u{�De�F��P\<@}��� C|��`����E���1J��|]��Pg��Rp�2���?�2@�ܓyE�M��C$y�
�E�!l�(�<�����v���H�TB�ti���^��>nߏ�y���*GZc�M㷓58h���� ��F���a��o#c^����!��K���*��wy���h5(�^F4�fN=�Oq��9�CC�ıű��@D���`��>���g��v@���.n�0zrΩQ��� 7�7�\�d�@�Y/� 8�uc��.�4��-\n�:�wz���Y��P�E��$h�iȐ���:��%��@�V��+n~��I�o��e&<��o�=��b�k�&�I��+y�=r��SNv�9蜢��j}2�"K�I94*��/����a��>�/�?�	n�o�Q
�%J��N��.��3-0vE�[�l.dU�g<臧I���lhA�'�q;��B�'a�B���O3t��?<>)Aڞ'�J���VÁ\���%z�%��kLZl� \1A��Q�b�ލ�����%/�L
��nr��@�:�����0m	`�/d�XP���\�(�jnT�/ؔ@�����>��4A?�An}�+y������)�A�G�qt����O���Ji��>����0W���
�:0������.i$]�KŘ���X���2��'FG?���z�Ifq�'�J�U�M~B�4�ljWj���
#YDp9d�F�F0&p^���H��p

c�$Y0��w����% �0O?[!A����Y�k:ۈ�&m���f!>�Ɵ?9�{򣹹4fs�j�T�.�p��
�Ri=ڛ�$�z��Y?��F�7I��Y��8UǑ�
�2;,|�9Li9�Z�F��1�ɋ��tO0j�T���_3�w�vc���&��M=��;�Y.��j�G6�wc�,|�˩�ņt�_��[^��
�a�f�{�{0.�_��Gys^�TH��Ō�r��"Xy�Y+�X���]������������Ps� ����Z���cJ�!��+�e��>�L��� �,P�[Ҫ�*�bA2w�'�~���m�����<إW�oS9��2���a��WS�,|]ϰ�v�v�E�EM����~�)��V��(�Z�D,Zs�0F�w/q3���F{#0-&��Ll�|�9#mF��5�K�Ce��嚘�J܋�ĖB�·�l�A�x ��:���P�D�;���|w���[-#��xD�̦�%2'6�E��'�SB�2[q�	i��}j�ܪ'Ԇ҉bc*��7^���(��%�,SD�4L��P�?��6�c�h"���f�j��xi��L�[���_Y�L���$+;7��xG�FeF���u	ڷ� V��M��	pf��$�8�����&W!��$�Y���2�eZ;����=�BUo��đ>=�ۈpn�rDTR��.#ҩ�B;�
>�ɗ/6�s	lpe�D����/��|�&��tu{�>=
涞�n/�ݧk��uQ$�=27͚?�~?�^5���)�nh��2���R��n��|�>��u�Z<��VQ��zz)n!_�d~����B�i�����z���4#�c��{O�|�����u$OφY�7�~{a 'y��^�c(_wM�����j�Dt_��.�xb�M~���y�y4o�"�����q�&�9KP�'���aV�o���$��@� h��r�I�I�v�<=�V ��ke.^�D�䶢F�����:�[T��υ���Km+��W�	ǒ@�`��U��R���@@����R���Gn��߬�ɵ������z�ʭ<[&�"r���TB����tF�}
a�z�����R���N�� �'�Zi(1�x0��~�4cdTKKQ��I7�b��[�.L���SR��evꔌ<mSJ9)<a���&�޴�&֑vl��/���U�L#�l:�#,%�fi���@It�x��x�cD�uAH�ho:z
����	/ONd�C��5�Ky���3p��+���fx~�&<�#�R}�� B����u��+P�J�;/���L��������2���:�bSi���s�ge �N�?��>Ȣ�ul�Gf���:2~��LL��n����8��U�(�1�������07X�b�@G�^���	���x�h��lg})��5���&�b���$��Ȋr8r}is�T��������3�bO�Wc:������מȯ���z�<�tV��Y�i����LY:��c��YP��ͬ�h&Zٰ�%������'k,oY����µp��:����a��ј�����cMRl��[��!�-�Ѣ�Z�d����FxFG*`aK_�F`V�����;_�Oo=��[xl�(�]����𤂵���=7�Ȓ{S�d]$�BK8��Z��  �o��q�gpFN;�~FWvn$�;!hhLqyQ�*G6KF�&�\�jH�-5�xP����UQ2'L���DY���d���]�vە��/��;��}]��k�|���Ͼ����]}5򸤮��tQyF��1 ]��7ـT�c����l�V�W�]�83�r8�QpM�9VZ���Fa�O\u�Qu��|p7� ϧ�H5�����G����:\��(����^�ž/(��Otf��>�O��"����A1�<Xy-��ڠ�y���ث���fv{у}&�n�3�x�]iֱ�g�"_�����TAJ�A��<p��A�)
U9[nLI��0�
��CF@�b"u��U��t`*Z������3 ����c����+�nD,S�[uq�b�����MD� ���
g�@vr�PU�0�Q��7���M�v�Y��o"m�Ռ[�"���#����fQw�X�wnOR� NA��5P!)��"�^7s<�B8�=M����_;ި�e(C�4 F� t�wN|:\��%@z5�`��&��?v5-,s���\x��$Cn�9.*6��T$O#Wǽ'�@F_���3$���~�VV%)��]�8�?�p@��r� ��=y|-��/��`���&ܱ�J6c���Lz��x��*o'B�1R�1{����d\�8�	I�vC�Æ���������[��x_� +������G��(�
 ۫ԛZм�����Ӹ�P��Zf�M������j���:"Sm�,X�����`m��ҧ�F;yV&�nNr�k�����XȲP��k�GCO�ӱ/#aS-Ӻ�3�wY>�7]�rÌ���_I�  Y�S�OΞ 10�*j$���U���f��L*��&Q��.�§��Ko2����S�;�0�-L��n����ĄY�>��BO;���f�T�zH�����F�9����0�-ƺނS0��� �km�ӡ)DS����;��H�Y]�!J�#H`}YZl��ɬ5�X'�A����J�kW�͵8[8�SS���V����Q��3�mɴ�XL�AN��9��sՀv��ؠ�#V���|���a h���NM�Q� ��:�fu[>���h�06��7�v�����dG��-P�����U�;���/�L6��*V��1/��t��|N�b���a�e#�i�[
T�W�љF����q3�0)�`<M����y�XQS���'5���E0���,��|���h�����rn�K�,W��0���mE.G�"l"�^@`�����M����X��$�]t��M�V�Zo�-m�|�,̓Ws�U��	l�(�KydU{&�Ady�*e�O{��vL��_�?L�6v�
�ùo���[��</�߾�uN�+���̀s7��� ��d�a�_C�~U;�]�ZDG5�ː
���˼��JZ>۸�H˖ڋ�;�4��h��S�S�	��	��$��o���Iثi�_��U.�m�V�wJ2O�E���&����0*��s�@���K][p��0�� ��%KM_?�L� �ĖΦ*<�w#a9��g�2q���̈́�K�#w��T��������>Y6�j�0���G���b;ʙ*���Z�ls�)�g��z��A�^i#7l-&�5�����ZZ�a0��E :r��>�8�Z�$�fo��3�f#[���f���ّ"�{��lN ��(ku��?��6�N�"Osi�*��@vO~���{w�&��Ğ�h��#�Y��dץ�5?�>�Z��&B������~9|K��G*	B���	��^lj�_ٶ �b�]�D��HJ�����>({�|Juj.�����紶��{����#�'נGw�3:�e)��u�`��`��#����V<��L�M�������'�;�?^ ��E(���;G�3�� #$��<����9_�1�<�zۊ��yD�������1qh�hN�_��2�����ਬ��a�0 �?�m'%��qZ=$N��}�}�#l�<pz"f�<���h�6�3�$����I�iְ�@ ��T�ۺh�����WG�Z	��
 $�ݟ�a�Am���n��_����2I�^��P�cu�k�Y��Z�������Z]�5�^_-k-���<�;�������*M���C:�{��&ރQ�����C}�' |��� 3�lK����LQ�q �s��|�j�_�LQ4���z���n�m��՚Ce�{�gt��,��c���/o���~'p�3ٖ͠���'5|�;�U��e��B��l4}��X�Ɲ�c�t�B!787�$'nȿ��h�S���<	Et\5�fy��A��&e�-Dɤ�RƮ��		`yB(�������$��)>N��n�~&JRS�����--V�D#�Û֑_Ə)i�zs�60?��2���jΝ��^�[�(��s�>z�a���v�����$@k�!�4�2R�|��H����&�?�3�Y�����/sD�*��`}��*��K����4��&��~�(z��a�)۵�
��_,s:�`J�:�c�
���|�n�j�Z�+ 9��ӡ��!q���f ]����o<褉����X
�Y8���9��4�I�خ).���*g�a�t\���c�M���j
�ĕ?��,P�yI�,m�mi\�:�<oS^�J��w�8��bq�)���z�*��e��u��m�c��C�T��S�A��	�����G� k�Q*�B��L;2�Ֆ�4.��=�xp.�*3	�����Z�?t8�g��=�ك�,�9��.���ݓA"��z�qm<�0�m�ד�K65cT�!�%{)�7�w���P5g&��:0g��b�{����*|�=���D�!�{�(��R�o?o�X���͗M�v5�lC]����=	�a
�A�����P����9R��jAFN�PS@N�!���j�	ƚ	�4>%l����<V���ck��P��h�f�۠��mW���_!�D�!�ֵ�p�~��F-����f�` {�g#���PՈE6�2�aLX
���}m���,�B� �z뷫<����ї����ĉ��_����S��
8�C��7&��p��'B�,x@����)5�l^ˁjZ�.7����r/�Ě�^`������?^M���W�$RnS�ޝpe�o�bDK<��?aL-��E������nZ������=k�%k����w0��X�Su�\�,N�Y�B�!sح5�#a��M�[����6�%�fv�1�H6���A��%p;>n��v�x�Eo�׬��'%_5ȱr�b_蔜MS_$�����"�(z���Z�	P�
�.�o���p��k|Gil�*U����%��>Ҍ)U�R�9J_��[��]�����E�FT< Db�R�$[�&1a�o�Q�}|�"m~�����<����T��� ��;@�a��@�O2�u�KL��gs�^�c�J-�ETFJs�Z������88�,P�uM�-���E�7h�r�b���G\�؇Щ kY����V+=7�ǀu/�.M�2`d+�B��R�E���qȾ�	�������.5w���+[���^u�(@~��������A��0|}�G�ˢ���^+�kj٠��9���i��M`͑�Rz	�!A�F�d�f�E���0�a��c��k��}���_���:!�6	<7`�8� v�(�6m-`ֶw�l����H[���e ���6�>@>n�J�{yQύ�� � U�a���V�V�q$3�8��ifd���KL��zsC�^�V���Vcp��H�>�]�2b�%`�+c���)�ׂ���������Vy��A5G�Q)�տ����DU��;PP!NV.���+QWW[�QV����}ɘff�Jq]�,��/:di�L\�������W�ɮٷ����F�&i�����K���)7nkz5ҭE�/Cd{����=F�Dh"ҜWs�'��exn~�� �y�*X*��(S����X�6�>��J�@��z��u��z�?�>"�U(Ӹ���1Ɍ�1�OB�p����#`�橉�����Y,�j��9�c���w�da�j;����6��_�[��[
4'�s���/ �渘;���h#�>�oJ� �fU�&TI�/ހ���%IG���H0�B�q����ˌ�h4�����k;/_��1�f�BzO�0�7W'H��Ĵ�y>~)�R���Y�]�ͽ�`���.��Q�����+�c�����I0��MZ�L�������M�Ӆ3a��\7���:Q�}�T��k��b+Q�����Y���7o��K8w���I߳T\�\�X3G��N��S��rnǥR�0��fB��ev�eҜ����j*5���$�Wt
�}����`�j�8�1/�\�Z�!�s�9�b�5��E�^�'� ��\بo9�+Tص<ٽ�����i9u���!vM(ྣ��=��_5 <�O\n��4�*��dn���XJ��|�ݮ~֬��^=��(2o��dG��\V�NBV����>Ɵ�f������(����L���ϴ�Žlf�5r��ӂG爪p�*�7}�K���k�	qN���K�alò�&�;FL�����T�6�Ͷ �T���/�n�)�L�(C�-��#R�����	:$eR���	���;���DŒ��Fo�H�*��b���bN�%ʽ1[8)�ӡdZHY��U�z�J���B������vk��MivW�`D�3��'ϙ:-�� �[Wٕ呖^Ph���W���pӭ�$���]L��T�'OC������!Q9<�d��f��������K���%3*3�Ղ�0�z�|����ջ� ���]���'��g'�!./���O��|!9iSl���&�v��֛���.UM��#�̒/jC׾�7a	n➽_��-��Fsj��5�4n���\My���;gqo)÷�P99k9AI�	� )������hx�(W���-��|/�����o&�!��)<�����s��$ij�˺M+R��X��l]���"Q�ku%*��at�u4�
�c;���4>���oo�8]�I<KMR��\��<i�*���}��-6_bT�3=4(�@~�Q�ZX�c(m�D�}Z5@*���]� �3/gXJ�?���й�,�`"����BΤ�<,��ʝC���?GuG�4�}���4��Qu��N����H��>W�%tϯ�_{*7!�����r���hG�(�Y��V:�"!dЏ����$�;o���>�,8�71%
[6	�����9�@��Ġe�4����8��]�������0爑������o��`�X�1&�w�m"Q-N6ri��:�s떔�N��h���vz��N�V��~�Ϻ�S^䁌BF)Xav��*���q�Z�:�9�����?wS�����4��	�<_����׾�3NF���a��m��^��Hj_�rL�/�J����_g�!k3������?46F�c@��0`SL��TN2����v�H/8>Ue�rpF=�K�:_m`>��ZMJ�8���=�`[�ꈤ�+��&�����+�J|�609���U��RP��5�͑�c��48������H��_�:M�S��o��)��nu���&+�8�^P�ȅg��B��v��b5J��_d�N���=>6�S	�R^a��t۱7|0�]+<&��Y���;8j���l8�����za�*FaO�~����`��+	����MHK�B�ڕ�^�t��H��� dO���oam_��B���݋�̒�p����ʋ��^�曡-7w��;̡F)����Ly���C:��H�/�_K�D%j�@�#ԬJx�r�l�ډ�ř<�ݲ�G�$bKFo��U%�G(¨~ƶ8��(�hό�E3��w�A!d5\���'�<lD-�XB�2@�vҶ���������ǴuB/Xl'K�r-�&斪�ߡw,�g��5^|ˌaӜ �c$����.%_S�|�����c���<ec���44��������ݫ���kMM�M����S~ ��`<2�;�sx��ύ�`�����<�O�Q����v�cs�[[�g�_}�q�wQ<�C��\ul��`�6�����_�t�,����`l��ƚ��R��S�L�Y�<]��$�6B����=+�
����D}�u�]-H���tcLWˬu8Q"�i5��A1�Pv��izP }{���RP�0y0��h�I-F�Z���m�Ef'z�6`S�QY}8	�"j��:�e�i�YG�=v��B<���RAm��O���G�9G�
l��~��2�U�U	�tI�r�z[�z�G�3����N�ų���Xi^w���{�`�a�S�Sf�6���5@a���Z\�a���C��Y�0>I�JM��/��֛f
��?R���-eqV��Ac�9o0p�8�W3e�MeS�!<��0���U`*m����Ar��Y��XlO>2h�}q�/�IC���s�/4�#���$Oi�	��\/e�e�kQ!a/j�:�]2��p!G&�;��5�K��#N���'�fM�MǇԁ���h�v������د��G|���'A��Q��/]h$���W
Ёϕd)��ˢuӀ8c���Ƣ�mjh�D�J|f��L_<$�����Ӈ�L�Qw����r��o�RJ�]Ύ��Y��4�n�xF_t-���F��Ͳ�[J���J����#_|9�OA���J�g�8o !K�u)Q]��p��V�q�c�H�I��Xp�,Y܎��*��&���gͪ掻+m4���6���_��4��$}��Q!b�f�$<�s_?DIKGK��螏P|Q�h��t�Ru�ϝ)��s����*jD�xW�u���ԗ��rz�����)�F�?�qq���'��0�1`X�tS.$
�E���B3�{��.�kl����"��T_��@�W9�QgT���t��x I�����Ł3�PH�����/�v��}ܟ�4м���Z2	jQ�G �m�Ǽ\ò҂�c�葅�#��2�⡰)S�3��x;��%�����iS��j�14�!����4��X���^����D�t��leE�?=��7 ���j"���:�x�G��������W?֨}�J6����xJ�3E}T ǒ��\��h����P��A[�U�P���u�
u�.�_�o)7[Y�&���I!� tjk�YȆ�¸���ݛ��/!��h\���,����;�k ��ܒ2s�xg2�	\��X�e%!�v
'�P���0�L� �2`��2����WK���z��6�Q��ܹK-�wMpһ��t{-+�fHq����⧵o]p��_V�,���k��W���wH��"u���ȉa�D_1���ӝi��7H�����BxL"m��� iJџi�0�r�~(�+�&�6�
�^��	^ �H4�J�X���b�֙�B����=�{#;#�ɍ͕&-f����l��+K�/��)(��_MCeh�s��8����Úr�zV�$�S@�O��4?e~��1��@�q�e^/�e��'��ZLu�5{��.`}�a�ܽo8�J)�As��Z�Fd5\T��Lkdyj���!Ѱ��µy�.���OD��f�鑌P���)ށc����Qں��*���h@��F���e�x�[�(��*n�����nۛ��o��3MF��K�M��g��-Th�έ�>Zۏ�������s�>�W]am@:�Q��8"/(e��t�ߩ%u�2^�]����K�����$Fv֤0�cM�s�;q��rRd�QƜ�_��'�dRl1%�!�(�/�ʃ���d�\R�-T����-��W�яü/a,�b<�x_jl]�;���,� [�z����壎�{5ɯ%�$�1�?{�V�7�us�~j���kE��7����Nh� ����v^���kX�����X>^X<	�0��[�\������HfKV�U5tJJdMdby�z�_��e���*��������}4���I�k�扱���y�<�
�]�1�9�'��DZdG���{�iN�F'0�Ű/�O�ч��,󼴇�\�I�s#��^�"+���Y�nz( ����ډ�aH2��f:�ٸx��h'oG2��b��x�[����m����d���j,NB��Z[�_�*"D����v+,^��xC�K���#�WK `�!��/(jө�͟8�Q�t~3�*�͠�N�j��0�F����;2�J�r+��L ���۴p�J��F�$�N6��	�����"0�ǿnl:.:�C=O{���(���`�I�'�/���1�H���o7�TG��{4�������Ɵ����l[��)	SL����vjp���P'���ƬI�\��"-$�]�(=��%�x	>���yDDZ�k�� H4�;t�̡�8��%�]�;~s�wes�a�9��ood�f�*Rަ4Gz��� ����;Z3���h����/��ws�	�SÂa��uM	����Wi����y��'�D��x�&�"ŷ�!���y�;� �A|���pd-�@�O�<�� ��fu����O�}����������%�I�FX�K��c�I�3T�fK�ňC5���k�f���@N�:M�Ϣ�3��(��'�����d*d`�|�"���h���v3�œ�O1ϣ#n[��ǰ�'Ě��D�_��Ұ�C	����e�g�m�-· Y[b&���)o:DU� �m�����p��梣�.�q5yZqu{:Y�qA�T��"`3��I�z�w�/%���@6�\Ɨjps\*����U.��c��������{�;�`'������ oa�1���f�B[Dp��寯�V9ȧ���4.Rʷ!�U��0�������=@��<�����,����\R�Ua`�q�����|��,}�s���t�#��*�n�a�1�f�[@&R�%@�:�Y�%r�,x,���lD��fT�y�p�r2k왃�5"`�bp��"0�ε�����/U�שH [�\g����,�7u6�Y\��,o����x!;䒁�9�)�f���ةb��G#l�c���`5��JbڳkJ�9�h��(C���J�B�L��-���lQ��ի�8u�UGM;�1����|H�k��1�
rɣ�1�Ȟ�X?a%΋��st����!����?��:��oQ�K_̎���z_�]�� 
��l%���
�ҍ��+ߥZUY��2#��,
��m�[G��"�oYN���K��EDɖ9��	���+aNַ�%ǲ�ktA�C������Ǳe����>M,�sC�Ι�O�!��K����N8Vp�̗�&"b���������r=�����ڭ�����5mx	�6�K��5�������l\����q#(�T����(�L�t��!��EO��^Es�"J6�E?a�j๦�{�]Nm��l(����T����`��I���ʀ�.Xi��UF�Eߥ������k�?b�x��pR�bJ��zX&�$s��3�Đc�>~g�i:���������-4�@���x��������APx8Ԫ�xK��*߰�Mſr�!m��ˇ�rr�F�pG.V&1��qsi
�M��u�b�LR9���n��7��� �	��h(M�$(���n�t9��ӿ\�Я�w�W�
�!��U��2R�L�T�?�Du�`R��*��>�x �$R�{I ���J��G�
u37?(f��k�ˌ=�cb�I�=��k�=ӗ}���\:A\7�ߧ�g�n�Y�:���Z�(��p�"���F��v{%�� ���V�?\�<�Uh��o�U�;�V�Ȋ*K�3�Ls������p�I��#u=�Lȁ6,/�H�Ƀ!��uvn�h��a�ۣ�_&N�ݻ�W� 𪼛-�AŮ�^�`E�h&)f�k�_w:�r��F�<i ;��B�)�"=8�f���Vrr
�Ί�>�n��.f+���y�.��rGF"���i���[`�uI��)��ob�F��Ø�����;����^{h���L�AT�-B��m�saP
��e'���j������K1{[`Yf��լEy[�����4eɊ�u��-|�}"D�!!4��7�:�k�P�e��+7�|�
�0i�-*+�d�.s�c������:/�_e�E;h}742����e�4x�)Y�O,7�%��G����'v
F���'��Cs-g?����,�k+���z�3d��+��e�~�De�zP�� ���Cǫ�5w����t��R�[=��7����A
5
r����k1X6���[��7�'��3]�z�Ï�>������3ݜ%@~ht� q$��b��;��L��)�XM#@�Ȭ{r>�ʈ�̊I,��n(b�q�w�	���*G�.�x��A����p�U�
3AY����'�v��i1�\���!Ѻ#Y�B4
�mJk��b���VG�-�?�I��x��B[jgl���?�Ľh=;�O{�~��,Խs��j�����*Ȟ�]ۘ!2r�/����f�l־I�^D(k�#m���Ԃ�&��CFJii�~q�±%a���?:)͵1x����7X����\X��,�#��ߪ�8�Zh����r,��j�������&F�Y��,Fd����Il��������G'>�20�O��#��JUb-%�6���.׋��I緧���%	��,�R�3�N��Y�'��h
H�L���`�t� ��`���j�{�k����w��c�Rf�
�d7S�t[�{D�N��%�0o��2���F=f��2���z���{�8�ً�3=�@h�y�uuqK����=�����L9���;���"�/�2���6�!��ѿ�v=�f YP�{�n5��
���7��=AS���xT���>�c���F�e�[�S�n�i�;fӕ-I��֡У���_��:��b𙁿'6��FG�k�o����{7��j��K[1h\�a�Z�ït���Z��r?Hy��m�R���//�|�vrYf���>��]�3b�)�-"|�bT��������Q'�yjA�`��s���5L'�܇�������w	�$
o�zz|��Y�KזMt���~^��jȞᖡ�F.�ܙܽF��w���ө
u�b<;��uH��8򝐞mF�ᏺ����)�
��l&<�aq��g yG�<�F>�����n�kE�+��wZ�k����5c�P'F�EG��<�q�}��Xni�q�YG�(��y��1'v��i5���J?"U��8�n��ltze�㐙�'�����8/�����Z���.�����O"i%f���0�q[M{�|)�]�)L�D[-�T��Q|���蛖�������A@X�M�F��67q�X�9AX5P�8��1����h��'|c�"���#�o��k/��h8F��Sb���&r�O�Z�ھ1wS��I���+2#q�f��>z��L�:�t���T��4vg�PH��a�����U�^'I��ܛH"�je�k�2�XSGUxM�[P���).�� �ֶ���n\�y;I����J�tj�E �>�M�ԍQk���*Ӭ��?���7å��UV@I���æ�o�h��dH[@�FRZ{�˰T����م�� �L�lݵ�pͥ����6noݰ����f��btVc�N��%��;HB�\4X	����Y�Df�\ޣ�HR1,�i�v8(+.l��Y���I5���O���
A�����t�L�75��&�O]�o]��E	3�T�+��"\�7gB�i�̯��*��ˡ�D8��A�l��ӷ����p���"�3���� mCl����q��x@%-�o�zC�v�t��M��[ȃ��4�}�z��W���pe7��Iyhe2�?�����%������%8a6#C[�Ϥ�/1�[2��=��i�|�>���g(��I3Å���6U� �Rsܤ>ؓ�hz@�Dd�Q���tp�!�NbƂN
rY
(�&��1&pvY}M�pg�I�����dO�����T!�$�xg��a�q�0��L���nH?��^�χXr]	� �\I/�NK�!�T���B((�2v���������+n��w�j~Vmh4[�y�Y��BX��V��4��Po�bG��+C�y���޶qh�@�OIy��&�A�*��J��~�`�k��"�b�>5�����k2�~~�)ޞ)/Sw���I"b�����2�1fЦ���S�|��'F	��NL�81�m��e��H�p�&Q���A	'7��9]@�^�:0�\�)��,�������`s��
��/�,��!��l5hS��j����Xﾺ�u8S�,��&\��$�H����T��	����d{�lD�\}]���.;qh!<�"z�;ua���H~������u��I� ���4�?��˦����f��
��t�f(�q�fB�*�8�kw�B;��s��������� ���j߳[�)�0M,(��A��嘱:��FSE�6ݞH��#O�Q8^��32�RjڒB �V�~`	G�6�@v�g�֟�:�q��V�A!Ć�V�r��m���14x��L�N%���-�\K��n�b�V|%C�%���G���B7�L�Vs����"��q}�L�X�ջ���]bMx�n��Fy\�.E8���"<��� ���d����I��E 0^��v�"�W(
���� ����s���6�d��0���ǌ�$91	Y�NR�?����>��;�	�O�]_\��la;���"Di3h�j���k̳����	��W���Z��P��*�.��5��I�j���׀��(N�7���p ��:X�(%�[Wm9]�o�s��9<�Pn*�����}��5c��G��r �cw5�`��/ z�)r8�䁏�v��ixU�(�Z���3
��!m�*��g~q%�"�n�F�2�PO�.��NC�]�f��}���:55s�wkd�1��gA{�kQ?"n��%],`����pXa����Y&쯫��#>O/O����X��J���,eƼ�����P���>)�|�0��Q��2?J�Q�U���rns(�t�)w��#rR�k6�7	ž�/
/���cj���`�����`2'ؕ��p��"6M�U1�xFT��1{�;o�n���X&F��I�?��_ă��X���Z�yh��MnRZ~��7,���-VF��*n*!���%�0��F]��|����F�}���b�z�Sy~�����_�f�.Y�[��P�/����^����v��{����W��a4�ts8d]��ր�>��y(��(�0*�u6�d�a)!����x��Ȟp���c{1�?^���CL�a@#��8��POP��~��=}�v����y�H�����Ez�sͳ���)��Ef/�6�9�E!G�E���>��_2!�,�,�n`�NP�g
 p��K�}�F�s /���}=�Z�R!L��+��(���h^ϲ��e�Q�ç��Y�Qr�9ΐ�o�j��I��I2f2n`���_�e���j���r6��{�ys�\��v�hm�Iy%��)g^�o�B3x�ıV��ϳuh�@5o%Ć�'�] ���$��֓����O�%���qo���(+�g�d�w+"�=GMf׊ڀ�6=0�B��AK�d8)�P0�g�6�I��Nl5�d�`�9�	۪kP}���o�=��!���5��5�y�&0�Ό�ʦ����Kf\�����Yf�Ld��W��l~1`�"'�����*
-�J��8��?mn�#Ds��r���&�R�N'�DѵH��"3=�$훸@[N僬SZ����S.�&���]�5z��%��=��@<���/���r��j!�C0��T_��H{�\�$�bt=7<�CA}���+����Yɘ(�x��o� ګ�e�א�E,cKRO������/�Y7i=��fm	a��� ���T5f���C� ���M�Xш\>2�R�Z(V%��{!� k��1s�����<{���o��L˺>�~2��P�EQ�DC�ۇx��lv����!+I<�r0%�v��g�p���z��U�{���NZ�kO�+y0�?}�g~� ��\�b�Or���oک&ag�*W��L�3�y���n�,�o���}k���_>�{i�\X��P#��z�wX�j��!�{�]�m�F�m3Z����(�(�~�p�oM;�,&KG7��
�[Cd
4-$D����К���7��hM6�Y�ZG8AuSꡊ\ο�K�?�[|f¼��B3,�fz�	��q��py��n�����L�"Q�N����%3(��F
�謏&�.;�f�3(�2�&�a��ZQ����M�ЭJ(K���G�3�x*t̀g$:��V�R-х�EO��GW���/2goX�D�D��R�Ӷg�YǍ'�g�E�U���kHzM0�`��ޮi��k\�Xt04��v�3����ߵE'�7R�a��+�$��%��b��O��SCr��K�R���F��I��i�^.q�)UqWgs��� ��`&�H�����l�� ZãD�1e��G�uҁ+���Inϒ���J�hFBv�R#:F:��1������Z�o�+q�0����O#���F2��s4H_z9���D7:7�(��)�U8N�h��A6��0_�k�_擏���q���hd�J����T�Q�i#�KswjǼ��Aaf/g(kTl��U2߾�����J𰒇h�.��tp�0ܺ���.|�?�����V�h��F�P@�O�b�s\��W���Gi]]KDU������F��q�-�D�
2$'����Ҭ��#��l~S��T������w�7��/Ww��1���`���۟ڎ4��DԖ��J�̙B>
~�T�j:�����^��r�E�F��E\8M��I�?��}̿l����N���S��̌�@~�=^.� v��M�F����d���b��b��m"E�L�_�U7�d��I��U'5<J��VVT��?�d�Q���_
	7e��K���W���������jiŔo{=���G>��e?s�KZ2�r~Y�JA�?������<2��vC��U6���ma��ZI���cB+�4��+a}�J��o2V�b���p��y�UG8l�x��f��Ycu��������8ٞτ���2���6�Y�r�U�vum���yjE���F�U|� `�4y�Q�_-K���m=/o�DIF:OL�Nq��n�П����њu����%��b5�@ڸ'�)�ACx9y�'���@�8�]q����@���<�K�¬�=$�Ƃǉ� ���?�#�ݻ�x����`Jqκ�%]��6���kl?􆝎x��iLl��0f�Ҭ;򼨳;�5��P@*��8��ִ_SV2�ܬ��s��"'�(��XS��ל(f+�-g\M�6�>ᘽ�6�5a�G��Ӣd��	�+�c���#Mx�AwZ/�?�
'e��� �LF���. �t�!������UD�oG�� #��,$H�|��^�e������_vכ�ct��;�8Q%ޥ�?����m��5��Ơx? �,��VLr�]��������):J�l"�I��J�xt���
�#�q����6eر�b/�*�q��Ȝ�sqWN`�6�����P�q��d#y�K��h��Rs	L�Lo&�B��~�w��Fq=�F�/
A�VeQ,����.�SZ*��v����1��s�hl,�8�1���xyիd>�_Ä���Mf��p��n[WT�)��<�{��>�[9+!��ު������z�-n��o�%A�D�oV|V�MJ�yS&���Gk`׍�3��+�vl��Q��!���(l�.F��s��ԫ�0��qKx�\���b��l�+?#tf�=�LFM5�R4��}�͈^���t.K��OGn��v�E��SZ��l�L�F��D�J��÷@�?���d��3|����[p�����tnEI8�}v0�+�`���,+G�e�*)�%��|s	Q������ݟ�&-k��M�Ms�c���
[.�萲	��*<��+$\�T�]M�a��3��{/�EaU�+�[c0&:��5�uӾ=�+�rI-�T�F�{�̍�R�|��y��Y��Q���0\!��t�ZҨú�%�4%ޛ?^-�D*PQ/4�"�i��ϻ
k�[a��ѪXc���kC~+'�v�8r�p�����Y�37�X�8_x��o#��I���U�0`�ƕ䡫����{�nm�L��
{Ͽ������ٿ��1��n9?��j]M��߇Xb0-�t�јWĢv�c�5"���MqY�Ӻ���嶎�$s��k�n�i���ڒ�|��1fB}kݻF�0ggQY �|��|iЁʛh؟ѼH#g�;�m3���o�󻫺� 	E�t֤�
�R�b���ʔ�C-���)�l���r��Pr�jZ��U⥃��mX��ҢH�P�=�G��W���"��<)s�{0ur�10�U/�;��`�lGIx�Q�J�pH���]u6�XZ���D�L̖<*6���#��wA���ټɞ=kݧ sj+��^�mz,��v��KR���3������5S{����r�ֺ�g�k�7�S����ƥ�A��f��	��� ��� ,U�G�V��~�W1�3zfȆ�?�P��[�����ۧ��(a����!�ܞ�(���-�m�7��G�C���&��zQ���|���gA�z���Z#h��i5E�XƟ�p�sW,�6mɝ�q��Vޫ��%�Nj���	1���?���x3<`G@;^<u2��M��:jx��.�/FقnB�5�@ePR�p*��\]x�hnP���{�倴�����^�E~��<�rk���Ē�u�#U��&䥸��>���	#^(Aյ�?0�9���.*m�����OL��$��TD�v�WwRҏ��/pP����������J3
n��Lf�ztR<�B�8��z���vQ�"�@���Տ�f���Ѱ;����!D�~�#F/���?�(�f�����T��%jO�RY��KS#M=C������ o����E`3ڜS�q7�q�6}���T��V�?Lu�W�_tR�*�`��r[[�Q�5$�2oջ��b�T���(������,�-d���m�@I��zB2��ƙ���O����ߔ����j�/���%�=�H�5Rl�x��i�/�O�hT�0';���~JE:�u��@�v��Z&r��!T�t �}[<1����=n�D��A��U6�b��>(nwZ͝��|3�݇:'d�k�i����[j��N�VD�����Wb�w8� �<;��^�΍��ɵ���+C%��"��Fi�3�t���),95�gk}�b/s�o��j���"S�N����Z�w����(~���و��vY6��Ǧ~�g&�9��e�Gw�~�Ў��Ҥ	O;&O��8��B�����[^�`i�d��`7af���}��Y�D�`���}DUY�6�+X��/�]�1��k;�:�T2\�X�"p$�CF��}]�E�U��Y�!��DD�
'��pƨU1�:���y~$�^���A1j�U���n��ax�އ)�8q�Oys�n�k#�^�F/� X�>���I)m�8l�����X&�B��fC�k���RYP�zD*����+�-�߁��"�L����뽾a�^���c�W���s���b4��8��!������i#���mBF���j������O����g6�2/M��S�Ā��f(x�#��]z(�vH�K��^��Țp���>	q"�#�!8��(1����G+><ރzc��R1Юu�(��R�}h*j�����ڎ�S3�8	�kY'�DlM�׏�Z�����;]���	�,_�=jp����R_�|CҬ�(n,-�����9:bT�7��Ʉ�^���n�(Xj��^���
�p@���`��khGʰ�I#�N�M���N5�k���/�n�f�]�{\�n|�c!��t!�D�Vg����~��xi�9�X��
��U�w�1�?�d^闧5&���(��Y:�-p�7S� d`���>|Ѵ�z-���=�����������`a�q�QL �oSe�E�H��4{,	��O�z�F��Ks 6S�2&�J?���~��,�_<��A�^P/��Q*���D�a7��%y����掖�w��a�ܪ=��d~�0�3d�0���>!ܾ�[ҷ��xG$�a���L�mMf�P.�-��RQ%�k��D�{�o?^jB���R`�D`�-���s��=�0�����ty�$�����!��c>qp�KX�iWUp{ﮅ<5�ZTfh׊���oW�<�T/bW��Zr/��+l����ږ�V��kCCkZe����9�|&���0%���.�S>o�x�#E�ToSr�N���.(�J7F�)���Fޢ�V��&`��,��g3|���&.S<{RjW�"�'P�h7��N�K���wbr�-��=K���1n���I�Ue�[Hb!%f0kB�����<�)f�)_�jBsM:`|WA��'�xNl�����i�o�����#-����1�,� /����[k��t�g�O��ݵ��%���;5��L��6���W`��\"������fa+[}��[d^`l�˦�i�U;�wR+���T?*^�XaCF������^CwaX��'	�n�W�E���rU��z��۽*.B+��v?��[caʺ�L�}��8�T-��e�Ӏa��0ʲ!�J��P�Ħ��T�I��4v�o����b�M@��>��]&F"�	�7����3{Z�'�pX'V�B���~
��=t�%A!b[�w�Vo*�q��V3�O�0WR��u�h1Θ��C�<��]a0i��|��=���b%�8��/�4���:�z��%��0/�`��Qwћ��+��E����������޿��C�sW�uZ�T�F -�D]���h8�
p{����Z�v��S�S����	)�"�����ǹ��+K�>��@���Ϳ��TR���TqWy�
І�9�+*o�qά)�	)=3Rּ/���%G��=Lz�՚G�A `��V}��`Ռ,VE��V:��s��*��E/a��n(P+o�;�k�ȅ���h*�n������PԋMǠK`�\�֟��)y*�/��p���.���v��omc�6b�R��P���ESR�ӎ��I�ʇ BWt.Ώ"[q�&i���~��o�;@R:&dֽ����qW�j1�=���%�Zqb~m����P�5'*��ê*�l�ڼF�A����̈�@�00��^C�,������2����}賩AB�OJ�3r�!Yus����9\\�����5�D���2if��F��u���z���~�ڹ�S���j�K�|��R�T��,w� 0 (��ٍ�}Q�/��N'��A�t�~t�����s �g1�~
A�ơ �/y��{�c�@�]q��(ni�!_=�ѓѝpLq��c��No?ʑ��Y�B#�B�C���8��K�{��׬�~0��STo� %���+=��[��wxR�6�]@b+ha�e�7�6��u�%�$�OƵ���3�0�}���J��}/'�Y�04���Z?�;"�I3�9,2�
�B.䶱`�q�P�J��O���7B���i�:S=8�G�u�9B�:?�8Z�K:��V���Ü�����Y;zk�ן<_\%���/�`R�ޔ�zj�W������0�h�ZM��=!��j�ĩ0z�W4�t��]$��x�0z1w�uw[��`���=j�U��|��Х�h�-�((+u�[:Mt+R�*���6k��W+5+���.R����#�Pyg+�I��p���g:�|�Ό�ϊ�������)�d�*Iw3�t
5cvJ+��C�F5C��ۅ�=nt&��A�'e$�U��5��)0ѱEtn�C�Ү�ٷ�}k�r�H�h&�O:q���Qq|.��Y���(t���B���ۉ��O��s3�eq+�7���� /qԩgɑr���M�!�S7���¹hB�&w��ߪ5�I�B�8��o���
�y�Vb;E�o7��v��s"9~��T��X�w-׿ꨵ�w�$�r�\��0�����ܺ��]����_�䳠��BJ��m`Wo3 $�z�NEY�~�ID�6� �9�>���,RҘh=1]�0�\}ٙˬ˷���JY�!��|���/���_߆�u_�n�+zآ���D�T������k���2}�hr$~��F��!ڎ!��{�O��1�
a�̢N3̘_�c��0ï��Q��7��W��C����J �F�擔�@@qy3�G=yq��ϊjL�X�1�&G��t$��m]�p�$@�8��9������q������i�le�(w�VM�C�>��mSu��6��<��� ��<X�D耭�*>���';����s�#1��V~�/@��j�iDD���*�;q����w�3�����w�g�l�+�Md �hK(�sL�,PтΫ���R9W�	l��@e%���c�B���`����b��k@$8�n.��pf�+��9<w޴w�/ێ�:�!"6�sGyF�x߮�r4��s��!��%)%�|���A�(?�#��b�8TD���?�+�j�Q5
j+<@���9�=�A��i��8Z�d�)'��*��]H����`c ;�� �Ϋ"o��V�5M�G��b�z�(��Cr[Bv�p8R����s]Y��7��e#�����R=mZA�U��h���Z΄��Sw�����[u��U�� Z6�$��c|�. �ת�ĕ��� ���%	+ϕJ ֐��{�e���EmD�H����l��fDg��o�os��X�ȳ�?�Xu	��������|0�Ti���+֚����R���_�L�� ����Dlc`�J�����1�|{���Kg-�p�U����w�Uw�3�D��u��5���b�ݺ��4:��ܫ��>y�l��E]���9Υh8}��O\Ԑ�U)x��UD�	_�Ǌ�g���ʄK0پ K-t���T�����)��Z͔ؐ��t��X$��]����tLb|��q{��N���(�ϴf~DZ��B� �F/v�bqn���+�w!�d���}���k/%qJM�������T_Kw�7�'��9���a-+�m������20�VlT�c*xu[��R#[�l�cKM�1��������Li���R
�ه�t��SÏ;&Ɩ�x�Hf�����t�^/�Xa�m���Ʉ�C��Ƀ���K�C�d��s���	��&I�@N~ѐSUN|� �\�"i�!ޤ�|-Q�>^
�r�@��4;�����З^���e�\!��~����RE�M�r�9��A��mn>�^��aYm�(Ĺ������5Q����o�ނ|���ِ -��~U*��x��.bZ��ad���L�W.�;�˥V�}64��ġ�K�#t�����ID6�ҐX�q ܫCӒ	)-7#C�� �x�N��K�"x�(t��R���t侑��٢0�q�D����:m�5&��s�����u���� ie¤b��&¼�����1[cF}��{�g�FaqڳB���O������8��"j}$I������![+�X�I6�q��ץ�{�2�g�)YZl�"�ߓa@��������	����~���J'�Ӆ���; M<W��*.���>P#���#]�6R�H��� L&X��l*[�O$�ːN� 饷I&z �{���l��p����'��tb���D���*Ny�A���gQQo��pD>��B��tپy�����i?}���YV��hj���=�m62�۷gU���{��!���3���.hբFAU�+[tba�,�^�d�%]���c|ê�1�n�D�G�6��<��ܐ���~����M��v�%X˵X��t��������$~���U#P�K��t�^eH-U���CA~H��]���7��ޯ)KY
���(�1g���=����E���Ͳϊ:M���݀��7=e�����S��K|c�2�sW {��/�V�<`����$�������NY�D���,�Yj����pP|p���|�as.���:i`�\�8�X�R�=��G,#��UibM�fT�fh��h��͵���`�r��'�yKkG��_��o��.�j�?����a�W2d���j���92��MM!�(w^?���=a�c����,�������Fo�^���-T)u�I0�v�H��yA�vS���k��F�Z�����@i�.zΓ9��r�l�
p�P�s�ܙ�
Z�n��w3V�8�U既!�k���w�6��׵�l!��M�1�kgȟ�'ӽLB�Epm@rr��O����~BEn �8�����[���tfD��W��V��^ǎ����k��}�tulÁ`y���	�.�BW^l[��hr*D���Ftw���*�[�]x���v�N=X����x�[�1Gg�c87��ÂB#y�Oh��Ӈ���U�&��ϸ�S��
��>^�ڦ�+~MN�h�o�ˢf.yT-2�Tm�N�O���S�̨��le�%H{��Q��%�����U�Jڞ�ڵt!]{�8(���
w�w��b���z}2W1e��9��ɃM1qI��b9��3E�l^�_�gDԙ@���㤰��J觞Ĭ{�K�����[_��ȕe���T��&�ȭDG��\2�$��l�t��@PH��y#p�C[c��e���.�]l(����oY�K���j��6xp;"v�ZB��0�7rے��TZ�?���f��� ښ�x�A��ޢA1*�n��:������!��������"b��fa/�0���u�|�g� �wm�c�ܐrW����ԕ�0�dT�׷�c��=8p�1Z��]�XuJ8ye���t�, ԕ��i\l��@]�ӷ���{r�m���?5)o�������MLij��v��|}6@9z�&��GZ�VӑI�R6��wY��M���e֘�5s���.�ۏ�x���05Gj)^*�.�4i@~K>�Όt>���M����h�@bvP��,����-�܎j^rF"=��GWK�1��������ur���s�~�i���-���)�&i��������r{�RژG.Q�ۅ5U�[_V�7�cJ�s0
Dfc[�T�4�D�'C;�����ϴ�]�َ�+�G����&ݥ��ǘ++�8d?ؒ"ȨS�d6�_�|\�!�\��Y8|��D� Y�b>�lSѻ��:����s����)f�
��k��?}�ps�m��*�"n�W�Xk�:�Ko��m�/��4N�uVV�bEtO�6�d*X�q6ծc�C��vj�I+���10��4���<t5���F$2w�J��R��;v8ֽ�DX�Q� �Un���W�uq6^�_zɅ�ķ��a�q3A��ӻ��(2�C���ݧ��w�z+��1i�#H��m�|�]r\NW�Kt>?����Ƙ} �~N� ����#�`d�c�d���e�F�4�e�����uG<��q�\:'�Ն�^2��{~bM(5R��X��ŔQ�7��"��»�5ظ>��s8��������cfL�.��DF�tKzV�����h �� ��m!��U9�*$��,�d�C��c�5|U-�)>\��2��u�n�u���cqGb�?��3���y�%��X�s6�|���3."��	塼���5�/���x9���4}�9l2���n�ql��8���nAo�u[BĿ���4���L@�?	��:�D��Z1�tc�5tf�~�7A���]h�8 Zra�D���<*��������S����}�>��9Э���Fv�3]�TA@��'|�7π�i�|d��yv��ʻy1�;`�7�;���(�I��������yM8��N��䢂�3N�Ce�F+5�Vk=h6$\,|e��#3�&	��:���@�s�^$�7_�	aN 7[<�@����\��M^ꮦ��k\࿒���km-v�6�u`d��X��dm5�t��
Hf�Ds�_����]��^NVa�9ͅT?�������|Z�5�<��q���5�Z��ò?.�D�B�3�MF"a7."p
r���mrp���3�9}s��|���a�(�[�(h w������g����x?�\j�)d���Dé�.�[E���^J���Q-�+�F<��nҫS��i�ru!sL,R�ӑ��ڼk
}�P�8�E��pC��\0旴O������B���ΨY�F��f]��[˕�%�J�H˝n��7<͡o0���F��
�As��淈�RD���j1�4�'�5A����ѯ����nf��VQQ��bN:���ֈ��/�V�ʹ=�(hE*��U�Lf�M(���Nۍr)Z 10�
�xl�eN�P#� $/�D}+b6��� ���a2U_v8^����Wۼald<�c��u3�Rt����he��,4���1�7��Cs�{��ɪ%< �p=�o˗�1#���k�"�l�>ό��F���w��N���Pxt��*�$�rgHE�)V.,��Ma}2��P8M�p�����kr��U⿗�Y�L ���R�N�I&�]��R8�Sܲxw�)w��ϫ։Y_~γb�m�Q;L@��-j(pIܩ�F���>���#���F%�~��k1�V<U�C��!�o�@)D�Wr���5�r�N,�L�آTy,�������Rt��g������ �~���bXM#�k�h�9F~�-�[��ve���g�^!��\��8���i08��b-�dFց��T�7064u<	Q�{���)ݲk�ۛa1�pq$Z�̛+YG�1٘�/�ޚ`�Q�8$��QΫ�6r��6,-5��0�Y�.���Jo���P��]4��:yy��`�`o�c�N����8^���^�ʸ��(��`�xʏة�[M%�#�ƣf76�[�~JA
�|�PA��o���ܣ��LBe0H���I4w:fYe͈��r#O�s�N��>��<͗q��^瓆�@�^<u�30l%�hGm@Ꮸ�4�`����O[MŘf�� ���8�0�M��k�4�h��M�V5�7-s�C.�"��j��ۚ�Ǜu��w�R-��|]Ԧ)�ȸr?�Ru}��N���.���P��Mk�� �)-���7�Ɯ0Ufb'��-sUx�<H����"�g�M�>�Uc��c��Ľ�o�G�=�� ��@N3=��ý��(�/ �������i�ˏm%�L�(dP�����U�����Eׅ��S*��?�_
�O֣�ZyyAD��j!���c 'U7vԡ�f[����dD)����-���ιŏ�h�+Ej�Y�Q�$��df3lҖ�иS3C\y�A�[B�[��r��-Xz)@زFP��*0�db;h��5��{�wl�@���ٟ5b�r�r��\���l�?��J�� �Ӓ5�Tu��~��XeIm����tZ���PvͲX4��jȈ� Eͷ <��N���F�T��YI�5`��Ja�ւ7mېu 0el_�����q�x��� ��.#sp��2�w���O� 3���>,�sh1�WC�6F*8��!su#I.�h,>����4��,��B���g���4���k=��f�Ml��v����Ӟ2�U-
̥4���]=�5�\�>�Att��\�Щ�b���|z����MH�H�d�;�jK���ִ�7�U1�6�kd���=����vR厀^�(:�Q����ӱG��^G�8C���}2C�8�w��$Q��MK�=�	�I>�u��%�
������I8�AEA�/��xA3��k�5��81�䥐�4��#u4�˿v�
։��j���ږ�@P�9o{w��*/����A�}��N���+z$6��G�B�r���D�����	��:��>�5
�R��8��9nn�t�n �򧚾���~����w�C�+%L�9�;2w�c*GR����F�tQ�e�Rq��Q�v\�pT���ٿUN�aL�ޙ���l�j���b��t���[f(+
��k��^�&�Zc������?^���Ğ#
ڏ3WMX�݅j%еd��P�g��[�lXqY�L��}���.#�ܑ�4�է/�b�y>�\���7�/�\��b�q��4z�@Pu[2Wu����pr�Ai��P�i�%CZW(	'-�[�mu�	�ͅ���W��R�h^�ϝcaQ��J�o{���-�!?����,�4| _�/ōd�����7Q��<tﳫ��|�,$q�^�:���1�<Lg�?�uiuS�%ߐ�����J��
~;@>b�W��
���_���c����R������=���t }�)�;��O@q�i�ó��:͈�x	k�����0Ș�.�ݸ�s[�����O���Z�є��H ��m0[%u�P��'� �_	�`�kM���x�9���}�62��?�����y��6��yX�[Љ��h[�ސ�#K����#ܺ��!p8�vc���tn�T���Նբ�#��Y !���ض�U����������kP�P�Z<q����w�V[��y�ӿη�>�����(d�4��WU�s�ֶ���_}�z)�_!H�D���"6(Q�`��G{��j�k�"���:nz׿��v���kԶ*!W\�~B~H]P=��������?�+���rEBX&�hcZE?3Hh���\�`	E���=�9�î�ў����ҥ���"0Z9'�উ�Hc$�N��2ڕL� A����ƫ-�Ʀ�b����і��RRr)���#19Â�h�آH�*�;��Q_R�.>lU��u&�Y��b-+lTo<�޼��ls��!��j���!�Rr���=�����X%��`Jm��5����>�e����y�F�H�۳R`k���I�jFYx��%��� 9�vkv0�u	��"��[�~�����#ٌ�Q#�<ci ��Ʌh*Uz�80�w�ͼ8B��W�ĽqC��;ɟ�\褫���;t\k�s;+�c��o���&ش���)y��9h `W��� 	)�yZ�BRՂ
�J�(�6�w���Qօ�2x-~�ש�~�@j���z�?^n��Ğ���E�}GNx�@�D!Xwbb�E�L����gd&"�UlR�Ip�eJ7Ѻ��ca�9�
P6��=[�)ˆ	L X
�YV�
��M�����db���<S��;FE�p�D�V��n/�F5�`��4�2��L>�r�a��������ijŧt��X9B��%�^i�c/іy�l��G	
�L�M��Er�-qw�s.vF�� `J�l%�MdR����%Zֹ�p`P��8ccE�>�]�W���3{�)��"	�r>!`AZ�搸C>�%h����Asb�R��y�X�m���&<~p!I��6+�
`�%�+)�n����9X=�e���8���4n��=�d�[c���iX�лvI��;e�bds��8���1z x��rh�x��\�k"o�Y�P�cd�1���-(�OWX�f�&O�0F������qk ̋Ք"e�!�iw���!�q�R���<�)�w�T�G���6k's�:�����.N��-YMu�}]|OL�"t%�y�q�Q%:���/z���ø�pYl��c���H:���	Qm,�h��6S���
�(\��8,O���4�3��7�n��}I�A/&	-���>���U,�J��Z�g�4{���P�W�'�;Тo{ę0�H�5!�?����aǭ�ù��Y�,�Z��@�� G����Êt����Nw�;҉v���k��_�+�*���c�-fr�%��
���9i~,cZ�m����-�g���Dx��6�<��3��
q��@f}����I<�����
�Hc��z6����O.,��A!;�|t����-=�Ԟ�2\E��k 25�.�<kO�_�PQ]�.Ƞ���R�n#gV]��<�� .\P�`(+0:��(�����c6.W��ɹC�7������o�Nʄ
-1�G����`Ù��z�wXr/2�k(n�,�k�#yý{)\��-�p�?JS^���g�SY���@�,M��ˢ� �׏��? F:��@Ձy53|��B��Z
����{gGL}���H 	gZvH�M:?h��q���t%w8��_	��˚ľ*�F''-���K#h�'f���ﻭ�7h��z��G���{Љ�S��e��q��\�v�<U!��[���fw#b��cc0��� �����1�����8y�ާ!f���k�J��h��
�'A�E�i41��>�����p6���8�!�X�픊nn,i��L$�4V�-�'�D�>TL��[�ǖ]xNG?5g&�"�sP�_V�mK������KbްY{���
�f��k�%*�T� e(��~i�]��sl��>�ȩ%D��oC�"����Bl�AI��l5�tj�d0b2p��Kx�p0W�^N�x.�+�_��~TU���m@��TĠ���O�!x��������PE�'�V	�G��6UW�E�C�t�&��"�5��	ְN�� 'IAE>��wo3=W�k\������2ķ����� kI�_����w�`�Qws�3�@++��=�Jŀ�2B���� ?z�&�4��B�&����/�f'/��Y��|8��b��f��'*����}�'�*���}�cT���6����?7Y�7�:_M����}Ø;�\ۊ%4�e�}��˘XەR�D[
$�v�䑹�����N��+ah���]b,�vf@)bRl�z��ݨ��'k��XI��.�X@_"�?��%�����4
���Et�LS(L������X��<����{h#���z����v��x�Ү�����yKV�j�}9�;�2z�0���#����H��УeFE�p�$�X��z��Ez�
c4�V
Kl���c� � _�Y(-�@z��D��E��,�(�e_�0�ڽ :{�f���}ٝ�s� �O�8E�)+���l��6�#R}d����?7.u5�8�������v>!�U�:��X&K���A�阡�1$:#'-#]>�lZ,~����%��ll��D�4�:�	��Zx)5��g�([ǻ��Slv����B����+��2�~T����%�t5�O��UR��o\���ƞ!�o���DkIȪ���N�� ��G�����M@(MЙW[.�?����0���h��� H�C�D����ig(�@������O�h��sXã���isO���zHP@�`u����iR}��_'Xw��f�t֨��Qq=����0OqȨ�J
����h�S�|r{�m uo2G�|�V��GCYPde_Kϋ�;{�t�9��ҕ�Ҟ,�z��k�f+0�B@x�1������浄�<�gR�g�l���5+��r�ݥ����<�.P%�?���v�y����H�N*B��̘�wjO�:^S�h1o�6=���R�z�|KN�nn��S�IN@��O�[���]%�����`V:��*�e@�l1
T�Y<��a#Z�kǉ�r�G�>�ޛwQ�E�����4h$;������( �`�]��@�&�x����
�Wu`���ݙ�O��gbe
���.@��.)���op5�r".�ǗR��:L� �Po-sC��\ .5��Hk=W��S7�n�<�)6\��d���$�t�`tC�-V���~�dXh$���kܣuw��Eu�ps陯�>V}���'�>��-��|���|j���,��m��8�鐂dHNX�W<��-����s�P��:��E���Ѐvw�d��t�%N*�]j�?�(������g]�v��7�t�y�)�/�P(L��D���p�";tggr������K}�X�����+޸������"�\	'yx���N��WN���PKrN�H�Ġ��\�\[0SuR<.&O�m�U
��l�μ�uE�Bd����]�c-ِ���i�X;L�e�џZ#�
9Y�_(�h�ă�oV��қ&�ڧϞLы�����?�4	����yÓx��XÜXb,�e����uLٮv���~im�a��6B|�˿\L5�a�n�֑�SRI�߸FkI�r�&Bۮ�B#���ѧ�h(Z.�(�C���i���Ѳ���|)�9+��*��e��m�)M�iim�'Q�p�P?[��D��W ��[���0�&c������V[�z�m ƛ���e�^�V��諓�Y6��+,[}p���DdF�t�H_S(~]�q ��	S{��
��\��-�[�焪2�(\���z���y��<ւy�c;f�o�i��a��'�Zٰ����C�~w��c�Z=*��ִE#$B��HR;��1��e_�ؼGXO�ּ��׃�
|%�͖���N�u�J��9Q�]�ie��Ur��y��� !fqn��
}1��{�,6Ц��w�榤Q�`0�������a���^���#ԖTn���l���N�;�S�a�dt��A�\��8�`C���J|��lZ; ��p�pD���g��K��N�u!pH�gF=w�;8SaΉ��
��-�l�؁���RCC�+6>z� �+�x�����+�F�H�����u���[���MGC�.u#R��G[;>79ϫZ���K�e����
j|�rH�VQ'��l�-�*I3qc�����G��ԗ�m<0tevir}�o�Q�7ɱG��	e.���G�Zy��{���]�sPA�tp07�ڀSv5`]��*�B4��n�3��]@�+��@
��0��z��bNy^Tɩ�_x)Xl��S�N����1���!�պ�� �p��k�\�E�w��h23-��O*R�WH%�"��l�E��)���x��9��>��[������=��*��[	�
�$��)7T.l؁`'��f��*a���Zʠ%�Z.P��������RHF����E���2~^J�������;Ao|��=Hc�\Im`�W���,���Ӑ`6���A׫�<͊��5���qt�)�:�t��vJ�_Uhր3���W/y34�JG�i\<�7>z����� ��ة>0#��I�:�pQ#�O��F�?t��D���^nww4н�0������ΧC��4����(���n��1����������'��u"���z�a�KvO�!�N�|�뛳�jbB������߰="����a+�?8�#����DU������d�a��GJS?"�
t��v�y?�˨׳�|�ȅ�*/�}ءޮ+D�`iP"2���{  ﺤ���0��W���\Y������l�UfD
�j�8��?a��w��d��iJ��/���P_);"�ٗo�SB[P�U���4_�!��F\�h?m0��\�%/�Z,�W��ԫ e7��h������Յ�bX ��٭�&z��@���_H����h���G�C'�2�x�yy�&6U����#8g�S�q���h��,�7ؓ������:+��%�S�l�h�+	��n��GX�� �p��	?_�!6���9���:��Ug$*a�B坉�Dx>�1c�E���N�铦���u���XHVK��q�}�Ow��"Omv���\1�T�i9�Ljv
,n��Պ�
7LNgӟ�NWT��[m��\�v�����N`	B��]�c{��҇f�D��e������_(5P���VP���J4=�ň�GGC�Ҙ9�C,S�� +-aT�4�n��p�]pE�j���Nހ�F������,at�Č����é(I:�ֺ*���˝�ӧ|���-� �M��T��>N�	�y�����$v�)@/�?�*Ch�0 �"�g�����#*�>���.���n�u]��L(�y�y˼�K8#W窋K����C�ne�ׇT%�(ru'h�&֔�,����aAYpr��4[k�P8�*5aH��V�Gw���yłQp�jhl҉��3�f�y/F�׽�j�	���+nߚ[yE6��\�X��� �ƫd��nK{�|�Vt[����}��5�6v��9�+.ս���u��n����r���G`��~_���_�w^2О��4\�G�O��4�Kw�7���F'S5g�|Ϟ=��0�i�Oq=��Rv�?6�\�tA0��w1�����F���I��u/_B�����kYK0+i)`���>���q�,�5�;1*��!(������1A�K�N��LV$�$�H���B:�h������Ǆ�~�K�ħ���fh�I�UH� =ћvqy��b��|:&�iJ;�K�E����_4��Ҽl�?��u�W{~2�f
�-0��a� e�ݭ,�~涞�kq��1yWI(x���EF�È&�n���+�M�|B�u��>�~w/�eͯY��^J�������Y�T���)����C�5��B�����)6�S���J�d�����?�ԚSuǬ
�W3�H�&�1?��4���Mkr�W����O&"�3��_�یK wl�������ې�������:}\���BQh/��X���Ã�˫3e�DǺ`m�흒>ŗ���Yb&%�E���u�U{�1�U
������q�=uK]���ǰ �bg�y'�8c�K��"����׃&�u��#U���A����i����p;�s|�ҷK`땐��x<�ǚ��9���0�b��z"�#��ԌU����Pgcc�b2O���b�j�����A�K��l�� -!�sMXt��� j�i�v6f�{�k��Ku�V!*��(h�� ��8䪫�5�J45*�wU1��ݒA�f[���e�`F������r�p=�����J�1&�5���-4αٔ;��M�o����
?�{���-�?�"5�����^u�x��t 3�z��d6\���B6~���3#��$d�ZB��<;�#K��$��R3��|4���1�GlM��aB&���-ռ4^�kc�ko����I�q7Ҕ4.�N^&(�y���tMM>0\A۫_���19�|?�,J��udN��.��=7��e^Y�X#�eU�+�7wF郙֚\ٔm��$���+}������ߥKQW��j���Q 7ylM��]c?,ۋ<�/'�������U�!25�����y�N�y=H����<��S)-!�}�����P�*�=�L�]����(h���%1�M+ǁ�Ǫ�H�T@��㻕þ��d��kb>��ۅ�&jwō�ʁ4�j� ��D"=w�a������x�6����G:��1`-���ؽJ��U� 9����0��˔�.���צ����$�A�+�>yxiZ�Bت��uB��͔p�<í�l�̯�rG����+3
ucuɷ!���C݆y]Mv�Q]DN$��y��<�0��~���8�"I���ه@{�?*usX��abK���l�L�{>��gW�?��o�*��Dj��i�����3�zmJ4�eWHY+�}!���J�O'��p���x�&�A�1��Z(r+��,�I~�.�S������o�<��&�׺c����A��e�G89�Ǧ�a@�;Bp�\�q�5�bp��y1�b��M��[�۫qlײ���2�f^�Lnr����{9��D��z���[�����j��@  P�ѷR#,��jGr��.�a�MU�װ-��K���%�r����?&��
�u��ա��/���3���4��o��,� +	�U)ʋ>��}�~�Ϻ���i��@W��9ı�3� <�F�K;�q��0��^���~���>5{���D褴�~�i����S����]x`��K�]�a���7T=�)�(�WW0��k����_Bu�^��Gmc�3�{E�C٣�v�F����D&vǗ�J'Y[��	w��b����1�K���M�$y��f[����,�%�qΔ�߮-o���B3��P�����m����Է�"��n�F��VVqsK!L��/�5GJ.,)i���E���h��ͨ��2�3�կ6�\m��=D���b����]��Ȥ�3 |�DY�j&Đ\�ͺ ,~�$Uv�n8��+�߭S��Xi�K�6��)�DTZQ5A�]M4�#����]��0|��}7·r �F���7��g6�Xp�{#^���Q�N}�$����#��2���g�|mH�aB���L-�~c)������٭���N�p�_Dܶ��i�Z�{U�	tu��IE�}FŹ��J6�W~p��ȹ	�����g\�ez�]�=��^7���9:��������LF���A�5Vx��܊r��<�~��G&��0��D�lx?E�n�9�}�	r,'�xI)FK��J'��bs{�Ɩ���	墺?�1^�����$>�8-�]x��x)�%��>ꋣ�&�`�� ��է�fYs���8g�i�`��1ʔ�y�8��q&��*���?��B��	�vN&Ҏ�v����5�u�������д��D���~G���G���`��=�
�3	�à�bŊ���g�-�y�lC1�.Jp;����6ꕆ�&H.3@_��3�Q������Q�!���f����Ҷ�9�{�x4O���.�y�R�pv�K�$^ʛ��Ӡ�Ĳ�F]�it(�k�?���i��r�JY�erq0�;�G���W��s~����ʑ��	����O�%Nsw?6� �ax�N� 0��2��Z���~�  ���
�T�xY��y�����еS�'�h0�Or��j�&7�v����A�����wQhڲ�YQ�9D���N�h8���^�<�+�g��8T���s��JG��͠�'�$j�D�f����KP8���>!�y���ԏ��:�8�[GJ�w�'գ!�z����\Ň�Lu`����S�	ZB�^�rP�*l�C�t� @17�.i!�m�6	w	�-��)Ua3㒝�)��ޓ����).VQqwY���bO�x�_��JG���ȍ���?I䙛�l���ɰ��dJq�2�<3W�Ç��%%� ���D]��'F�⪩݀vC�e�%}Y���V��xm�G,"��m�/?�C'����0�-�)2^��R"̵z��Q�(�r�wc��C!���T}�!=�2�O���4�x5��`ǧ&X*XV1"�@�%�m,��ӽ�Z��aOu)׹�����FL��mjp��)�f�V��r����bu�� �
�R�!�Y���tW��(H����݇��Pt~ n�3��Y�Osc<�:zk���)4�O*1Mv���mO���Y�G<�5�`a5_r>c���T}򥈺�ڳ�>�E�Q�+#�pjM��w��(��U�Iԓ�߭���c� m�Q(uez���6%�k�0BQ��6��[y �0�ɹ��T��f�=��Ȱ��4e����dK���"�W�xΓ�hi���ï�+zn��ǡ5�<���tS�ųj�!�j�.QC�I~���Ĺi��)k���À'�J�k�eYb!�5��ңB���+F"�&��T�^�M��+Sݬ$]���,�~h$w��lJ��u��� �5�V-�݃0���H�Z����;�<$_���:*pU���Xo�z�a�����;q�Χ}�D�W���Ѹ��,y�M��J�"�wc:���j�8�{¹�F�m͈0���B�iTR�ZȌ[$���r##�����T�~��b+
��|*�Y�/	|�������~��.���SOD��M`��n�OC������SԜ0ʼgd,�6׿T�X`��0���)��S�߭"�� 7�{�\�����<zgw��.�����D��=�,$m��`!H���4.������P����j<�cȈ�ʏ����7�	D���-]�!�,�,�Q~(~Fg���+l�0�0o�Q
��+t��7 μ.��ծ� ��$2�W�:���g��"ՠ~��������^���V�p��n��3�wj����	@6�#���.3F�uS9�����Jyԑ=�culA�m�t>b�K�$�Vr[�ikԗ,����M\~��/�r��B�MOx�O�HfD.	�[	�`�G�r��d�20ڍB����d6=��2t'����W��@iw�<��\#�6w�gΟF�/�Fs�pR���\N18W�n,NkI��؀i:g���(߶���}�q���&!�s��!���+7d�,)�����#�$8oI<U�o�F
em��S�FAk�± �G�z��]����;Ή���
%���|u�S�M�{�_,�	�y��"���@�`�tw���ʍ�'T<������Ɣ����a���/o���2���j���19�R�<�BH>Z�rƱ��X�Q�[��/
��,mLy"laS��v���p�g���Xr5�
�3�0�𜇠4���4x6�����q��	:W�p�7���7�����}�@i"č����C�K&�G��U��	�6�F%�EGSaK��-tS��%����O/�^T8��2
�>���?�3���@�z��ʘ��H��eUJ+T�Ir��O�\k��*��P7�0`�u�O��44�L7i���q��t��Gs�N�������i���:��j�P��2��(r
	�����������h(���J�K�E?��/p��|����Kg�b*xE/`�D��m��g���x��U�~{p�W��i�V�w��VV���	tVV��L.#��#5�_D[��i�ƂΌ���� ��4o�*H���
����z��T���̻'#C7������OٚA�E��Z��j��[]L��7�&���G11�/+���AϿ2 �E姍XЕ�~d�O�y�k��O�U�;[� �P���Q�y|�#�g`���.A����F9k������"6������E&[~��CY]�'��C4X姌�$
��Y�����	�~@AZ�WUS���A9N��c�c�*� ���1� �p��i�%'I���Hrj՘)9� ה[�Ǌ�?�!P$ki�l�ګ
�1Ik5S����������+�jy螈g�r<��ya�`�Aը��Q�j��)�.�i��<g��W���q{n������V�[N(��{�L���]B_�=�s@�4P }lS�\`(Oo��f��J^�d��d�[kH�D�)t[��Z����\p� /4�1���x�"N��v��Y��!tf�=��<爉� ����urGU�oͥVa~��א������X�*������x�}�p���%���B������.�]�u �s���ׅi���N��1����1Q�e�� ���|[�2+��-�''~�JR��F
D�����)۲��4�1܏���%g/G-c	�(���0����r��ޏ�F�E��ì�.�&`r,O�n��?�Ys�A�i�es���a��&�m2!�[NA�֩GO0�͟��$6a�#�y�B��|:���M���bP��o�����P(��F;���"��������
�`���wO�wa[Jh�ًJ��̪#��F�/~�%�q�/�YN�)$����	g�V-T���;2E�v�	���{>0^x�Pcjk觡#��Y�����@/�m��VԜV��!�K��m�	 %q�q�|����B8��O䨵��԰�,�S�ZYd��w�=�˪����w�$����/��+�9�:y�}8kU���S�;d���_r�h�[q�~g(��gο/�h0[���E��3u#�4l�T������<�z-ꦜ�!�.�����ũi�LhZ�jU(���zvU�>�u�[�W����O2 �s��2�b@�aSF��f6�fF��s�z��2Ӎ �f�F��NA ����_v�O�.��0L�0?��W���s����	�w)R13닿 c�!Phv~U�I R����(��d
of'���1"���R�d��#7��
$�-d��bs\�b��K���o��_,���~�z����Vl� t����@΀?��)Z�:��<��J��Mv�R����#<��)�"�5��Iz�>�����T�� W��ƣYN�Q�"U��8e�0�?GM���b��Ě�aJ�dv�B��V0f�5���b�į`1RZ��?�-��
h�1�<[{�3�5W����.al���lbf�*�3	c����2�7#�qe���[󁶙t�n�+5���3_G�e��K�4���������*��۵Yj�ߘ��h������X^`���^�}'k�J��c���=�l[ު�3!�x���V�WdO��b&�BH$&
OHոKƮ�ǽ�U�P�CL��g�e�ȱ��PEN�ӱ�H7t"9}3V���e���@P�Me䚹��zq���X�(G5 _�,96ը9m���4k�r�tⲡ$e]��w�mC����P��l�A�2Q�1��A-��T�=��]� X����h���K���e:�-��問��l�8p|'��莧6F��%���4�"҅�����IV�������B���g��Wt':�I�:�$�Y��k$PPJ��������q�c�7��o��2P�x�'m�O
5�|�L��:,@|���41�<��{��b��	ﱆ�����vr�.	V�Q^��V_�N���I�rY��Lܙ4��_��F(�,�p���K����N��x�XyL�n�yH9ń��]�y}�ݨn��kP�6z;�>�U�	a�k��߾S�*�G����+�;��K�T@�D��r;����o�H�����Ⅷ�A��bR���[p���$�EFR��i\�U���c���`�_���B�������i&�Z.��~����=�һ��V�4��B�^��C? y�(!3� �=��Ī����R����Cf#} ��>]NL'�W5͸Y����t����P7�!C2Y�%|�t{�>���?w,'O%�4\��҅�||��x��z�&5ܰ1��mB#�/��L3�-��;X�r�0����o�x���KR��Qy��R~_G
���G�O�2��(�|��g�{����(pt0_F���XO�궗:�% �p���t����Dex��0RL*�
\r��*˦�I�A���pM����-�������8MD a7�����T��Pls��|��70�w�9L$�FD�?ވ�ʽJL>�Bn�; nN	��¡s����������#���A�Ϟ�`��;��tgi���»��B�^-�*s��p� {Y܅g���f���ֹ��8���� ������~��H��q��� ���>R8&��:0!x9$bo*�b?P4&�jza�4b���?�y�2�ʩ��=��1��Y�kfބ/�i����1)��$?� y�0dxv�-�;^G��rz�}�~�˃��|�nQ\NCG��oR��=�!�	�a�0��!c����3,L�04��+囏|X~�׃��w��ݤ���x�)��w�A�N[�&f�.grGd�dh�L�q@랈c$?fѧ
z�M����jz�&&w4�6mo2���{i8˝D^V��ǅ��Kο]�����g�[r���ܕ�M�N���$Uʢ42��}j^�/����ݚ�!
S:ϸ.Ϛ�r���~��A��A���bu��f�����p�n!#�)����$薗 �����İ�`�-/e|�ߨ��w8hyB�;�0��2���|��c"���]/$6Y��܆_��9@UfY%�Yh�p)YGd̨���*h
�b�T�?�S9s�,/>�ŮTD��� ��{�Z�ߐ�HEd��nv'�j���ԯUqy1�	�9F{�52�_�y�f�t�x�W�9��y����(Qk�!Gg�A�9)�!�a?c �=�K��4=\]x���+76���.+���v@2��Ͻ!��m�G�,(��瀶��\���v����u��M��kP�c���Q��ڽDy�+�{�k���B���ք���S��f�~�K�fM+��_�[�U�,����	���NB����E�l�Yc�+��1�߰2N��k|�� �ʔ��ņ�ѷ� �fT�|�u��ޠD�R�R���"��R�N�͵���`A�3�8Mq�؂�G�4�p�Q�N�sx-3o�%k��}�v���S<�����*��,p\��1|�� +�e�wM�H��O��u����O��,@�vJ2����h3��Q`N@��|��8�`^EZ.
�#_�\���M|�yD����L5y�j��MG^]������N��]�7���h������N..��"d�?�`:��Z�M.�LZ���Gk)�.Uk��_��o��񵁘&�PVh翄ñ����iT�9�lO�&y�ٯa����4�O�8�[}^�u0s�`�<�K�K�7�J�/��ņQyF��ofψǻ���kI�p;b�����C���=�8�6����J��T5
ʩ�ܡUt�����'#)�t��j
����h���-�ҟ;pJ��X8��&�| �Cí�2��M�	i"ȄGm��d����=M��H��v�n�t��y��$�ͩZ����d��	�a\�u"�u{zX�Oe��.W#���L! d����|�xil������.�'(|��s�=���P�����ǋ����`�O*�]�p�#��f�d���d�'"���6�]��~�>�@�_Q�{�r��H��ڽ:��z�a�����J^�εB	A����Ć��v���7(pt��|���l	ɍ�8f���9b�F���u����1�������GJ3�̬&��$7��H��#J.<C'񊭥�`�ܥ��9�%u ��֣��þiE��W�.�IO3̵>B5�<C�mzwG���o�?�,�9���&�n[��U��X�"��	d6�;�i��34W�).�>��wSJL`|�0o�n��qUaIWJ��nԽ��B�lC�&<=�oR~g_�	�ѧQfOiʌ����b*�r�99g՗�u+�#a�l��Wv �n�����L��"E}���PMROd9��3��N�x3
r`V}_��hW��I�h�H#?Ѱ7mA��f�e�)ncģ�X�-l�R��Y��#�${�a=�A�4�:+�Hw��ڦ��:}iy��?�7:D���5}!��]�x�e��h�<�sLuv���׆Pt�@��(,��9䷂~;�v>kH�X	'�#\�������;MZ@�����bSe����4+S�޿�ɼ%�pec���5g{��6E!��V�pps�7��;ͤ�u$���^>�(�9���T�������%�t��&�/@+SӖ�{��C��~����ɜg�=Ӟ�7b��q���I
�a�e�^�̖i1��~<v���RY׆�Pi���(3��7I��q�eDH�~��.�tD�h�L�B�M�բ�#ͺ"��������<V�\]�"`:�
P�B+Lo��lHӲ;YEG>�c���/G7ݏt��h-P���g���ݫ�݄�X����3aIz�u'l��m!�bQ`߅fh0�ƹ�LNt��5ɗݳ�w�����H�q��\�۲lk�������x�d�];�w�w��x�̰e��
�\@,�#ā�q�,+�S@�h!M$Մn^�c?\�����D�9��G����:\������G�SJAC�d	4�DHtؘp����w�F�=�N�h�t]��@�ݨ�bzP��c'4�8>�R��W#�BMϦVC]�ڋ]D"r���
�B|z�,g���fX9����2HRz��o ����a�'='u�t�X��A�㨾��(&{�[��5*��m�#{	�ުmUm�y��{��!*����~�q�)i�g*�O�G�O�/W��l����$W�e:���T/+Q���/o{|���]cAMR�z��mKa�f�3�{�Ko�Au�c��0p&��!4[0��"1���� #��M0��e���"�G�Td.���	N����ÈKgq�uy��H�hpK�ߵ.��3;r�?��(�s�:��b����kG���l��WJ��Mg����t�n8�ZKs0C[���!Y�pPü6ĔK/v����P����X����a�Z�����ap�R���R���г��O���u��r;��R���� �_:�=�j�M�2gȻD��j��},���6�>�s�K^c ���1���eQ������B���눪��7|iOC��g�ZU�[�ڗ�W�K�6����R��2�zd��TM�ZP�$!�V���������6 �ױ��K�2>��.y8��,��-!�"Z^ɾ kZ�@��3�L�<<9^��I���W7�Ӫ���/���9�t���WySi��:p�>$�T0��*j+5��a��fJha7�k�������Kb5�� �^z7H)�h1N�&/�u�ۚ���2�����}�.Ѵj�~��7���~�y��b���X�%XI��}z<�\&�k�LC��,������d� ?�5X���4ۜڦ|E�b��n���EI���.��-a�ڈ������ؾBX��X�s��i�s7��4C3:�xI��,pca�����;���Ƶ9�����5�6wK-��;�M�:6i�R�O�������A�K:�l�D[��E��BL�{�����qD[��=l̶����m���T�U�=7ˣ��j\\-�뻪��2�5;�|��@�N����|�E�A4EW(�$�g�~���B���SI�KE�^���u��`�3vO�DhI ����46g
hy2�b�$�A��Z0��s�ĕ�{�BR�8��8�^�-�Z�Ht��2!��EKy��	pq�O�X鬔A��EK���(m���<��N��70��iM� ��9�#4��o�<��%GQ
���+l&�����]@��q��|Ìv���10�q&��$U��j����h��!;;�g9�y{�@k��tӆt�kM@`��j����(o�s���0�����f������Ḻ�����?]�c�"�(Bqk5�s&�]�[��>�ߵ�:�f����N�q�!.x�h3E��(����G�$L�K��R�#h�Y������:�C$�s��J�Ca�#���S4	�k�f�*�z@��
�_����\݇�8��逷*���%�f$�;��e�$�S�+5����U
���p��M��g�zs�����f����V�uV�/?��E�b�2������n%�+"��9�L�w{79�kԙH�ӓ횧|bB��`�����H�^�U۠�I����
q$4�2R;G�jɳ;R�|�6����׺e��� $�x�]��~6�h6�纷+�c�ꗄ
U<Xm�R����}�]��ꩢ������,\�h~l�E��~������)J�p;s����T_�+pu��.�<.�!t#��cK�S�l�5*�!'�EI�F�G@f��[�����o�I�H�.���Q���;q^��''�B�T�'�.h�.Mp�®��ܜ���}�v�eF�3�:���%U5*®���������#Urj������]ܽ�~���'�Ѱ��iׇ�;���'���`��V�ז]~��ׅZ�L�#���,lZ7
�kb�=!-3��(</�E�RM�Z�h�(t� �X5�X;-��]h��AJ'r;}Z�gq����DX�Ba��O�X?�	�ۛ�Q��I� 2ʌ��y�{_qu[�>7m��[������Cn�3��]f��
�N�|�?��bJ�g��]_ZG�g ��&'<���/Nbʸ��v:1�R���1�YT�j�;�P�B�-F�ae��j1�2��5��B���;�S`�r�?�*>��߫�� ~��I�bT���^Bh1��Ѫl�1�uo�[+;]����а���gZ�ራ!\��n��=��x��_��4����ܟ��:X8íJ:�J�Yn����:ڕ%b��4�y�s�����4ǶJ����rV4��^5Et�k���_�R�ZB�cU;���78���(�&Y�LAD��6Zo�=�	�mj�I"��Cfh��P^��W�:>��CY���'�y,�����_�3�М��Wr@KH�.�����.�"�Q�?��
ĺ�m�͐d>"�� ��w�l`2�τerS�F#������SK�,�HauB���эt�0�8�B�8:dZ'D�-� �Bf4.�U���xl�C�����7�>���`��Il:��Q���}��
Ԟ����Ve�L
�^7@�~�a����ږ� w��dZ�� ����\��`����i�	�Wt;3Rd��.t�D����N0wK	��N�Mx�7�Y��� ��;V�Q��]��u��i/6:@=�.q����*j񁣞d$%Ïf���L�ENP�}5H� q<�u2�פ���7��9{;3�0ײ�C$�I��4�le�"���(�_�q��֊F��e*}r������DF�6���l��q��`��q���X����1�YR���mf�=��U���]Xjۼ�s\��N��X�G��YU��<���۴��h��{�fq!#lA!�O�����p�(.�l���ƚG��GZl��M�~qW~g�b�e�v����y�2�'H�
�=�C����T}M��7F>n	�������g�2�� �g�t2�b��<zγ���d/^������E����d]e\,�y�pƉ�Վw�+^�H@��0�#��2�f0�����#�8��%'�iP���^�Y8�AӀ9$�nK��3C�[�>7�Ԥ:�����`�&�čޢ2]c� ~㧐M��Ĥ,)�����G�tIW����/ǣ�&A�o'}�ױTQAW��O��ma7P�Sf�V�3�q�6̀`9[���V�G�v�@o��Ӭ��Dխ��"'�4�@ř�<���?�m\D�Bj�Q�}�o���)�6/��kb�\#��j=#��V+��P�K}:�(�j�[c�6�F"�*����"b�w&-�"#cDG��T���K�����=٦�%�P'T"�Gρ(�O�J�CpV�N���ş�Y/�[w���E^~4�:�@wW���O�v@F[�ZQ�����n���[ּIm4�|��z$�����`�$!s8�݊����\T��,�Uz�8���N`�_C-X/ʖAb�DM!�>�@���
�s���޾��;��7����9~�Ձ=�������q�Q'Y�>�ۄB�8�x����B�"o��OD�W��6K�J,#A/ ���È�#�9*��
X��� 8-5@ :��^b�!�w�V��h1C�Z����M�]B��3�͟Ke~�/�-��Ѵ���i���/g__���*g;zgQb���E�Tq�]��v�m*��?���|����ŋ�2��T�C�
9�X�C�����\��wrs����aS-����K�!Q�w����.ضq�Bp����p t�7DPfGY���*�^�{� ��"�U�v����f�,,��.��g��L���1�3aAk�7��7���{<� \�����![aZzk���"���K�*��n�f�[�ӟ�<�3��QY��0X"G�(/��+C���L�
����7�fm�k{��z�G�+�s -��9:ϥ�i6���[�]E*D�v*'��~NS�f��<=�ˤ]\��i�󑞡��Ix.��C����M5�JV{�i�{m[����xne,#�p�v��P'*B!%�A\w�e�9<V<\6�^?

#��gZ���2�{�;*)� OA9
f�G1�c:3�N��`���;E�e%Z����u0L�!��Ňr͟W�%�{��C�U&� (��7�������AB���1�v����B���5]LeP�k����$)7ɩ��Z9�;K��y3Q���Cp<�+�[4���c�za~�D3� �y�\�W�� ��C�";$���3-ޚ9O���˿��K�'���=���%��Xx�<+�m̓�nנ��q��a,N��Dxp�,ZhV�G�`W��[ʢ�֊����Y ���^�2U���8<�R��C�2ƪ�a�k�����2��QI#���2	���<��
֮��Ѥ;^�|��X�@U�Iw�k���lr��@1^7A��H�~+?�g��c�Y��	Z��U^�;Y�$Ưx�1t�
{�ԙ�^Rg��Ϊ��#��9�'$�!�~\�`AH����ƵmZ�E0�"S"4,V�T��F�ʵEaH���ܞ�p�'��'�6��&���<�	4���m�-`��6Me�e� ��5�P��D�Y�Q�y���}+�����[4N�?:�ӏ*5���fY:	=��iy��Q��ԡ�a��ޅG��-: 5�� �������w}	�S���T`!^e���P��U�Y9[��*��O�o3���\.��� nvQ�HF�HB����
��۱�8S�͸<�U����$ 9��|��%�P�iO�Ԙ��J��PnI���L�Bb@���Ef.�
����u_<^��@R����2`"0v��"�8��^��?�L��V�ߞHe�wVH�Z��Ծ�73�D�< ]}�˓�W�[%�COTn���^��a��ފ��Cϓ�k�Wg�Z��,-���V�Az����/��̯Ol�$�D�~�5u:��
C\�q��+Ψ7C���O�|��=�$w'>���6��7�v+Q��ޏ�_^�u��G�Sާc�)�����U�ݞ����Jϵ`��6՚E>�܆7�h��<��{Zc���U=��tz�)�G	b&I��.�4
�EIf�{4:npY�r��8�������};�߻HA�nտ��N��t�7�*U﹃;������Nŵ9|�4��/�[m�3b��B�\�w�t4'Q{N�ϲ��8��-��ܖ2�2@��ꣀjA�Y�Ys��8!e�uK`)��.�?��!�
k���r�1_�ف��uȶ{c�x��=���R�D�n�l�̧Q���64��1�� �K�^����s�.�D�]"�Iy˚vԬ�����`dl� �ӝ�*+7���wK��7�]���}����e��e�u��9"H�=�	f���ȹ�R�6%<~ۓ�2�G�fw������e5����%�'�.�����P��N��W#(��/���Va=�@��0Ͳ5�JU��XEt5Ç�;: �>"j���^=��G;�M��UX�?���
$:LB+��'6T��7��
 ����oh*�s��H�N������X�w��9!;��G*�є;}1X��|��
��T�Ծb?x15��b"-���1�B����W"���>�i�h�o�&Rښڞ��t���֠I
W��S�fY��83+'�RR�ن���PC}��dG����"��^;]��شJ��bD�������,.m&��S���G��]��3 >RV���N��)�)�n�X#��� ar��jb��!�_9�ˋT0��)�H̬��r^Ԁ?�qx��?hF���^#���!���W���J�??V��xT�>V������1����mw_cn;b�tЄ[�53�Y��\!�)ֵ��\�Di��Q5����^(
}v�>��u󚔷>+����Yʄ�^��J�
$Zi�:����мjS�\����ebJD��e�+x�e	.��B��c���4#�r�Lޭ����ٖ-�Euc]�2T5\۹��CE�n�� �V]����t�S~�ֆ��A�}y���w[\�$�9�����zn!�X��N�Zu��)+l1��8�֛��4�]�Rv����a>���P�(`k�B���CV��qd얷����L{�,���~U� ���?J�����#edbc[-U���cw@�P�4�O��u���ǈ����*���q1�O�u�0�7�#�{`!�P����G�n��Ew~0��Yt�3��-Y�2�Y9������a�����_INx�E�UA�ܖ��Q��:-�JTC����*6E����!t�|RU:1I�䭟������hӮ8�N�7\�S+�#]و�6��d���=�zx&c�d	L�9�偂�yG����>�t\�����"�����\n� g�-L9�K �7Sc���?��ѧ$��#q�mL����as���%����8H\��	�e��P��<���<~ǀsd�ڼ����3�-��y�t���5�2x����z��2������j��b"�����DсY��8�|�i/��x��X @��V��{;z7�?���)�5;^/l ����L�U�/Qu)�g\�),�j��a���;��v�>-�օ�qRp�A:K��қs�.GVG�����sC��rZ4�8բ���܊�Ժ);%�3� 
m�燆V����2�Z�I�pE����D8��}�}�:�R���3�1���A[d.���J��473�A�Xa׮�Y!~iF�j�P��q���r�o5��������>�nШ�8P��G%j
�P���R_1�ִ����	m��Z����n3��(���]J�ĦB��2��'���,���C�!�{
beM���(�2�JM�~�2��)��9���b���#�(1ִYÐL���LT���K7�Ch#e7^�AZ�t��iWb��Ň���H�
36˴��C�>���hv6U��������xiyo�c9= MR�zΔv�'H�G��!�J���&���W,ND��+�H���2c�_%�Z�Q�ݧ�.�^��đU7b�[M���k��W940u����[��-yU�8:4��Je !�f��9�8y�	8d����O
�ΏC
�E�)�zcRɸC��7���Sq)ΖьT�nYw(C�l��]����[J�N�z)N8���#o�+�� '�4//VT%���9�� ����V�8���rZ־���B.��x�w3e��v����Ʉ������2I��o;��*����u@�xK�^W@1̨w�4t�uδ:wF�.�y%ԃ{u�����-���>��R�-^*�����_�x<i�8�B
R%��Nx�d�Ud���P!�Wһ�\��Ss�)n�Z��g�ֶ"�G��F�膺0<̫����y���"һo3P�H���3���mn���k��b��I1쀛y�{-s"T%��UάS���'��d)�/� ύp��1���/�JS�����d�ɰ�R��f�'�R
��6����J�>�>=|\�S�Q��IꡞHM7�S��v|[C������:�PG��>��u�s��\�u�-�ށ	�J��T���:`ly[�frY��YҚi��
�[e@�7x�4+rf��Y� ���M���@t����5�/XtN��J�:~Q���%�,ܧ�^����`�SP�~���������"��P@�����QX��y�mޔ�s]m��i$ݠcK�O^��rc��[`۠=��)O�#��%4��������{3�H��״�j�X(3����F�Ws�T�����er������KDf�{����<Q94u�@%A��b"�wք��N/�jg��M���{6�v��l	m���AF�N�R���w���]�oe��m$�짬C\�t�Zx@�G)�����I�>���VQ��<�?=e��j�%�u���
g<���RMsD�xأ��]IOWX���L~;����ЮNgت�����\��?�#�k�m��ډW��F��֠��0
>�$rr	����2 �<����-��E��0B<Aل㖛�.C�0�a�r~�x�Z�c����j���a��JA�S�q Y!N?Zŵ�^G@�����v�3�����_�~��̋�PE~<+�kT�����6��aY��+��p^L�T�,��~�{:�'i�J�2,�m����bV�ބ4@2�)����b=���Nr��>�Fz��@�o'�n}��wV{IH�&�)jNmk=���"�ϝ}���2��'Cv1�;_���R��������{�D.����s��]hWf	����q�2�
�y��N&�����L���#��I�A���q��ѾV\� 7�3as��*��x�4M#P�>��,{Q}&p���4�:�l���	������]=/Ъ�_0X�}��%�'G��c�4i,��q�U�p�@bc�E���b��c�~����A(0���s�>��S��i)�)�L��)��\���K)��u���g�|�"���f���cǆ�x�`�~����eWW�߉�d��^{S�Ҩg_����H���Btk}����B�C�?��`�������, �T)��������M����'�˜V|�$.��0��t��lW�K�����D�HS�?[�S�B6bK���u3^W��N8�C@��%����|~/f�Eû��$����Sy_�/=P �¸����KH��
�l���4oH��f@hwv�ok�g�Μu�J�o��
�\'�Ud���h6|�z�%	ߒc�Ճea^W�C|2�.�8�G�+2��i� ����5��C��D�)�� A�,�$e\Y�*��  �N�&��"�Eze�iQ ��b��R��O�n]_G˽���)>�!������%�H􃒄������G�B�*Q19��N�?��@�ՖF+��0=͚�
����R[ B���,i���ds���`�#T��yz\�Z,���[ޓ�\;��ٍG���Ժ�'�n��n�L1�5UDT�so�ڭ�K��S��%yjIrݶ�o�~ó�,��?�vi��6-)�*p���-U�����݄Jː-�q�R K�@쌥�Ȩ����o�� .�_I��HZ�9��g����U.��=	�j�[(�G3��qI*���}$w����� a\�vr����n�/�9�閃)��vHy�V� �-$����p[�n&xۄe�@H�Ї��;A�6EG|�WM!"�*��[����X5i
_�y�l��f"eM�!�n�����ܦ(�"���CTn��vVN���S|�!+3��Cٔ?�[V�����U��:�Ia��J��s�>0�����@?�Q.� CSX��q�[W�2Tv�q6M���^��}�dN_<Z���@-ʢΠ�2����̠�Z�t�˴`����5�Ue��ҝ瑏���T���*RΖ�[H�v���e�[�h��]���LS��	S��u(�<��̭E���`K�M��08bR�Ķ�:4��6(���ỏm�aҲ[�˟�����H&m�ǩ&%S���٩��j�l���½�7_�΃B8OL�`�z\S�U����S,.���D3�{��wY��&F&��
�.�D�ϼ����/�=u�񏢸��a�q����h��e��i�LC��^ru���&�?W3M��V��)p�)7ݲ�uig�$p-�[��e�+��H��8o8R0mo�z�T,�z3}�#�?��r}p���_��,�k��=�V�y٥�A�x"J�M�z�u ۍ�	p�����*�pcHf�r�W��6^�P7����Tޘ�j߬ݗ��rj�Ԃ{��Nzj���{Е<�S���_���U���r\rSG�/��X^��U�~�'O�3gP�٫(c�"�q�Tu��`����"OOWZ���������X�J 0bؘ�/m�����s��-S���y�׋���Pe��{�]q���p���$Xd!�h�+��L�k*�Հ1A�:��@2j�د�b�z�=�'	XV\pf,���`V�[��t��j����p2W_,F��yW��^(D��N$�� ��]�ܰ�~������茯���H� i72 �R��Ζ��	0���Z��2�M��K(�P^¿Bٯ��	Q��gYcs�
�]�$,��5��P�!�$%���kxじ�d�0>��J ��c8ͤn�.�Yq2��v�0����9�lb+�*��c]u���x_?�p�TQ�!�@�h]�|�v�M��wR�W�h��&i��&Y8:��-�fr��8�bz�2����3���0����j��u����CC{���0�Q�#�h0�աJ�,�T��\��,s�&�G����Q���`�@̭�q��)<T�rJ�L�m�;�ݜJt>��V���7� �r�iq\
sd_H<6�l���¼��޵NJ�}G;6yX�\Ln���US5�^�s<}�Sї\�P������K�AX%`5���~%yʺ5�f�
�Ώj�Fo����rFOEj2���f�a���.�9�	�	BE{�8+H��!T�rTo�E{��d�]֊Jo��W��(}~[�##�=�5m�@_���xn秅�V7���?�/���i��[Mv3X��:"��T������N�k�T��g	p�R��b�k�=��-�3�=6�ˤ��rY��~�����d����
D)Ui"WL^���|�#��'E\��=��b��)	�P#c�'���Ŝ��%��vk/]0y�Ū����`T �KLz��d=��a�8F�j� �B9���� ��$�7�%��ؿ7��?x��E�Gk2@ʆ�� ��V���ܶi.PP�, �$-ұ�������oW����H# ��ЧMT���{Q��7?��`ɩ������R-P�bÏ��aH���|��~�Rݼ�cD�FejM�eD�K�eC�b��$��Ђex��p�mGm�'7^�w�B{��ΰ��PU��r�n��ܻ��T"&?�T�����%�_��>���Q�N�F.�?_+b����1�J���qcD��X��h@R��f82���&&;c d��̀E[�a�kF� ��:~��Zם�BOW'H�w���,\!�����؍�5�b�_4�8�n�}��I��^�@���!u0��RPD��_���ⴆ1R�J���d��P���",@��R���[��࣓�x&5��_�pɼe�U��<:-��=�!}�$t~2�������p�v6!���p�VXn'%k��Ce(��Fe��a�q-iGh�M;�3�<=^��p���� �O#F|lb�3Ɯsj�!������sL�b��?���X-�I̐H;��}Ne1i�z�<��D#��mo��2�D�A*�~򣥷�f;�<x��ނ�����-���Ci��9���c$Q�m�~o����"5���f,�r� ?����V�fhT���˨>����S�J �xV�܌N��&��h{�'x�P?m��[�gσ��X@��9��[J���Dm���s��B�3*A���R�e@����wIt�nWE+P��n>��1�lp�]�;NafmЋ���%��%C������'W�.�3~�P�3��`sO��iK����#ȲC/�GJF��T{!�Q�HcJ�x�I\x)�gn��3�ו�vɝʕ0 �FUtB:�0݌����Xqw���#ޓ���-�zg���FމQM�~�㠣�q���a���E╚��B�wB��
ˬ�n����S�������ɫ������2܎�n�]L��#�#�.6)�PB�Zu�'�q�᣿��DSP/�Fh�E�ζ�ʢZ��I��ӆ�p)�n?�t\��x.�*���p��zA$ϧ0(%����N���h��?����Q��s�p�=(�.�fZ�s��C&�g	�N%��<km�V7����.�[w�A�[���N<�z=D^�"!i!U�}�(O4v1ِ��G�z�l�^Ơ�x�[����ytbq
*�.�yI�t�f?q��ڣ�W[��<�,Q)fP�3�H�E�޻���ƌƁ��^_̈́��D��ﳣ]Uu�[�`(�� 1K˙ݩda�]N��쯊{��]���q��h���ʁ�Z��q�py䇜��d������r'T2N�K|�ѺS�2�v=�1��"ۿ<!<.�77���[jל�I3B�=�����)&�7'Y�!�㻹jt:ż�麑zv����#�<n;D5:���yu�(�YX�D�e�����y�y�����l���R6�1�b����Y�հ��F�������\R����=;���[u����9�BW�P��y�y�٬�N|�|�ok�Fa���Zr��G���W?-��5�$���𵣙a2(j@���}~~��u_��]�ڧڀ���g�B�w\���f�*0Z�h ����D?��|�b����~��{�Ait��f_�p|f8 ��B؛E-ǵL�96Hm�P���vL}���5�,Pc#��cW͜�ln��b�}���W�0j�.@�V<�D��:��'N��6,����Rީ�@ʮ����SC��`�C����g��U*�B�B�\ ;�>�����D]��|�-�=��~lv�mD=��Hh�2�����Hi=�Bԡf� 7����q@<I�(h�ާ1��r-�h�ϯͮ
BWuU'j�}����[hU 7α`��;u��!�g��J-2s����V`�R���F�}b��	mlV�<׋z�����&��_��1L��6�GӁvO,l�S`VÜ`�}�]����1FF�㖘pu���n<��_.Aa�P���u����s�����a�*��j��%�Y��"��oBp�,B��cv��a����i/7�ϒ,B�Zx:���-��C����j��( T�T�C6�F}Ͱ�o	�gl��dAT��H�csK&S����cR;�Uٕ��.�oL�o�Y�޽�BF�!x7 m���t�r;<��v�غRhX��I#�
�w%X&ȣǶ]IYtٻ۱�ݔ;a֞�:�%�Ì��.�u��
�ل�or`�m�D[H�5�u��w���v�(^Vi
tZ��́�<�[�n/F'{v�P4l��d�4�G>�i��۝��O�&OH!��BY��2b3@5����6���w�i�l<�&���lG���O/4V����=؆#�. �(ki�o�Ry��,�ү.��`7%���cѬ�zJ_���(�NL%�ausq酰%4�y*jp��S?oN� �����Q˖3���b��o>xm)���YZ�3�œ���|��|~IB���mV��5����;r�Y��Q��a&��_;{��T��n	�Z��MVdp9�H�R�����9������pt��:`}�c5G\\Z�tl���UB��Q��JM����8M=Gtħ�;��EYe����ScA��dZO''1���eaM<j�%H~���/-Z쨝�!�S��m�n_��	�:^;��*�yr(Y��C�XϞ��H���W�tx3=X��s�a��;>u��h����¼̐b?	H٦�A��!��i�|Q�'�G4
���FI�������מ��YR"f��߃�7t���l��� ��D�M�OD~=��o�K�\���;ǌ�Q���u�I��H.�?!�`|����>k-Q��F�K#N>*�o�v������Z��*��
ʤ���e�*+7���}����e]�G�0W ��W�!��.4P`шc!(���s�l�X����+8y���k��4c�/�{�s����O�����Z�)�d�c��s�ڳ��_��5S$�DUn�2-���/	� �!!��/�%�>����߄�7X��mX��d��L����Z�7z��CH~�K�"hR���8"�N'�7p0�k�������K�+"�nx�2�8�� ��b&�"e�ů���6���DS\��f�|�w�Ӯ䷯[����f��\Q⁪�b<����PP�	��x�}�|9J���5�H�����c�KX~��!Ā�}@1�R����ڦ�U� �#g���8��k�@��j
j���Ө��Ϟ
\�'X��!�����\N	I�j�A{{ޕPk�8�JL'�2
Pt�-�;.�gN7���~{:�En��ă��˞��z l�R�t?M�I�-�χW#��MN%bM>D�� ͻ>9���iX����1�2_O���� ��(&� ����_N�!��y�`�1/?'�F_q����#�R�Cp��Ձa�'�� j�rI���^V��I����o��p�"�ׁ�������JoD�0G����h5�iIGܭ ,NI~�OU���:9Ug�u9^���Po��W��VQ�!�<��g�V�K�KnM�ȿ٠�����Dբ�3���J�9e�5�4w�,�?��­ZZR��H0��K�)�$�����}Z��f�r�-�!��JȪh�]e�jd�����H$GC��@$�dݲ'�-�,��!�׼)��&RĻ��I�tm�D�]�@h(��.&ak��n=����ߞ����sˀ���e>u'��I��EޱB������Q�=�s� n�s�S�5\=�JSz�_1�&j}b/V`0*$���]6�<j����Q4���\ԆA���o����q�*P�*(��a������	_GHB<X{r��$�t%�V\�e��Md�jx�L��T1��pHl%V_�G0˼�G13�X��"z��/�i6��֯��0�
{�wJ%��]��1�S-��R=��Z[�/�W^�r]�$#Z�gu`5DI'K�p��ϲ)b~M�'��B@p�~���O(�v_���H](��t����a5��}�%��41�,���1�jy8\�;�$\����5���3���Qo�b����vG�VC��K����[�����n��"$6���يlN�'�����=��\?����l/d*��$�^�?L����R��J�q��@[�F�����ɝ����`!�V[mR(�p�1�nP��/z5(�:N+x�&�iw,��V.¢Bh>�������_�_8G
a|�/�ޝ8[C��i�e�=���Y�ǽ�,f���? Y���K�>��ʺ�|�F�>���mѐ��w��!Y�)|�!���RZЏ6�X��'���'3E��ŏ.ͪ!+�a�֋�C��vg<�[��qWy׎5�b�%��7�`Y#��gX���L�Ȩ�	�*��U�`�:?g��8`Dm��]3^���&ױhzj��ȭ�/�ue)x�$)ZA���S�����U@�%3�H8`�%U�RL�1�҃��7qh�M�gh�+BU�8ϴE�ſq17I��P�+3���ab�"��X35Km2�mI&���-Ac+ξavຶD�����X��  :l~�	Ti )����������3M=�i�E/����:�� l��z�
X�%�%Y�w+=�r�6��QB(K���7Ȩ�3q*W�SM`����ԭ��u�E�ɞfc���� ����H��-��|��:�A��;��Fpv��Q힟�F�p�>+e�0S1S�x��,�+N�G�/|I��~Ro�S^A������q�S	��
�5C���1��z�Q ㇢�(gR���2=v�Մ��4і��b��X�F���¬�G^�0Y��2�p�~	���B�_>����pr�*���2<ы�m^�g>�˅�mb�*+9�P8	Cu�K��'� ���x�0ќ>4Q�4�HA �ݤ�ymV��u#�h��C�WLl�/�;�S�� �0��_�ɍs�@�F�GXd��������!ic+�S� �	տ>��Ǳ��T���N������Z����"�5��Ę���F�*О�k��S6X*Q?ˊ g�;�bb����,�����9�7�.;��<~�;^�u���&��d���5�p�K��4��(&�@$plqV�|�8>�/k������0��M�^���F^7is�:�"�A���Osi��Q'U	�m�:��x��/c��>y�DnT��q3�i�7d���J�?�� D��L�.��(q�-�J�|�wID�_[�g#�
���a�^1�6׾o�Θՠ���t�-��Ė9��s�@�D��o]�f{���6`�A���9H����I!�taI�ɞ[��O>'�d�-��e��!<Z�g������9�t�����th��l>���P�kzE�k��
,�_W��E����� �b��J�x�ף���ba��Ac	��$�l�hT���8v寗z�[>M�{<�V���]%d!9��@���7W��2˒�z	`��6���Z}YX��q�61T20�\����u~p*���z�hp�Ov�OЩaF_���^x�gB8C��ܼӃX��>y 2_�AC���(�y��|=	�3��Ǜ�� K��M�h�r�
B�k3X�l�i��R�[�њ2�>N$xd`�Z~'4������l��:�#mC�~�M�&��@}��x�.z����=�c�c+KGR�oS������JO����ZT#	+</�2AyNz�Ћ��Dým	*�{���H�΂h ����2���x�%]ɷ��4���cn� c<n1���%���5��|C��9�i\Y��'����)58���9ca���)%����<��.L�o#{g���z������ⵐ f��O�u ˃Y�~�T�G��HY0⪟@.���jw�Va�ۤbw���d���s�89���E�2]\
��sw��~b�ĀU9{9EB.;Ҽ�-�&�nY�~��`ğ9�c�SDM;E�R��CC��+��?�&�f��ŷo̥\�� t�ؒ��H����m7���I��&��b�wt�����Q�I��="�8�j��ӿ��H�  ¿� b
z��t3p��乍9y�E�[�wm�������o��т���|�%N�v[�p=�9��5[��H�#Ү92gq�؄/�0���eu�9�B��L^*�P�A܉�-L�P�q�:���`n؆ϼ�%)���RM���n������lS;�T*#��8͞�HzN-��8â���ss�����dW@��ϕ���ko@Q9Bs�P����m��ߋ��^� =x��O����^�52q�p�
�r��|�:�s-�g����&�
�NAz)F�b>k���:.��ɓ*��f�)�3+�&j*�FĂ�<��ߞ�%����G�[��gՎ"�"��ʠI�S8����D�-�	RO���Ӗ?����x��s�ğY�Ӭ.�_jGT�؜j��	�q&y���:�ͨ�/y��H�������/}Ts�e�Kd���S^�xtWH���F�՝z�a���s�Ly�0\����X=*1Qc�,h�]s~���?��i�����"b�������K���#: :*�^�Xǜ���z�%�����=G{���9iQ��ЃR�QEh���)w��q������~�@Ä*���-���^�)���g��2�������V�6�� ��7��h�_��WI+6I����H�-륡�PS��+E+��j��i^j٭!��vx.��������MS9��˒-`�ƫ�L���6͞��lSgA��y�Z�*!�k��ѐ���L�p;��UG2?�(��Z�ÜX�v��cʻ�;0���!Nt� ���i�
�0���-O_%ıd�a*��
�N�6�R2e5��~���b�<s�R̔�+p��@È'�����_)/"�;���Ba��=(�\������4>���P[�-�������S�G�RS���v+|��j��軮��_�j���ꂗ�R��U�UT�r�'��Q�L'{8S��Z_����1�*F7h'D��8�2��,��Pw�.��_IՆ�o�_pא\覿'Lߤ��;�ﴶ��H	��ʏ�6���X2:2��4���u2^�E��f�B����.�u|ѸEv�+]��<�_�5����Fמ���e�`�����J�f%�"_Ÿ��.�	���*�����Ͼ�P|���ׅ�����7����E��n©�Uv2���b�Q^�ZB�WZ�n~�����P�.F�9I�SK���O=������~Γ��y�Ԉj�b��35������h���>CQ+�=% 25��3~����x"�AQ�C�Ϳ��R�	��j1 �F:3�k(SG	TR���n�p_��ض����?xS�OC�9��؆����f-7�w+�4�b<��\��(ɻ�� �M���-~����q��z�5p	;Yyc(A�X������'yO@n������u~u��Ŕ�R����uhx��\�)�NG�x:t����7wsܜ��@3��b���m�I	{�q�e�-9�o��G7��
_�)!��=�ЈĔ���<g��@�c���qH�մ�슺E���=�L��z��oT����"��2r	�W����W���]6�� QNT��F��BI
uM���2]�A6��Q�elY��z��S�����͈��D�2�!��g�+<�|0H�wm�j�ϋ�Ӳ�����e�,pl�?���		���
q#���3o,=�Q���w�E��D�y&��K�)#w�Xc()U��i��Yf@O9A�N��u�Eպ>�S�@�l�<�=���b$��Y�꾔�'�l��obzK%y������{/�W�n�h<�*w2q��j2w0��]��:���#⑂�S�����0Tۋ }���c�H$A
5�ڐ~Hq�=h�-��ѶG)�[�6��@�iH��ʶ�QK[I���l!��Bu����������OL�BY�@�D?�L���HbvK��d�"1<��r����pg�[*��u���W�R��=?EB�����aS�����Dh��X�k�rK��܀�GoI`��[��~��c�;pk�G�$��P M��m�NHT�fԎ:�O��!\�ħ���ݰtueS�Ht�3~TQ<��W�x���,jOJhй��OB��
o��� e:J���j7�*c4K'��޻�a&��23�+�mZ�l��z�k�pw��ǦέZ�Z��T�%���<���������?u���\"DL���k.�GJ���u⮝��������6g�.�+m���7�J|]����
��p�LǶ�0d�E�vr�f�|-��[m��јBj3�z�6d� qtQ�*0 ״���b}��Xݵ�����C0���Q���C$��{�c}�t?�3M�|�L��D8?�yS�Oӡ[۰;������A$���R����V阁x`lr|��<��6���,�J�R�'�c`,D1��?Ż��¥���z�~G�ʛO���� ��s�9�z�T�n97~S!&�����D�~ �+צ'��:)	���(/����v�@��8ڏO��}Q��Q�����j{�(3�<�v�ߧ dl�u�w���j���x��9S��j
=�n��r{�θ)�פ���Q&�#��<���6��,ƻ1u�(S���j��6��*�@q?֧���q��6����!�_p���V�nz�\ e.���w����3]����8a� C�x)a�|L:\�2[���I`@R�sS#n�ΐ�9?څ��b9��_�;�&�H�ϠW�3�D�tL�3QF��#BG��3쒬�6�l|6'\ep7�����Ήg򯵍��+v����1*��%G6��M��?�|�0���"��[ۺ���ʟ������I�{Y���?g5�� S���چ����齕��[�tI�4�_/^#6��A]v������Ȍ�;��O��n��x+��v2�V)�N����b�X�]��� J,�m��`��'�C��wXDk�D,�d���?�g7zT��@Z_;0J�:FA�}�(�-p�(�ss�������D>~ϒ0�L�
�;1�TS��-<E3R��@�b0�}(���9"����4�s�Dt�U���k�V�*�a��l�S߲�����8�@!�UCͶ1�uc_�[����]�������u޼�>7Y�U��x��Re���Cb��ܤ�oDx���qFT*���V`��0���k5[2K�^k�QSrkQZTG�����<���S�Y-;��~�Qi��B�\S��!1�l�{+*�����������vW��PH���5	ᕇG�B5b+H����׋@����n�  7���A��I^�A��z��M���xӦo����(g3��9v�B���%-�	��3%=�f���ǌ��Ȩ,`���Ҙx��8������i4���l�W!�H)������\�v��j����0�!8BX��n���|y��k��mB"r�wȜ��8ɹ)bY�����������8A��j�gC��\L��)�@��o�ӌ�B�ނ!8@�I�(��N�~��t?�� e+�<���.���[���
4��ǂN;��H�ݖ�b-���' w
Ry]l��i�2}����JT��U%�	����*�]e��4��na�N�< Kt��0���e�.�M��I�Ĳ�ʙ��A+��§*��@:�@fv���"ꂍ1.�����w��M�U))D�ɂ]�w�2����PA�K��j�?� ���~o��]b�Es����:.GʟG^��w����v����������M�Q3��٨ 6::��f�	�'�,���M<t�R_��n0N
O0�(uG��=��#O�ynڏ�f�A�y�� ��hR��U�)��S0��� Y��)��-H:���FAf��u�+��10�^l4P��X*[�����wq�� "��%��z�����r/�6�չ>a{�|�a=Џ�а��� H��������ǌ(s�裰��pi�����T���&�O���|
���O�~a$<*��O��NH��-K �yёY�[���~ui��y���T)�����u>~�������N.⯎�0��'��h9>$��WZaF[gߎC�s�h�m�a��>�
s}OB�:��vTd�-�z����wo�m�*��!(O�R��N��D���y_tr;���}4f���n�?�Lg�0UDմ�H��u�I"����zlH�VP;:|��n!�s��Ñ�8�)ft<��#ah��3�+��Tp��.oo��t�f�|~í�fX��)�E�
�;��l� R\r��D��(.�1&^��φƢ׾>�{GT
�����D�vڽ?_��[T�{ԣ�0�vJ��F���E��8'�w����x���(�����
�2QꄓAh���Ȭ���Q���D�����_R�Gʻ�	�lk������?�[MT�$���s������ �QĜ��	P�ݰ�m��r�^x%�Y��\���<Vsh��T���AGI����`�Rь�y�e���$ ��~�g��<�ʽ��/�/�DY¿L,c��*��h(\g�{L���)ḣ�х�����vH�]��Ҭ3��C�@yJ�'%�Z�?�(��U�����4�Jj��]�at��G9awv�T�q|B녔q�ْ9��!���� ���'���W��gv.�������ί�� �s6,؄�k�u�D�M���3->"�+�� 6OM���ie��T�lU�&�|��}���M�g$�T��4�>kRM��MxnT��4_o5"<�ƙ{�N�⬂#���"�������sNٍ�<FWJ��$q*�u�����/v������BnS��RS����)i#xJH��J$t�qص�Q-�_��o�+�i���da3,�7_��T��5��[$�Ϯ=�C�]05
�6��{NC?�q�ߒ����r�_�敳��O��4��)Ԩ��go�M�ܐ~f�`0i��B�{3�%��܏ٶ���xn���b�R%�k�*o�"$J�8�v��Kӳ��f����+�Vxų�J4���>����	�8�E�p����Z�לj"�kýZ;����w�oPh8��a�"F+22��ϻ���V(+���z�S�y�r���7St n����HT�
l��S�ԝ��xj�m(>o+��C����=�k_M�d�ބ����vǾf��Ŏ�qgi*���h�V�SD���~nȴ�T�>�ξ���}�sq0��*&Y%AN�_c�M4BE	%���'�3 �̰�عz˸Vˇ'�^<��T���au{u���h�#|q���6��>������:��
�J�#f��ӵ���I�î��yD�H#w�^WǺ,��>u��')�իS0���ٿ��ɦ7�R��B
3�B3�Tw1��m�+m�Ұ�2��A�\m�W��&�Q!r����-cS�;�����zɄ���B�]s �0��6@v�X�[���ا�W�i�U��m�H.z�m]������m�0��S|�'ͪO��gV�4�8Hzu���/�eFh+�N��W3�?���RUx4Jyv����}�%���6�5ϟ�<
��KM�~��\�'���a��D�Q,0�lV86��6*`��^(��{q���o �.�O�z��C�a���t�R�&|���VE]�	����
;$R��Ke��\�c�t���'�Y�U�K�Z/M��
��3Q�ћ��~��,�P����03+"��&p�9<���#���PW���L�|��!��G�E��-�D�g;�g�?�JZ.��Vۻ����9Z�H7+�
`Ӈ	�*�}a��~���f5B&��^�
�#���6u@d�}�L%���=��l�ī�����÷�Y}k���	TOΫmu��Թ��C'ݫY�7���P*O�����2W8,�V�H��
6j�����笟��l��`~�.T�.dW0���gc�pR�u~���"\�R�&S|�E	ZMN��0-T�nS�5SK��sx�A�K&�Zĥ�,sø�`��|s3�Mۮ�5>�D�)?����S��@&T�+=�#��s0��*!�E����A�� �J��I��}`�n1	!l�B��_w�?p�#[mȺ��w6Z�,[��A�,��i�`��N���j���j�%=�r	+o�A�D���+�B��������P��8�
'ē.�ۚLE����Td=k»�-�El�A',e�%5�u�{?S'db:�Wl�ᓩ]�������3�2��XhP�{�w�Cڲ�#'`vh�hyJ�Uɴ���5րs��V$�� ��ߨ�D�Q��_^��b��8rۀ�#�[�A�7�l͈�ޟsm �7<>�l{,:z�.���
����ӊAڬ��Z��ӊ���3��	��)�B�k}�/@���-�p�vS>�C>z;�p��îBaP^Ӗ*�W���ϛ7)��g�)��o6́�+?1���~u�Ѽ _]d7[���Bh�$�����!a�p�~�]�#����j�hֿg=���7�{�����v�9�����i�������\'���8꾍�R�1z��&�K��ن�]V���������T\_Ⱥ�r!?)-P~^�����uqK��e�������O�b�n��T�1D�p�P!�{�
���d�֤��o� �gq�6L�KJ�D[s|ӝI�= �Ҭ}��F��.���U�&���0\J��A~ϲN䅾}�N�6.r.�^� ����:K��G�`c�Fq��w�2ś�_�^eh	�ӂ���-�E2�� q'�������aE�8�o�����G��s�'Z�Jv�) 7p�-�t-��Ⱦ�]��T���`z�B���]+�;?�r1����ϴ��HFA���z<��CO�c�C���A���P��H�-������	���Š���4h�$l&_5[�贆����I��}���Z�/Lo�,� lz�n9�F�n���լI����w&��		������ �v�g�/6�����m�����S��Sݛj�w8���j��$��i�fxn1ZRw�E�����H��1��9���5��t����1�G�����C�5�@~F�*3��M�k��9*.�G���#�FVB�lB�>�$�F7��S�o��� +,%��}�q`<����<k��+���k}�&�XJC�mJ�p�'CD7��*��ҋ�D�5h�����i�M��A\�)[�E�֩}����ԁ%�g����y8��j�u��L�6�@�0��=��Z�ts]����ڐ|�ʤ�$�u ��� fS�O�68+Rr�V�]͸K=`r��5R|��5o}��}W��rMI���!I������t��̆経��q�+��ar��<WV�qb5�	��̼ɬTzy'#i��r���,�6�h���Q���D/�A��%�^��Q%���Z�
y	t�)rܴ%"�'&�DF����i�h��4&sQ���a��5@��@g1H~�u�K���g�ʳ�o���m��;o���$�g1{�7�)�
E�c��-��x,~�:�	殛;_ 멾eT���:t�h����ɰ(Ja�x?X�r��w��Ɏ]B��&׼��+b(�݅��$����PXu���4����b��:��olx�����Cي���`Z(rx��M���һ�
ğP��r���7�U��U{"��:���g�-�cF���V�NQo���	0�����ތ��o����㘖��d�ia�d�}i!��Nn�t�]�Dݵ�ʫ䗨��Rk[�Rk3S��d�S�+�8[ۇ��s��}_��XEVv]t�ԇ(�K�!! J�,1B'θ�ȁ����,�ۇ��U+�'UF��g�)@r�;�P>;�-���NA���������So�����ݤ_����^l+�A�>�������W�}1�Vȓ%��r��"���R�[��ucU�Y{�M�N2����{m<����e��W���z?2����9���,t�Zͷ�C�b��{�W�7��(�D�٦��m�a�ʷ�1�?9�7N,d:dʳV�9�4|Y.N���oͨ_�����Z��.ˀ��Q	�SI��;��0�L,!n�ۈOVk�Q�����ҙ�'g�$pJ��6�� כ��R��̽��~.���7��œ�^]P��d3�����ӆ.�����k��ߎ�Q�ބ�/���~{�Yڥ$F�zdѱ�ᡩ�ա��Ҙ�++�Q���P���-�R3�C��3��K�9ԧ8�
�]�Ξ��2�
���~�[X��Dh��e���#�E��W3�/�{�±`���?@�g��������:��}���tn�ͯ��HQϡ�W׋�������� /`��35ٙ[���=��sl~�]��b�ni�H�{���y�p(5E9�1��\2����_/ñ
r����b�C�w�*r��	�?�,}�"�t�=:F�ɇ���F�����kV��_�)ӋG�w��N�0���B�?%)��R���ڍ��!���'��{�rB���H��)�E���u� �IM2�`�l̻����P]����>��wk����^uZV{G��ѣ�T�!�����'���9>���Vg�M"8X�&)rq���b{�/Z�-����@C�l� �V��T��V 4�Ă4��:����zM?��۳�hj���<qX����H)􏒇�(Q]�U��b�X8AWK2��B����4L
�I��i��Vm�}D.=� A�2C�Z��ow�}R��A OV��$^K��)�9��ɨ��%>���/!�UWt�3�DѲ7i���Gk�X%��|^n���GgiX9������Sc҇aeAf��~g6�u�7��~��"A���(�-�ۧ����!A����O��i��E��sw'����l�]�CpW��k�N�7�cZt�`,�H7bD0�ؤ3���( �x�r*4Ax<P;o�_�䐀�󂎣=i~����*�u��,���LG���Ŧ0�7���~�V݆j�d<0��pzB���)C�{HP��^3�8ֿܟ!z�A`pac;��'xb#�D��{/@@ ��@����e��F"1_�jٮ�7eR��1��mqn�.���R��	�q�k_��J�OY$�܊�"���M2��e�k�VhPj��FA�U(T�(��@KoFd���>��6&n+6W���a��@t���jtͭ��rE�vI������+��YO��M���u1�� 
��D|@������*�ߓkm2S����L�WV�tS#��b���8����y@X��m�|�_ľ�ŀ7�9=�Ye��4Gf�A%�5�6���"K>ֿd���^嫰,0�^��l+��$���IO���|<�/3�Y�|O˧M=�;^$yEQt�$kO�ŨN�L���A��#��ԖD��y85M��dK�-�|>W�vmY��9'H!�&�3#S*N�d)a���uI�����@��ӤQ��a�~}M���
��E.���Dot�Țp&�Jv�6����8�R�8����,��AZ���e�c��ݳ���>�G�8������#�;��/�eD��=�t�i)l��9�6�_et�Mm�)l��$4�-_�e��s5���#�;i!���!r3�4\��0sA�n����t�]`8���_|��3S��VƢ�,.#�"�� v<�+�R�SO�y��Sӹm�g��EIԶ���?��>9;a��I�9/���gu�"��7d�J\.�7 ��4��.��ik*/�V!G�%`A�/�}ugdʕ��/�e �s�f�Ʀyѥa�m�_��棭F�`	��ϭ�
��ne��|�8�_�5�|�&�G\bU�(}u�����/�;�G?��_�^'�I0���i��J݄1�C
�j���.?������7,>ȇ�����oJ�`jկ�0�Pv}R>Թ���/��iNY* �3	_��y�ͽ��f�1Ǣ�*|��������{=Z�8�%��D���F́m������S:�H��T��]魄��G�༪�'��49�������rUj]i�mm�~���]�BF���m��������U��돦ɏ���t@i�%L}^�g�,�e��^��%8h
��dC�ue������ǯ���	�Bf�MG0�JV �fN[f���N�T[T�P{�*���g����:���_a��>����/m ��WC���]LK�nsrHy��L�J7�ӄ�)�b�e�S;넝�|�R$3~jp1������L��6aR䮳���-٣@�����P(	��4�s��8�	�NM$:ş��N������n�Z�$�R���1Ѥ-/{ژ$�;�ڧ��k.�� �=��ɺ�\���t��8�A=�_�dS�y�"������� �lW��݃nժS혪 6����=�2��6�J��$�+����D��7�V��F�㠹�N٬�OƋߺ`X��+a���7����f�/ʣ�5F��hH�`b���^�ӕD7�'eI����>ckI�ᩀap��"ړ�E��mI�>-��E��>8�*��vg�fGO�vs�;h�L%��ry=\u/� )�l���F��*B�,�|�<|b��<ۼn�%�q�f��K����<�[|{�������p<�5��Ȥ�:�t���w�no�x��ϔ({����Ռ�K(@�����5�T��q���Cd�36g��^>�*`�W���k��ʡ�~�'��S���H�_�T+������Nضqc��Tq�1n�̚��F���0��B�7���;��H��	q���^������m�)��&�S�Z���*��e��� ��ҹ��-v[X;cat�(j��$\ڭx�)�6f)��<�t�Yz�Ԃg�B��~Op�US�`�'�v��ޠ)<����
��UF.�o�6E��UH�ڬY�b���=F�-��|@���փ;���>���Ųf�ҭs��y0�R�n�Z���b!_�V*�X�����O�VX�sV����n��RΎ%
k��	���P<J�,Z-���r�ͫ=׮�e�F\��������#�&�`�隐6w��7L�ɟ��g��p�U
���bܯ����>ak����v�>>�ลt��['R�����9}�?J�������WwvuF��'����������w��Oמ0<#�4 W� B@��3��@{�4�,��
5m=�(��9�.�6M�Xv]�2J�T�:KD�@�$,MĎ�YV3��l�ð)W�1V��q*���ǯF��@�cV��%c\i�@G*�3�䓮������%�w���#>��9k�M*���ΉMYȣ�Ӏ�xU3��^RhPZ�q�sdU(먶�N�u�1��yu�6�C�/}f�4���]��6��d�	0}}����u���~�W�4b�l��m�L��l��[�����ė�����:j0'��UC^4�U��jd������;��M6��S�$������A�Ը���F+T��Լ���d@7���I�{���<�c+��v�l�G�����O��72&�@8��̓ٽx��ϧ�D�w��F�q/k���<D�E��Kۮ�_r���9� ��S�;3W*�>"[kz�� @4�b)=*�N��(�#��/ �� �oK�O̾��0���E���r
1��4���n�s���b�dJ���A�|��d�8���P������<�����u%��N]�`���w����X�k*7������Y�je���> �~J��v�$���@�x��x��g�M������]�-:N��"��a��M��&	�l���f�����njp.�GH S�z?8�E��B��=0 *��<��w��KɄ���;��"g:g"2o.?�&�㞐2]����7��a��.�W>g�]���ª��x����򤐣�.��.��ˇ���.�9���ٶ� [��#Z�nE�rn�,�϶���B�(�&Ƃ�kM��4Ƣ�ljV�-}�7���!����KJC&D�!}g^�q(b	��{`���%�e��>�|��l\1e<L�ZX��z�)\�8�ɚL�u�c������s
�>�	�t{K,�\#�Z�+:ܜ�a��D���Iy�җM��\��(B��������[�+�$����c ��W��c�1� ��?X�j�ƣ�倨-8�b��L�-��+��`�����M|M�${�G�sAi�.��8z"�X�HϊD }����b\y~Q�e�ڎ%��4+%��N5�N���v���Zb�:Y��ݱݾ�q5G��`{kD�z��$?�B�� w|���!hԙ���9_�ђ�]�0G,��%lu}��3�	ZF��=ҕ���ԅ���۹Ё[��/��<T�{�);�Q���ng'� ����I9,���T�UI�+�Uc�>#��+%:�M�\ѽ����S����I�)�����_{�$ms�b���@�-`Mh9���;���aL�B)O�twł�\�zα�>CG[]��:NֆP͍~x���!�G:��x%��O����.�A� ���$�B�7J;��YW���b�P�'�N��N�b~LC�*j?�ǝ�f�yK/�x��`c���A�Y�.��jz��k_����2S>��Sn�����x��U�v�EC:Fs��n�7�f��	Z/F�?0�H�����ŉ�2b���4�2rA�VYi�J�V����[?�o'�����K�}�$��}x��R>��O����<~��z����Y���)8�M��������Hm/(�0V�� ��~4T���!SU�
D��QBMT�a�<��F7͕jg$�o`�,��c�.8kwm	��[���ݧ�h�k=yU_��a]g��^u���h"��27.�5�CλP��_�m���f���ל&OC����f7,�BE+p� /}D�f��:�s���k��2jz��:9$d<�7�2m��?��ȑ���'qi8�����g�Y�� ��|P3R�z���}��W�����Ad���&����,e�r��]�A��w5ݯ*�Z�l��9��eh��T#
��%��V�W����x$O�٤�8���a�}K!�9�����m�V���?�Ȁ7�+i�j�=���*��h0;��8�?�}���El:���y�[�|(w4گY�#ʩ������T>b�1_,֬0q(�\,M�4א�;@].�p[�(a���f;�(*��[��1X�Y�S+����J:lp���{���arQ����h���!C��Z�Heݽ��#���@�2F���P<V�a��E�w_lQ��3�t%E]9K�IlI}ݨs[Y����u&��	��WT���5�e�Xe�S'=�2ZX�	�A�]��9Q����?��C�᤻�-u;D�tr�u!޿�Z��c�K�k/��6���;�1(���jV�ƭmʇ�ݒuP��Ћ�"�6�8V|�`�LQ$"���ʿ֧WJ�`�����{V�<���yHn#�Ҵ�/{��}���)�a�� ��������ZZZl�-��ɄX��@�'�Ti%i@yI��}��J������1a�����QqX4��R���n�,�ɪ^}b�����&��m@��o���e#��1�a�y5@	�K
?/�ԉ�.�ۊJJ�ix0�$�RvE؈�6mC�� Pϛ�c���d�M�!&F���~��\����b�9��!E	L|$�0Hj�5�<���g���3N�7��j@(�½t�������Cm�r4�V�/ZmU<�~眺��A.���8Y�v��*�7cO�v��QS0!5Hم;��s_T0+F]��.L��i4PT}�KS�$h�f��5�TAe�d�ͳ��D[IY�Rr��д�*ٕN����ԭw<��}�b�#�sn^3s o�	�Z�H*TXr����&��uJ𤎉��"�.6�\_fd�~u���v����z�A[7���1ʃ��4��oݜoV#�TA�9*��U�SB>�D���#_�@�|ٿ��tf��)S��q$�Ɣk�$R�2-q��b\m��º��`H�m�Szk#�tF!3�֍��&4�]*�/{!���P"o�-�r[���3�����uȠ-����ŋc�@X� ��Y6���M��6�� "�LL���'<��=!�X�=�8��a+g ��M;[>���+��#w'�{�I.�Xǘ&U6餃|�8-���,Z�������yR�W��&�OT7�W��@&��s!���Kˡ�I�k��Ϗ��'���ÀJ��nl��m,�n�#��R@���ָ�Fd4��0'F�ĬͱOh痾��<
���$��.�\�{)M��3r�X�B�kI��@,� ��BD$�N~�<����a��e֜덷�C�zohxG;Q1�>a���~W��ɼZ��,	~�u����+��G���ƍu/�[��[%���5�i�Z��:UU�B��	��hx���۵0}��a���Yֺ�w<֛r�؂[������1o�wVu����b/S�#���p�j�Z��z�3BRUE�8R%�h�8J �,�Цб���c�o'Ep�������K{���#�A�ɝ�z�D*�8Ӿ�+���2�T�	Y>�=�~>�g�2�(%cN�:.e6g)��~~����9'�	�Q4��"*�r|�(1T<�a��g��U�X�
eef��_��u�:,�'.+P�r�ʺ�zǜUgU���O̲.g�j5�.y���(�rV� �dJ��q�l�*��z����jWUH_���{/4�֭�����|7� ����k�!�$wQ;Sˉ�e�V��@7�	50PX&�4Hà�dEK7��ݛD{M7?t�Z��#�"���-��Ւe���z�k�,w����;��b^����+�)��R��y�w����(���N��[��Sb�|�w�m���q5�����|7��K��=4%vGt�שI�{?�-N+��?�]��2d���cb6��H1��KgWéyJ�����\�|��Z?��6��n�\S�����D���4����i~���~Q)b	%�=*mnV�~
r�§�E�PAJ�E6�/����ԍ±0n��kGn��l<N Q��w��o[R�5j �b�3t�A�`��\������+��JƝB
�����B�ۄ%|��"�{�+�JSR��S	�v�7���ο�U;7��=�P	w����{�?'G;�*�eQ�j3�K�}C�-�����^:����U?�#�0�%��A�t]�&x����@�K)�@$����њ���[o+���Ӄ ��GU�P���4�J"qs��T�A�y����������W��S�l�����<�w�D8�*"y�]���)`��zE��#�[U�(��zc �� ��̮A������*�7e;����+Xb�g�J"9c�8:*3��I|�*�|u[CU��p0<��H_�r��ǾXy)Hlf��n���b<I�&�hf������:F�ϣ��}�$ �_��C����z	�<�!� r���؜o0�x`�vTBd�\m`�!�Wjt��0E�T�^argQ'�t<l��RB!�ON}r�."�F�)��P���?�Q�8/�&�V�ID�E���7�}�bj*��ՙ�O�ѦJ6�:��\�!2C�N])$(���-��@����>��Z���]����$p.z݊Uo��:�7%�h��3=l/����N`���B��߄ge=�+�{9�xuс* ��W	�'�5��Xx�	�>�2����:	�<�~�cƉ��Ƅ�����v�m����(T�Ky�O���N���S�k��ݹP~��ɽ@g�������
��L�z�)	~��zk���j��<���;���TkE�"�ǣ���B��D��F�ovr��J~~���
����Jo��ƅ�\�X��]h���&���,`�4&��E�_�3���c�_J ,8��\����akDY��'�2L\>G���}b~���7�6���BF���H�vx��l�VVy<�l~GA^�&�{��KN?��8ug��:C��>��R�N�_cPdc�=.h2����*d�5N��nB ?'�ƀ~�UD�,�R�A$�J�� �:��R}�r?籌��������9n�m>�.ˉۈ����������腜�����;��A�@
Ҹ�]�m�(�(��U��ϛ`�>�h6���n��d�����6�d"r��։6a�����z����s���q��v�D�4�K�>1�@���"Hb&ʕ+�H�^2��Sa�t��p��&��Sd�X8�°e�8��xɠ`ҌYi��X�Ǖ�oC|�3Fz��Ӫ��L�d����ɡ��|8�<M��#�ڭ-=�Wzs���&���J�X�h���ϻ��g�Q�0]9jzu*�EU��c�����g�TR�;�%�����tC������A��A5�(ڡ�{<�T�U%-�.B0��
�}�Qi�X�0��s�i�0Eœ�Q�|p�Vu�Ȓ��HTF��㠚�*��M��s7O�1r�s�����nݷ��	x�����VG�����.|Os�Mt*�x�+d׳m�s5!k��}%5U,{P�6��%{��L���r-�s�Q^�O\AyND��H�pA�0��L�57�Į��+���0� �J�w�?�jME_��9漜�&n�vp a��7��f��+Z����	0&?$+�{�j���A�Df��?MW��胦#����8�߳�tw}�0Su�	j�.B�W	�'q�TU&�IE8TM�W��V_m���)&�幎�h��O�Up�Q93V�T���:Gƀ�͖�U'�'�@J���uvnJΧ�~�1afd�H>In58���[��VTm`WM�����@r�k~�n�',��j����G���*v�	րf 4z/$�Ç^ ��c���c_���C>�B{^f��(�q��a�B��{KxZ6��f܊��,��_><��ѽ�'�Pp�c\���[w:f����9�#x�L֡�mF��*q����M��`!^���p�h~��&�K��3RaG/�`V�o�M����RpKf|�-]0�L)y�"�
����Q ��jp_\+>)臚7t�(�zx�y��8�T�؏�N��
��yHa=)���q��{��P�T�J�)j���8:�>��;2��>�"U!�V�B������K���kI�d�s��8� Iv�0�� �Vy�b�l� ��SxS�kGv����+������2��u�#ܠ����}tܓ�~���S�?,��Om�9�YD��W��R�7�e���1~ĸ�m�/��J֎V�t�͔�,���:j�z��M�9d�2�~����-���i�P�sX_ ��g!|�)�|,������<��¨&�c���:��0F�ҕ�z6T�gk �+��یиo��DG�]º9��v����";y�4����:c���rl[�0t����Ɏ[t��ύX�I���p��B"��<x���\o���;���F�?��N�y�,�d���G���v�n��V?*�o��8$Ԟ�b���B��FlȺ(X��j6�ܟp$��P��k��Q94Ĺ.�yǦr5bn��	�k�i��o"�D�	�T`�SÈ�,k)Z�&��v�����oV��ˍ��(f��J]��?� �M��D�0Y%�Cm3{�����)�-�F/�t&���t6z9Ԇ#��L�D���}!�T8�M���׻kA�Ȼ�K�]vn���6�<�	;�u���,_p`�Y�i�	�6Nb�F��Q�B�u�ʬt;U;+�#�ќ����w��z35����+��l�~���:��ş>n1����E�(9'Ađ�0EP�`L��`��u$��ā��+iU�=�N�4-�h!Z���}������_�X����&H���gM�k�$�^br�^zld�/ڄ3�ϫ;{�����
1��dz�&����>�h��W�@c1��Ȫʽq8���H������'S�3;�u��DK�"ڂZ��Zٜ�W5�X��ȸoC{�I����6�K�{�\���fM��G�M��R/ݞQ?�E�7�o~�S9ѡ���S�w��������j��5qL������Wq���F�ü{��XR0���a��\��w>B����ceP��a�Xp��# $I\�u��=��cn-�rc��{��4_J��_t���3	e���A���r�|{��>�Юs�"��Y�7f�U0F�t���B�tQЬ6��Da���WE�gd��Fe�[�R���^��l�,��G��ATyވIW����S2b�l��8Qbk��ʰ,_�)ѭ�kÿ|]	�)������H�@���ˋN�c>�_.�Z�q�V�E�`x�(�{�ǋÓ<-�=��ǚ�Ir7�<B@���\�����,������kD�����D�$>����e|���|�1N��fze�8$�B����0Ca��:��ǶceX�*�ծ@������N�)xB@7��WO���]�+NR#c/��R�II�a�ךOe.D�|M�a�H�lk����^m޶�<A�)Tg�{2�Ө�ۀx��x��Ԟ]�����O�Cg�;R���{G)oSʾ�ߊ��!q�Һ�,K��2��#W��ZQ�]�nCz߮��>��d T��`�n���v�W�X�	��H}W����!�8�	C����;����i��^>�(C����'���@�A�҆0�7*ߛ���[�WǟߒR'�
�����9��?D�^WV�]O������38u�n�&'�`��)��:^������TF�5��ՓqXjcg�a���/䍏���j�D!��8�=�}��f�QKcK���I�)�9�l�_�s:#:��j��Q���T% �T]k 	�Yn{U8�5���?��.l\M^^U�$����bnZ6B2��n&��+�a�O	�{	Ts,�sc��$�J�\�g�*d�;d�����[d�Q3���ҽ�|��4eUc��zL)dr��i�Y
�cO��^�q��Q,��*>3��5j3T�kM�.v�Ϸf�M�j�����䨧��#�����#� ��|�-V�\�P	�����GDm�T_�X T�_]�
��^;0u��-�^.S�,_(b�_�	�P�ƒ%��բ<5E9�-!�ó/t��L�u?"���iM����th0uj�:�ob��	��Lc	Gze�V�������x,S^|�T�}qx5���>Gq����'
���C|G貭/L�r��X^M�"?��&�[�{J�>��H5L`�i���^��2�0�d�ogTq���t�lϋ�sڎ[r�	�-��2�)�/��"�F���AC�١�xB#a����k��9�u}	?�*N���E�:S%Ύ��Ӝ����h��o�є�۪Gvr�OP��s��tG#�E=[^1�H��$���-�ċ���y�r��4ϝ�Ԝ&�8-�g��C�J��U�|�x y�G6���ݪsړ,(-X���X��{�����}�2�/�T�����|�u�uR���'X�5g�!�,���G
E�H瑯��+A�
�#��j'�n�L�ࡡ,��v��ÀnZ��(z+<�)uj�"��aBK/�-��W%1�4]Ij��>H���%���\�f& A?Cs#��᪶�I���U�����ZH-�M��4���Mӱ,e�uȧF~ZѭO�>A9�m|���mꊚ�O|qV?��%�j�+F�!�rsu�MSkC+-;��r��'?CŃH.kmH(x� �Z�I��P�:e9ҙWa*4���C�."fU����#�(�1�}.�T?��&�.ߗ�_�_�r"�?Ɩ&���G���(�}z��&ɕ��&4�$D��R)��h\��m[Sp�21�� ޑך��ʖ��{.�zRZ��Ā�d�Xz�ȯ���~�Nyr�og�O���s�t?O�T�*�m�#kةo��X�/hs:��G}#pb���=��6T�/i�7N8wڐ��ޢT�@@M�rT���=!*l%��_�<�ɼ�?��&��co+Xf�xq�'}�{9�J��'9�B��8n����d--C�� �7=pb�'Ԅ��k�I*�� Qh�@C�"VX=<��׍�/I�n�J�� qg�L�1��L�����W���)��Gzs2_���ef�/�?�C�_�א��fh�FA9�a[� �j�A��ų���[0��(�5"
Q��CQ� '������T����vd!����V����ߣj���9J
^KN�OB<�F�N�����	`;����9w��G�<k|]FHF���!���eZ���o�"Z��
!�bGQ'��e�Z)�474����ތ�."�M����MU�+8���9p�	k�0X4�!�0�[o2?�:W�KR8#ƫ�� ���	��&��9�_�7��){�a�8k\�b����Od~�&�	�)!�����жZ@
�|>�g\����k�ź�N���;�#�q�g��pl�t�5��V�,-L�f�Ml�孡~����L��������{ƅ��c�7�p>�;�S�~e�Qݟ8i�b
X��ҿ)dCő袀�ϗn�?���YN(Y0��������Z&���nF{��Q��ڋ���Z'>C�`�M��\D�)+�p𠇲7��0 �ã��ۆζz"(��4����A��W��/�2��w|��Ӛg�`Ҡ��-b<A�4�XZe�K�vS�a��g���b|d�$lg����(ׂ�-����:�!����`�~E�n�8�C��p��˭��ۏ��?�WKT|Î݂q��x�_T�)����/����w,(�jм����F�Y$O��k��k�'�'�ʂ��Z����:sL]^����ա	I�.ܨ�
e�!���H��cwV�ag���Yd2EY�'�E�%���~ h��	UW���X��#ČB��n}�U	�8�L�H
���:,�mt���U;$�|��`�jKb��o���|v���"���w��5�Ȃj��Z4D��y�����l>-(d����z����{L�����fa췉��S���۴J�Qʀ�@�����a���r6k���¼�Kiq�r�a�='��=a�d_���K'T�W�b�g�ڮ=� }�7d���,��1��s01��Ѕv_�m�NSY+���$����a�D�_l��N��g��)����)�
ɽa�L�'�b�`�~����	�fݖ7�9ƂTm�ڧ�祑�_�Z�	O�#����#f�9���6���$�Z�!J��i_<�ѓ=�qa���S���Ph"K��ͳ��!=f�*����Zr���w7b���2�}@�Ĥn$�
e;���7�k��y[J`n�GLPL�qQ��E���Z@\0{;&�m\<2��Y���T�m�Ė������'�B90Ռ����!��k�e�<O�i�P\m�=(,vMog����?ne��x�l�*�|�-8��r���9�=�@Kv�8���T9RSSÇa	�_��,o"wʱn"����t
~��~R��Nu[�6s�SC��4��_����� �'��+Ƭ�E���<��k��v�Fsu�/<ELnITVW���IBqw���iH�	T��'86Ɍ�>��D��yJ��D>��k,�p�1Yn�Ձ��?M�;���w�a���fv��_3����u���b����yO���F]pax#��=M�^�͞X�����;�+���Q�+��`�TH6XY �o��\7��{#�o3=�pt��u\)F�p�1ǡ�T�
K6� ��o�$����6���.݀�ym�aw�ל��,��[��s2^�@v����'����H�P�&xg��ң8�?�u@��qdd0I�6<���1�ܚ�f�Z��)~��m��΢c�D ~�(>��f��:��x�G���~A��?�I���~��"�uӫ�9�lz��g�A��i���bʇ�����yed@\|kȒ�5"cd���/���?ÒyM���yv��lV3�l�0J�0~BmG.�����$l�d�<��@g}���;�����EdE���w<x�@#�6$]ͱūw�C����aѸ�q�n���B�i6@&��=�"�O0E=��`�=P�Fq�uo�{���A��E�IP9?|P�`#�ǡ����8Iti���dď�)Ѥ�j�D�	���q���!��R�&���S�HW�0D����_3@'�������p�$��q���Y�$�[6�@3vaV��r�cTȩ	 �幝�~]MS%
n3�ʱЄ��ō����e��ݚ ���[�>f��َ*�����+ؚ0��^��8L��rUfT�E&�~��S��d�����Ak���̕ �} '{C�z�a�Q�6�����/-��������"�Д��ʙ\n����UM!�X��<"��b�_�rख़����~�V��K��m�f��B�i�G��
I�s���X&Y��=8���cG6C*H�v���">��y�d4��et5) ������X���� �w�b���ql��>t����KQN�u���tW!(�]�N�-�)�v�py�c��6�@;i(
�:vN���D�v�QK����CPXg����������(�N��!�8Ճ�L������;IN䟬�3R�d��p�е?�mu��Qզ	�P���T����Ӂ�9������^�#3�Y�\�FV�"��~�t���g��R�f�\��Z@Wx�����9���v��<#�0�����0�
�dR7[��Rܠy�oW=	gQA���}ߵ*�G?%$��f��iu�p��RE��6P�v�a�,��Ce[��1(a����@���n6깓# �4�I�e��&���H�,6I�h�����;���EE�RG�~�x���k��~���wj���ZE)�@�[�L���W��W_�bO���>�%��l��a%�0��-��f�z�����!�6�w��1��nܼ��Ͼv���y�*�N/�iVܾ���KԢV���}�B�))ͣS�sV�7���|Ұf�������%�j#vR}�����0�����$&<mz�*1yZ���A�ネ6�wL��^`���\���"])m�&	6,��HV�e�	�``�6�E�ե�ޜ�a��u�m[�AT�TO`��B��Y	
����Z��/O�����A6�QdU%_}�mC�� v�D�l	��^R�����X5�U��*������cs�7�0̩ȓZ<�"M�kD5D%�Yȏ��z�j�Y?:|\�~6�ɹ��5s ��i:/"�3,�Yt�]�ܜ�/
 Xף�ܮ� �&�#�� �.��<?�go�yi}�n\�9����&��	��̚�і���� 6����
e�YG�s��H�,E(���/��7<	�Ij���L����ݾ�3#��?]v��I�ʹ�Hb��;PJ��H��'����O�u��@es�9Z�����0]��bY�]C�sE ̦}&�n6�řs�'Ҏ��I=pO�J���5R�ië[U<o�3;{���|}�,k�Vo��Κ�+�A��'�kKf����S{^�ܫ5\`�4�=.����l�3�3T#L�n6��Ջ�#��Y���N_�b\����^vv���j�������j� �R�D�i]�@t�hl�*��
M�!t=���Q�3t-��y��|�&~�|Kr��`y�a֜^z��+�~E���-���<���Ɖ�GU+!U(Na�j)8���'�Rr�G�V��+��r�cT:^�EDQ�Y�����EG:��4�!�->�Tra�n�}��������O�֡Ti�r�$��z��?!&������E�`��_��t�cc�L����#նX�ה��������±	�&I�?F�		��솰N4\�X�cj���B��� �`�X�������� p��*֬Q6�]�7/�L@ɉ��8��qƕ1!����@�Z$��ފ�f���_����W\g<��(=-����Q�G�h\
��́clƁ����4KD�W*��?�+>����:�dE6������N�~���,�������V�U�[����v����ޥ�\<
���0;�S\IA[X6�Z�	ng��5S�o.�2`,�)�f(��-���B�듰N�^TX9��Z{lb�l4��Ls�5��g�/D�Y�☾�ת���J�o�O-Z�쌢S�-�����w�,�BAO!����Ty�����?<������Fե�Wi��=����;�|���}�/��B7�$j�ns���Bfi7qO���"�X�Bl�.{9k�Qs�:O��T��-�Ƚ8_V[n�s��`���~Zp�7�t~۔/��<��r�Tl���+�n�đ>�l�I,�P��m�\��ټF tzUQY���  Pl
�n�z71�Y�V���2s<=*E��ŁA��^_���b���P��H�^������ߤ�2d�c�龎!�a��MO�ɮ ��u<!]*
�������9��(�AY^�̓/�!�wU���1�$S�d��J?����dX:I&���(<��� �Y��C��s��`+9�����=M$�TW�w �8K��Pe�����c���{�m�!{$�/ȿë{���Z>�O骨�g*���u���!997��]�+�X��B�j�s60�e��~'M =d�c%� {���g���Z2My%�U�6��
�h�T�ʡ��I�2�������� X=Ԏ�7��c޸fSp��iP����I?4ꢇ�)����Y.�L�D������#x����4�i��p-IKľC�ґ��8rj�L��\��^k��{�%�x6�4K DX��.n=p]x׸J5(���{@k��>"H�>�h��«��En���1�G��PZ��7�����MTnÜ�K�� >~{A�9�X4��-��v�ir:�l9qv~	�\������)#";��o�4ZrD&͗ڲ��+�Q�/�:V|T���d�N���&_.���u�Pꮓ�'�d ��=2:M|}/�9�:��t��o�Ÿ�{���:e��6�š'�=AL�~|ceڤ
���TeL��i�#B�b;�ͤ�{�1�BѰ�$D�#�>Q'�ެ� �j����8Y�Stb��0j��L0ϧW ��*�>ޑ���INmٔ�Pπ���d��୪�{�w��s�Ĕ���@�C��#�T�Ŵ�t��$��=�����4��V����^Hi˿w9��.Lŵ�9� x��:T��uvD]�EW����[hL�zSZ��������5�����#@7�a}}�@k
�"$j)26C-gRSGnwK�Uv��rEM@�*EÅy�Cb,#$q�$�
%⩗��_p�r�	v�48c���r������U
�mJ�;��ZW�w��r����-X���J�R�e �!�X��S�^�%4S7�����1��F�9�I~o�s���t��!���nrU�@��o�q�cR�-j��tv���ϥL�K�{�- 뉳���31��TO�P���)��׹K�K1���������N0���M��&�W�Ԣ{�xjc<��b�X�,����R�'��Q�Ba�A�XWb>�یV�iB�l1"�P��=ͧ�.�!W�d�@�y��^�[�� �T����)�p>���;	z��p�O�9a<��SEq���J�&�~��;���/:!6c��H\�uoaֳ�鱔5�@��p85'�$�J������ɑ{���3���;�H���^�gge�D	���*���	�A?.>���a}T&'�����>��7slj�m)"3���h��X=�Ǥ�L{��`/���FPk��?`x���6�dS>}ψ=P���%(!0;U�9�Yy9�=���n�C	X߃�Øw���̘����SZ&�n�|姛BUU_o��DA��nw�u,o�?�(�o�����3s|I��+H��vta�1���2ㄎ,�z�ӝ6�QF��S��mUO���֋l"Z�FFe��%��_�l�kl��Y	���
�������|�oC�NBq�2���R�l��a
�q�>���a��|w;�k�N��������ڜs����L�6'vp���ʐn��j�j�;_^�@!D��S�_!�������YY���j�PF��E�"���UVp���ߏ��l�T\�'bAh/�g=D���P�ҟ���%\=h�����ۚv��M�~�E_���R�|�AEW���&�{��P��av��C;��1���0xs�u���̈�DmP��\��P}7@����\�;���#�sQ���6�܇��MQ���<��\��F�^l�%bO���#tGGp=szװ�[Q���u�:t�����bnS�;���� AIޱP�a�5N�7؝��0����0������"09N�����/�fx~���6��A/|R$\�r?�4H�6�a�|�Ղܬ��As(j@���G����b�I��d4������MJ�����Ҧز�wE$�6��(!�<��+��=�i 
y�a��4�;��4*�?��WC���$�R ��9�E7�"6"��O7���-]��Q��.�4�����|X�ͮ��+�{��Gaxɷ�, ��k��([��|��XY�	��?q^$8���aQX�Nu?д�q/�A�b!߫�J�|�����^(�Y���Mlֳ8h�.�n=� �'��4G)c���`7�^�ǙC	W�ߵ�"�:J�R5>�wMAMX$��ثgX1
w�Eƈ��#�t���6�$Em�Vq�:�l�Ν%�)~�)��̆(��co졘yZ&�cZRh
�(W;�r�%x��ԝ��<��v�C����،2���A�FzJpl ���(�2 9�ֳ�H|@�Z�1��&wGb
4]{�~��J��#�g\
�4U��<Kt�{�~5����`�: ��� ����&M�!o�+�JO,1Yk��j��|kf��<�)a������olq�NU���ca�-6=�&�Ϭ�_��ٰt-�@��Fv�6���۱�U��8>��;��F��)���1� �v���-���a ̂�p�U6�_;��$7Ly8�2���g?�Tϳ�Y2���ݝ�́���c��4F ݶ������z��ATBB9H��G[�+�8�H���9?nH }��]Õ���J��J�4`�#&��+�i��Mܾ��MH�\�����Z�nm]�=��/�S�t;�J�6q�`_*)>p��	���m^��ګC�K-�A�ץ슱��ɩ��4���O�8@�� �����>�%Kd�z2t�a=��o���BB��,H�r�?�ߒҾ���ʍ��j�)P��W��$�=��T@mT��S��dk�Z��dm���T��l���,��Z4E�o#������ع�vTC�+�X��G	J� ����\��>��A�o���P�z�چ]�~���B���vk�2^��+��ML��̺��Y��a՝����V��rޓs�����_Ȓ�h�}1�谲t�ǃ�/�����͉�{����,B7E�~Q$��Y���E��]X�&�����Md�<������B���5�\y��,��ǣ�`���������«�� �H�B��pMf���_S	�YD���D��� ��D�Z����B6ql�e�v�sB�T�2c���=������K&r���b"Q�;�����7��j}[3���)Y�Ia��\�	G;��D	�堶{@�_�shK�ĥ����;���I�-"םqc�n0�C��cϲN%��`D̻��x&(�/�C��z��"�*��?�奀���w"���Ϡ� ���������/ X�?�����qS�"O����E��|�]&��Y����E�j���L�AZZX��G�d��g��`j#��#�[�<�� x�qўC�c���t�+a��H�6����{�"���x��M��"�C���2�湟���_��,Õ�����/��;ņ���|
*Iܔi~�� ���t���Ě>�7��v@���{�⸜F��ln(P8��m�y�d8�'�v�\����Q@D��y룂�;�ٷx[T�jxw���1a�o��n��ƥ�
��f=�B��x,9�zQI]h��w�v
����!�nl�6�8��z2`�1�eN@��#�:N�>$��J�HS�j����N?�;��}�b������i��'�tה7wi�}�&=�3Cft�[K)�!�N�<�ߟ	�	���ş�S7���,)�0JS&"
M�w�1���𒧡c/�%\���4����/^���"0�򨟉�
׭� zO��{�أ�v�V�ξ�qX���m�k��g�g>C�m�۳�@�\!2�H�������٪{�u��̹8�CN�[:A��4��B���V%,�F#�����ݭ�j��0o��I�� q�=�P�dU�u���\�L_ή4�:��NN�%J�J��q��:)�统�qM�p�J�.dL�[�������n�>�gz�d�G�}�4���}�v`:��O5���N���2}�7	�\x;N@?��!`���/��?��K�B����eL�P>�����5|�� �/Qr&��l�[e�����A���y���H��<���a��8n��ً ��Y�� Rd3��/]���90c�c��z��/�A߻(^,�c�5L��Ȥr��O���/�l˟�ˌ�Frʡ<���J���V/���z8��6��w.I���iw�ĢU���e��x�S�ĩ�hVv�ݮ�a�X1�޴S�]�N��H"
��<�m���TU>m+"�O�Hgf1&�H%���52]����_�^u1�Y�{8$�V�H:��UE�$Ο�[��,�����.��{[O�D��TP ��(��6]g���+���8i���0�O�4ɪ��󠔶�(�7AF��m����-��,�*�KP��K�)�T�(�5N���|ݔ����x�B���{�
���AO~���*jT\��ʩ�sN�\m��Z��v��5�RnkJ2�͉4Y��ڋ8�?�%�6m�p��!ز��H�Vd�K�N����7S�h�ˊ�e�lp�	��|�pe 
y!3J^����=]�ׇD�3D�mq����\yy!l̠��K ��]�K��L&�{qa�'��V��fMZ���"�Ӎ.pf�s)Y�m��R�&V�/���R�Yi���n�1���B��Zv蓒������#0nӤ��+V�!����C��/�6<�p��oG����O����ض�c���pաN����׵�v�h[V�A����:���6f��fL�6L�~��\� f��x�/���
<��Z�[�o�}�b����ݸr��ѣ��]�YV��*���5����+ع��:Y��<k�v�~�.�6��F�%��,UP��O&H�E�����.���=���*�U&���[�i��[
!<nm�����|NH]���N=�_�%�s7H��&�z���=G�Ce���ykv���CL���7.�Y�ߧ��!
�Z``�p�3 N�L[�����S��%W-��Z1����/����R0�%�Կ���c�B�/���"��uʳ�i��/3N�'�$M��Ց0#=n�CaHq�r.�D�缱�n]���:����m��'e<��t��?���q��+&*z���v��;c�V���3��Φ�����"���Oڤ$˸Z��x+#w�Cǩ�[��4U��g$"h��� -��M<:0��O�c��yjmaB�+;�K_��r��;�������9m�"J�G���ʼJ�1&�����q����! �~)�ǉk�A�����ڤm7����L��k୊����6yz@�I�rM�i¥4��W@�0�O��أ���_�e��F>���>�-'L��\�+U�N2'y��W�6��[���=��2�db��{\|s�6���AyG�Of��L��2�kX���H��֐�+������F<o;����"܏iC*o��l�*�$`��gK`a�t���%r���֨�$���=��}��C����U1i�C�`���j�K
�(��`3�����hB�xLD��+�~���R�g���3��HE�b:��J9X8gXK�E
���e��!]�*�G�� ���Jr��d��]�/�9�G�|���	DE��\��H�ה��͑4�M�h���K|Ra�
/hu< &�SY��%�-F�2�����\%Sy����s�*/|
�N٩x~��k1�\ri������v�35��T|]�����B�"`}�\�{��������������&y$���H�0��H��a�Sԩj�|=~���D��ZܳKTC���TP$#�^G�.�'��G�Ct�"�2S��׻��I����,�������˵�7PF�j�=�$��N��0Vf89�Pe߫�*k*T�%~>y!��������	��:�"�j���݋���C�����a7�_"��>?l�l��N&K�/r�==UQL��Qq�^ʒ�a��8�A�O��O�2Eƕ_1%p��0U�F˻��g���ŒLo���&$�Xzt̸TB� u��D����OV��^(�/Ew��~����颛b�ZQ/�r�%Oߙ^_m���[��<��<W�������1�<0 ���6��7��<����V8�ۀ��Xcd��B����]�2�YV�:�����-g}���b��u;��*Pg'��\s�F�N{�'��ҮV]X)�֋U���#LR�HH~�"���; ��r	�@Xv�I@eCe9p����\��d�=��e���� i��O��4�'Ng
˩�7�^�m��f,l��	`�'t�|I��x�Xi�Ab�������	%ղbes��� �"�`33��a��,*ӵΠ�
tS�C~���]��d�����w̲59{�<=%l��]��f�]c���m[�w������
q�I�i%�?U��O�p6u{���&���Be�0a��g�U�54���Gj5��j5O��^� DC{Wظf�:�0 ����*��˯.Wdư)!%�c�$UuK�o�dha,�b㐫\^�/��7ݶ���W�$�s\�:E��b΁�z��a2�]�:�3,�]��ك���dTE�;1�fC���F��oc��y�Ǌ���Q邙f���ޤJ�����'��o����>��@�;����BHD��#U���̕3g�p�B|j���O�OÅ��[��lՇ�`
_rû`�5�ژ�)���j_� ����a2bg�vƷ�o/z�ʝ�][�rtڀ���M��y302�o���s��O��=��z6��N>a��Ɏ��� ��`S�j�M}�;G	�{�n������C5�L}�f����uZ �9+���Ը=��uD��ܺ�뗘Bj��ض5Q��1�l�{�:�Dkh�~�NKx��x)0U�!��~�����J�����'!������.J��U��9^�+v�ݸ��L�?�q>Q���;`�C��_bSv�������S-�����
%�IV��ל٦��gx䄛��-w��� 
D$>[I�N�T�����-nD�|�{��(�]�V�xI�Uq�< ���U���#�o�2!ʪ)	e,68֗nX��G���4G��p�L<��r��|I�i�N\<(,Ɔ�f��v�X<ʿ����>�����5ח������m
a"�F����wQ��9�B���wE�#Ϯ��6�i�������dR)�-4��@��f�n�\�[1�`����A�4:��Jm���T9���ېf�S�/@��+$3�Mթ$g��!ЫN�'�!K�=F�L�{����5L����f�?�hV��KW��\�`�޺n�E���J��g_��{,�G<F�|��,�Zr�fLqM0?��{�E����ߡ1��y�+x��
����I���z��2^��&qm6���f9�x?HF#L�8%-��ނs ��%h���k���H��G���o�0-�9}E2�8��$G�@�)4u*�z����c6���mx��37���8S�L�,	�a��J1�]/M��k��Q��[�E��W�_x&	����qhOD��-wW�:֌׶%H�a��˕^M�
|��O�=�?	�_���eHx�c�I%�[�2��	�����8A5�=M35���@:_����A���敏�6�i��`��"91����}^E,!ޥ�l�h�ā�:���$a$I�i�NP����]Yib�}!��j^\�m��M�/H���c����Kp#~�q"̈Xu3�,tA����&)ؙ���v��1�M��8��0���cDa�1�!@����Ɗҋi׼������J�b��3�퍼=_���i���l�I��B��{�:�VcE�C?t�0w2m�o-Ki�69���6��b��Lp�t��'�DW�P�E�����7H?�����'�fCe�WL+���K��=(�q��Ǭ�ՒE�b������4.�Z�����%��Z��N�V��}�l���i�)#t����	� �8'��y
̞7�K���#r����L)?r�y�3���H�1 �p�C���_�����Ry�9�8�0		���b�}H�2�R��;Y�O�&�7���D6�����@���Wq�e���=�|������P�6�vkR�..��&�W� ��`h�����������j�[���p)�NЂ�<���S�PD�cB�Ga�'r�Q'S!6����-R �~�;���g/&���S�ѧ7�sH# ��c�9���ib˗ 	i}����y�}gŒl{*Vǧ�ҋ�fk��(��%�瘓J��N��5β;Z<��d���?��Li�^3w�k/c�JW`N'nj��G�[� �!��c�Dnc5�̠��ofOw�S�'(��B�]A�$bګ�|���s�8x����X�l,TF��PP���0~��%�kj8��0J����m���Q!��8�4�o$��	1��p�ܶ���W�<�#m S
�^�*��M)�:��@	�O��]�t�`�;v�H,����F�9��"��N���i��Pi&���w�O��V��Om�:d4BԒ��*�|���K�J��d4�%��_
;)ա�ȌD �$�f!7Oڜ1Kě�N�y��W������4|ܧ3�<.����=� �̋^v��8F'2�;_�mh�$��Y��
�]�p�Ƀ�p:��$��}�-�, ������z�N�h�p�I�wKE��	���|A�;(��\��V����1,&���lR�N���忨s��$ko9�ע��A�p5�^rX�a�}�lC�6s�=w<����!��F9��V�LHB<3MvK73N����|O[�|g"%1�����Hgq�e<�B�Wl���Ѿ=ޥ<0��U[ 4�TFj֖�������;��e9���D_`>��݄���[�����b�Z��b�Uv�y�AJ��C}'%ƭ� 5m��o�Oh_#-C	��z�5�1�<��}����ٓ��V{��A!��Z��(K!��>d��Q���%�`6m{�;8������7.jb�ƌ�Y�hU��L�%??�t?�j��[����C�;�8$�����9w{���S�?�X��x�(��f�Hj�}_d6��}Ϻ�l֡��!�4<��\���}�J_q	chƱhk�Ѯ��om�'�<����7�W�l'����4C
�W
����XC}F��Ɋ��ڄh��|�v��e����^���'�k� ���-��j2�B5�%&���3#���-�;�mbf�0?Ls%��ί��c�MD3��>Ӡ�;�^�Q�)�����p��i߽���D\42@(�+y�āe����^��t��/�^��^���T�MG�cV�������z���D p��:�?:����8�/B�?�CW\)m\^]S�����#�^P�l\���$r%�y�鲦-A��3�}�ؔVS�J+�y3k������<۬����^�� >�m�X�泑}`�z,���İ<�X�۸\N�(&�8԰08��=(��ŀ�p�r�DL?e�j�,ܾ���Cԁ8uc��Y#{�F�&b<����W(����������q�4%�bǥ��H��8�e]IU����>���gα�h�M���G�#��{7]���1��+Kk.~s?Ƿ��I��Gh%�'f}�WK2� o��ͣ"�BUA��kqa��
�ѐby<�a�jA�)�1�k�	DxdN>��g���
&�iB/%Y�k0x��N���E�lb����DN�m�=L�~�"�'�b�R��)1p�w[$��GW�x�a���^�����`�~g�wj�����Ȧ_M�V�kNg3�}��Ǡ�/�~؊�%h<@ǊI�z� ��H��T96d���J���'��m��l�h�S%�hM���͕����	��@�����Zq�����?�u��.��!*����f��}{:_v	譏�H��s�E��0!�Ʋ-Q>7��1+�����ER��
.�������p͊�.�.�;0�)�b��[ ��S�b���%(+���̈N�u8H^��ZiA�,˵у8)lRe�e�R����A�qŎ{NC�Sۺ�陬i|G,�,'�x��ӯy�7�DEPa�ZD2s�uI��Z0�6�����TR����s�d����
n��ES��5!��X~WXW괽� ^wd�;z����7��Q&��8Ue���	���R�������*��#+l�y*%uK�&�Z�_��5���ԎM�w��׼�"7����{�|`#w���gߧ�Y:1�kz_r/<��	�GIS�ؾ�
#����-v����#h/��ǃ&T/�Y�3Ɯ�'�n�j�Gψ�7��f�&v^lmWƯ<r��9�t�:�;�x�r��$[�t�Q�f���bo��i-���ѷeҝ�������ƫ��3Z9]0/hu8���ێ.�P7{�CG��7ؚ*Ʃ�� ��G٨w�Q�&$1z�0�X������YɅd|jn����"���<����d������!�(�:p�BLPwN:����!<RM�#t�'k��(\1ǿ����J����h��|Uh(M%�q¡�>+�/�%�
 �#��jz�Ro��׈���,90�I� �n��ED.0	~[gg60M����t��һ�E�
�P��fe��}� �1TR���|��{�\~N�6�	��O�����a�G�[�d��%~i��Fr��� �X ���bE�+�W	i~�jx[��#% ����������慔W�����41?P��%�Z��­�d����3h{�#��R�"R���Z?H�#�v`�Q�c������9��44��ǥ�JP��N�����ͧ��>��eH��N�K�j(,�*�6�wH�*�n�{���BZ~�5����l�1���"��:u�ͪͼ��_6���$���2���:C��&
�Iy�Z0?�����c1VZ�\��2�5�k �6�8)��͉��-q�B��ԓ�?޶���̩{֔�VS��a�v	�'W�����t��D�4��R���	)�$0x���~<��]0�M?�8�s8M0���B9;�E��;��߆>Ӊ}K���v���E�2Z�P�z���p�ЛF��KC�M-K8J`���J�G���D�������u2QL+E006��;������e�<��5���D�H�M(~bY�c�c�2����"CE`����3%����gQ� ��4�:�\�ᦝŉ��O|q`�P#�����
� ���_!mo��(��1��i��7%�y8T����w|NMܞ�j�5;\����6�#�-�g�&�⏅Msk1 S���2���_�ɘ�gA�KfB�c,>*�ƿQ�.���ϭu,���]f٥ho�ݕsa؋��,�������vX�6=���N����a
��5���;uܬ��`<��`W]�׈H�@W'Am��zw�ՙ����s5w��c�Y%I��6IPSg�� �!�>��}@��0���>�쯲�gO����B.�������|[4`�&�i�.ȃo�Nҷ����쯋��l55�t�7�z��>�Qv���� ��q�iէ
!��Xu)���Uζ��
���Xt�#��F�ty��77�� #�~��Ggv���ӷ.%=]3YY��Yc��1핿-iib���6=5yM�M�、-h*�w��g����ښ?~~;.��WPR����0�Uc>h��B��(v#�t%Չ^�[e/�������������k��8��mlQ�?��O&g��w�-��z�q
�L�?�ƀ;��	��p|M�v]d��˟�O��~{�h��C�s�A���Yj1�}�ί�Zz�4���%���J%Ga��%����"����u˨{Sӽ�D$U��M W^w��:,-�'W���C�N�B@�P�K���kg�"���"���;�~���	�_��sRb��%�epĴO9\-��JlJ:kbF��U7�`�ypS$��� 7�تobP�'�4�^��������f3={�����}�c�T���H1=s�Sf��e%�D�4��FM���G���}�=��%w^5����#,f�Z �p��A�N�O��L
5Q5���f�";���J�*����t�u�EVQ�
a�V�,�m�]"��6=_Ԉ?��G����8��1x蛋�w$>!�#�����R���f�I|�</F=� ��x��Eǎ�˓$�)��se�hA0�.���*H"�`g����sطO�K��Q2�,@��h�rcZ�ɪ]*'g\we?�!�K���2�l�����]�kW#<0	Qơq�-<K���-�J�g��7�;�>�	�j7�ht�q�9|���^`@������'X+��EM�¬��e�<u�-Ǜ�܁F�����1(m*I=���8W��rh�x�M �
����ߚaJ�"�<�1٠�Ԍ̓bw�ɀx]%ď6�����/�`C����;��L�~�g!��G�� 5�_#xz@J���jl�E'�����A�a=��0�ړ�Dui�;I��^Y]�8�!B'����I��#G�೬���hw
Aԉ��{c��oH��S0���]W�6,A����
Ir�qP��o�FhFy�M��5��r6��y��B��+�&�� ��kR���}�a����Q���]��^ێ�	�'���Ф��=p����Q��>u��A�gɤ��N�%�$6������D�x��W��8��u�n�;d�d��E�e��|I�H�J�f����_> ��);��Q� ���:�����/7Ҏ���_i^�+���{a�eR9��:�c��] ��&�iAsBu5�r��"�t�Ol'�=�����aӂ���S���v�O^L��<4R�z��jG�c�i��=��_���,����+lJnÆIH�"3�&�@{���
���2j<�v�_Ҹb�\U�n�k6����өcr�\��W�eE�&6* �e҃��$����c�E�Fe��y����A|Oޠ�2[f|�q��Cኪ%�|�_��ͱG;�x~{�7ZtBu#�<��B��\[���X.������ؼ (¯O$�!E��%�K_qicҐ�Hw�J��k��T���%)�䔆�ʚ)m�3i������㏼��*8Ҹ�ڣ���p��*�SGl�������X*����!e�u���׋X�5��2�[�q���}�^�BA��E�^�mY�ೀѭ���ˁT�&#�4c��Ul�	�Q��:I_D]�Ӂ�������T��3����<�:gT0A�P;�,1=�!7�h&܁nD�EZ��
�̇ȗE���E=[�<�>mg.��P?����1���v�W���0�t�/��vh�Bga��^$��\��F�7K��3������Q5V�u��z��U�_�����$������_fxIs�C�Y��ҝ��:K6�&v)����x�V�� �7�?+-��3$g�b����B�ϑ%n�RK��"q=0��Z[��3VH���Ѕ����2��R�]{��m��4�]�Oz�&�Z�n[s�QdX�,�_7��p��{���2�S�4�j����fƢȏ��J�XC����qJ1:���<�	ֱ�<\�r���Bz���y��Ҁ�F�T��6�] ڿ�z,0�幇\�B��c� �����+�V�����
,��U�N�H�`k}� j'����k{�1u��!�б�Y,%).|�5�<���Ч�':�$��?A�H���<�ÒIwM�:I2���}�w��IpT�զ`p���ȲZH����ZCB�'����.��v��@�3� gx���.��v]\<k2KfK���Q���0�R�bR�U��V��9~�T�&ƔCgj�/������eW��|���4_Ө�,!��� �KL.7Zſ�t��r3\@�nG��(�����	�X���V�	2�p������~�i3 ��M��%�#|���	����3n$�0�j Y\��-9�"��»��x��6����6`C/�����B���ws$�U��Q���CS�,�5H�C<q@p��-�.�I�R!��#H9 ��[�ȃ���?���A�q�A@���;�=k�g��
����M~R4!E29t-�j�t���Vu�.��J�j����m������JJ��C�*�ߑJ��#�Z�JPؠ�������g{k��}� f`z���t��葡]�ž��3��G���b�7���^�Q&�l��mA� K��H�k��ύ��B�����;���|�G���u�᝝ǰ��{y�/�$i����%����A� � ���vl*b���V���T+\�w�Hj'E�O�D�j
������Q\1 ���1�Pu��W6�pZY��b�5�. ���TۗL^��.�,5�л�5pU(��^B�J�{�����\3���P�H&��f�����%� / 9�(*��s�3�^p����9;tu��om�,Ѝ,{[��Y��͋�_�ڠv1	#&P{M��Ō�.A�#3�{ �v�Q������,*#��WP�	���I��[Jz����3�4���'W���2h� E�����jz)a �J�`�6��*YB#:rM\�Y�F��%���� M���+b���V����\��KȊ*L�X����S;��\U�^���"t�mX���F�{>�y7��f�U�6}���L��҄ ��J���r�ٳfN����,-R9+^��i3�N��8��ѱ���ś��O�u�~�u`��"�z,]�DV
�z����o3��]����ǠȪV�5�����i�_S�s�����hs��o�e�څ���@E���E?ͽ�9v$�����dGiA8����S��zС�� ��r�s��6+�[-9�k6���zZ9	��,���u�0���X�2���%5������������d׾�6k݇�P�8�Q� ͏_8�3^j"ѫ�QO��x�\1N<�������n���&#lµԐHKB�iڌ�8Q�q&!=}���=X�U�G�Y(���7h~hB4Z�үRY�!��`�S�4�Q�hD>�r�x
���+��.as<�>�O0��=�"��bu��:��Tu�m��=��a���@Wa=�j���h�s�3��)���I��_���c�\��{5��B�l0'�L�\	���.�=Yc��r�	�5Ьm�J��<�-�y������ǖ�;�Ӌx)Yp2���X���rK�#�"��U��*����҃��-y��%Ns+F��T���_'x,�]?P835����>~h��*��/l𾺌?�����_1:W���L�Q�*��M��H��D�9�����;@�dQ�)ȝ��Hn��J���z�| ��1}�W�^������w���C��yH����0�{c�P�@�]U�/�ijH���?T�V���
�:��]�~��:��ay8��:�Zݾc���&�1�{*�iB�ćӳtOo{x�ix�(�G\�套�K5��˄Pw��K�B��4g.pKS����˻�i����2����g��[��-�~&^c�[�����Z@O�4*�%#ݩJƱu��Z�&�Ͽ�:|����nR��q�w��E���d�q�D.x�i�O�KI���\cg灛�+�a@sQ'̳�R�9��\Br2���o摟�U���K�x���	л?��k`����פk�p�hV�OK�#h�*�5���2��!��I������%Zh��$����[���J�b�Y�l��+e�9ڗ�PhP�<�h�eh����=\aҏ��9���%b��|��Ś^I"��]��0�o#p瓘���%�J`����4�E��ٴ���q�+ڪ/LjЄt�j�&��I6V|�T5tA�q�����tۖ��l��Λ���:��K� sD8�s.�/,n\]��Q�Z,�������	L<H�ZFj�g������X�!/����N��Ď��
�r�f��  V4�=,#A���,��8�)�
�dj�U���>����&b���K>4�u��fnaɁ>�0�7s����n9t�4^p?޽�gà�3�ڜ���5_�ͯ�,��H&
P_��zbA�ܛ�~���t�D�W��KJ��	�oƖ[�Dò�y��o�i�v�>(j_)��03���ݠ�0�"�3���F�Ɂ"@�C�(�Q���*Jh��ůt�\q�� �l�����3���w�;�~�KZ:�.����$x�D��ތ������N���q�0_�Lu���x��ӈ+��sП�BD=I�F������W����X�0�`P��G�(�[�rp��7�3.n�	������G�8|�vD઀D"��(���Z���d����d<A�<�:����V:����8�MN�bk�x�(�U�B��{�}�m��H�?#z�,����gD��?��Z%a�? MP�Np � ,��J7�H0�,<t��bv�fdn}��0�@%���u�-�z��H]�"r}x���"��S՗�f��~�	5gMV��!�-�3�����r;U�2�Ü�=�fH?-W&�5��Ea��?����;��!�$��Y{>����)t��D ��K�'�S� ������2'���(Sˀ)iMΤ��잔��t��+�[\W�_�Xcʯ� �=ߋs�,&�X��tt���M�� r��|l9�q��[�������O/�	�&]���d�����]|˦�vBYQ��2O�O)�1�]�=�S>�\��lw�Z����&y��M�~��:�EHj��C����Ə�)ߌ��p�l�5��b�qQK��u�ؠ�����Cs&{���ڭV�w?�B$��쉱w�-i�.>P��(��F}TG�Xsƛ�X��h$P<��hA���Aܢ���P8�0ę�r�y��I�x�T"�vZ+����k`�倌���+�G�;U�_��������)3���ބx�)�lYЖ"&� k�*eI��O�;27�� ]1��u������
���w�bA�#K}�y����#B��q�out=c8�@��v�m����u� ����Pi2s27Zܮuz��;"����LyN����S�h��24��.��p��h!�QQ�l�Fo�����=Ƌ� ͻ��y�Q�;܀�>������i��������n��on�l%_Q߳����XW���_���J��,�T�2�^���j/��.��!�b7NV��$[�dX�,��$���a��At�lH�FkrEq�t�$_�g��"@~Q�_�.�>%0�-4�]��&;�������t���~%$�?m�n��Ԭz�Gk]�{�AFF/��$���f�3mm?c�I�N#þ����6ŁÁ$��5z�N�A�}rX4�����'[ݐ��5/��G��kz =�.g���I��뙹q,4l�!Mv�����|�?��	"Gg�a�"�BD�I�Zϧ��_�-?[a=�c?7Y��MʂT���W~�g�H��E ���<�V(�$J6u�˃$݊�h;g�xAȱ@��x/��g��6���Hm���b�dV���ذj&}|��ۥV�܅���٤�D�lj܅;��;��Ը�n�W�T�Ù�fGeNH��QzJ�q0q�^���ܓ�9+��W���(���$"��1�0��(;���7~�*����0��1�8$�����n;BĂY�.���YPR�0w��ʂ��6�v��	,�/�H�[�a^��#Ni?e�`���:Tp�e;�Y]�P����08�lVskZ3LvT�tj�.�E�f�qiE_%ZW�\YVAy�����(�O�K��ϝC*�m��-��oc՗ڃ�&:�K��!�|D>h��`rX�n��T�oLp+|�5]�I]ܜR��;��`t�ǚ��~��S�������ʞ����k;)���g:�޸��o�dw��X 
XpL���Zf.-l� �ƍ_
��i7w��y��/l���}��Юv��v!����dH"��'}׵ч�R�5��rf���Y�I
���{���"��|܃��k��Q�[)?�<yp�~�ω�1!lm�D��*)��q���)�,�/��a���'� xL�E�+Wl��x�!$	��Ϗx7��WS�����x��%����'�埊_�r�1H,J���iV���ݑ0����{SX�5� �./x�/pp��+���*�US�Ϗ��L�;�I��/T�R�2J��,7[��=\b%y
B���y�t~�I�ٽ��
������:i'
ÿ�l�Ձ�̓����@9{��{������&:�a�:���KW5�^Gs$�ǈ��)�0����{+�e����Q���Z����29z�� F�(T�u�"��֫�O���,{�Sݼϴ`���S�rư%C���}���Nk�0��>�V�,�W�+��'B{r��G!0��'A���j�@�No�!�ã+~�О�8f��y��A�f��i�x]�7P�������*�͖:�l_�\�*��Q�d�H�Q5z�T��=a �b��|s��z�+
��웘X@�n�8X&���_����Y��q]��%�	���i:����A��%��؜�i|�*y��5SM��L�Ε�5;��pI�q�Y�	!s���ޅ�H�7��m�_�e�?n|�"k���0EM��j�����_%��f�E&ý@��{��Ai�"��6 -Jm�AK������bT�ȟ�Л��A�C�#嚎:l���nK%�e�ó� �m�ԑ$�Y�AM; �D�2V����<���}.�vZ��W�cR�s�粟�5��<�W��!��;����.��~_�=�1��JX吒]F�f1U0]/ys������d�%���>���Q]`0�q<
�=��q�4G��c��yK��{2�]��>�MR��G}��s�3G����Y� ��/�Ծc1�Uo�S��n�Ǥѻ�G��*�ѰJ�먖���2��Ť k48������3�})=>_A~��¯FEb���Mڪ"����X��]���I}EHJs��%��,'��'�����3�g3���T
L�V�a4��+��س�cz��@,�j�[T�'�f!�J^�ټ E�;��a*�OA�t3\��I�z��ҫ#*>C�������%r�ǝ�kg����[���d8�x5p
�����s�xveh��ww�a �@��}�;7�=�L��u)/��u�*��(H�U�Q��Z�%�%��׮A����Yt�{�H��<�/:�9���&:�u��~ݟx|�y�}�u�4h<_��w�:�ѿ�L�c��4L���o%x�Ն���4
>o�N\�x �Dwau�\���T�@pe�nYh�yA�*�%����}o�zT��Z4�_~��ξ�$������S��Ǿ;��5iu<_B��mheW�T�WAz��-ZD#BT��
�=e����/'��ܖ�ϴ�e�~ܽ䒋PI&��l��>�Z�9��&Ł)Uo�ڪ�F�冘�h�ae�/������M�-+嘙@F�q#蒻,�Ll����kg�|~��h�7�/i(�}�����3���nf{0c�k��N�uS���2X�b�'�����[�%k���]������7��C���h^���"f��l�Qh�u��g����
��
LE���6��Ŀ�0�E;R�.�;��Òԕˤ����ZW5B,��2+�1o�3a��<z[�cc�l$j�o4]B��n�j@7}V����+.�$�[����Z��}�h��Icp��*7IdC@����\3_*ӿ�
zE��t?��<�=���+����{	�p��Z0镜E�s�|�i�G��T�@�/Y��T�C
o3����F��2��n*�P��n�O��ޛ��Xүv;x�,p��V8dB��p�[bu�M�����ΑB�⦥HϠ1���}�-;s.�雂���0=}�_
͛�f�?���p�5k�13��T��Ҭ�\O�,(ݸD�>vF9�"�N�K��H#"�}J�*l��O��ׄ��(�w*��͡��j]Td���udc�p3������j�:QT�ǳ?r�u��8�'���z�#����ͻg�B�0D����R���TE����JD��0�V��M�}��%�0Y�Ǉ���e��E�Otl9&i��'�}!T�dY��!�Ug��ig�+ ����)t��b3%��*�G�Ce��M���K�c\���FI��z�s�&du`���V�)ˈ�)y;��~��S���[#��|YcΆ�ƩI��S�Qy36��rW2�777	����:���e��_.��`��A�w^W%\"��Pz0�wP�p*X�˪�i��7��>�9���ħ���ώ��{:z�龸�ӓ����M���bC��I?RiX�k�E����s�}��U�#e)@7�7Y�d*��"���C��A�?/u�c��僠��2'Fb�wo�ہ'�u�c��C�E���_VUD�HT�#�4�w����1fO5[��O^��.$;����L�G$���/��֩ӁJ�H�כ�Ѱ� l���X���]�D$E�a��s��)�IV&_�"�l�=� ��w�hv��]�X��!YQ�(�C�qй���R�Ѷ�1��z�0��)�|�UW�[ y��T�p�hݍ���� ���*�& Xg8��D�s�<��p�W�}��8�y�������Z��IW>��\��=����t�GjK���©;@ońq��g+���^霼��,����:I����ai~R$�{�C���eK�<��t���h��F�c���ob<pc����I�Z�� �t�:,�Y-o-Ѐ弹Xa69w "U�!��g
9��?�0� ����(ǌ������.�_²��d0��զ�Q�	�n�2�����b��i�<�H�e�4�f3N)��	����������'��t�"ݼg�5��Lon����ڛ�(�Y�i�b�W�x��U��P.�/r�,��Z��k�u�C�d���'#�_��2"�޿D�3���oQ+VP�����K�T�vk'��Y���Ԇ=ݶ%�b乑(��z\.֘��+�y�q~@$h|�G�ޖ�]�f��Jqq�:��G��!���ƃ���V#�.r؄ܗ$e`�Hv�]����~e.7����]C"�&���eM�*@����H�K9�-���j�����U�x.��2h����؄�K��?I�B��ď�u�Y:�l��;�<��\R*'A?��:mS��'�vab��vi��[>J��i߂�䒋��Ȍ�$�~�L:D��W'h5�h��
���[����W�q,�>Bi��Ur���i_ԖM���������+��a�9� G������h�*�! `�=k�py�偕�N%}�mO�^WPg����d��:f�v�b�P�ǡI�z��a5�0�1��,K�ag,٤�t}ڠ$��28�\��T�u�F ԼX�?����<���OPO,
6��M)}��kC����I�U\R�N�����:Q���q�U�4�Y��طjg_���>��{������&�;�le�B��������8hZNF�c4���#R� ;��)L���2_�J<�B-4��E;d�����h�mX؄����%us�4�����i��Q�69� ;\a��3z�S���6̸�-��|���d�����#��i�?j�0��[ 9�j�	���;�z� �0��������+��L��f�g)�&�G�
K��?3�p��F�1&�Ds�+�FS
>�|ӫ)���c��>�5۔�/_��"��<qÙޓ�+F��&@��M����\��h�K�P�0������.�#Li����6I@⥉Og`3�[IS�ؿp���1U\%Ʈ�{��5�"ZR��y����@x{n¯�حsJ�;���(ǽ]�[
�Vx;�S�,�������j9�Dt�x#�C�sW�Bu�����P8�})�c�1ꀰp��8s�����1뤓0��)�����׋e� �%���|ʵb�V�������Ŋ^��-��Ċ��/�0�^k�$�f���s K�(#����&���;�N���>�C��~S��Ȏq~f��;�Z�}"�Ur�4h����k�&=<�kk�hK��=��_�}�^*�$m�f��~�Ȅ�J����y�5ئ�"ٳY͆�G����p���#i��7a���6�j�uJ�rj��,�3V+ $Mm�%�O��S�Z��}bduf�E��06rԎ ��8I;�p�Χ��c0M����a�?s�j�0�:�-'�7#����<r�f+���lp$Zڿ��C[qܴ�]7'�(���3bcm�ǝ>$S]#�+(�_�)g�<�I��Qހ
�n�֗.?Y7-���!�&�NU,v��].��)���7b�m��	h�b����L��G��T�F$�W���9-Y45[UbpQ������i���կ�����YH0_].̑s���ְV��吮6��R9���I���B+MT�5�O�e
E�R~��TN q�9��mb�aF�U��|��'��T�'���<�`��"�ꓐ�6��]����;^d�8�D�̍L��`�M���P51L�|+'���m^Vu������';r�����:�i�.��#���S	Zօ��&�4�f���C���Y=�p�;�{^fG�	�^Z*�P7��^t���t�g��q��w�7nT�
M\��4�E
޴Wܕc�x���X�0vK�va(Ӆk`	�o��WWsEP��������X�G�y;}����g�#�}SyOI�ꖜ@(bc�( �|}�o��mSI��'Js Δ��CD������w�C�q��Fx��w��EЭ^r/�X��j�G��&í�#~Hqaɋ,�C�&�L\*����6h\�����=��i>���>��5�� �}�,�ی��G��</tb������ڞd�u&��ާ�]�ʛo[H�l�/5<'0GU��:���9��߫����e�� ����eECyԡ��(+!t��^�����>����T|�"�?�ZNJG�'��Go�t��;q���)!d�^F��I]A���)�EسW��@��]��1��DΕ�_B�A\�βZ6�µ�������dxoP����^��)Nɧ�8ǲR�)������NƐ'�Aom�ic�}S�K5U�14�Ň%����l*W�_��~�ܷ�a��f"3)��(�� �������^ ��mT���p4�d����K��8s��-�}��I��EU��؂�M��D�Z��1^h/N�=�q�9)���p�}+MscXQZJ�f���x�Q�c�2�$G�W����`���k6�9���,���O�����������%�O4����}�u����P���l&9�_(�5�[M��X���Na�z����_������2��� hUU�5M��+@H�&[ z?���{j�(���$�B�F�8����@.okiߙ�j $�{��N6���)�.�W?@�!q�>bG�+\��\���?B)NW{߭"x����~6�ڤm���2Oy���T�Ro��w���,9D�����t�w�8m�ɾ��̆��R���E1=��A�J�������SV�Q5y6�$��;�F��T��Y�7��:��CA&Z�@�O�kU�J��_���_0�d}#;�R�Qj̘*�����nFIg�Q�̶��+7'C3�|{���8��'�[������^����Ƭ&�y�� 9��h|��:R���My��ŗ��c��Z�|�^�C���|��iv왖ue�(�:�ns0��[�u��]$f����QwK?��rN�'D{\ꏽ��|,�<4;�.���H&N����b`��?x���^X֒�
�.�ɝ1�j�y���p�4�O>��Gѱ*��Z~߈ 	��U�IN���ƩZ	�G�UE���I%�Yt�uXu��'�H��Lz��t��&�J"����a�B��;���7���yW��J���3������>q~A��y}�����oV���@-W�Y��z���
�A�m�ᎈ
֔� >�( �?y"�Z��R_U��w�0��J��|0bʑ�;��qIH|j¡R$�P[��g�QV�@V�=�
/�ޫ�B#z4]ع 6.�4y�89�P��*8��K�w�2�;�)�n��u\���2+���p���?8J�l�kDiF󁠿�lV��i5����D�z�M�"�I�2�![� ï��U��"���yC=��N��e�v�t��N�W����O�oS\�Oa�nQm��!v����5f���5��e�ώ����&��I��%�H�'#0�;"}�č�� �ge&�NkO��l�セ��^�G�狖��<9���U�0����P�}�@Y�7�6a~bp�Nc�ܯΊd��n��7�|&�y�F��&';�3�'1<7�*�!c�+Ѓ���H� m� �#vE�����=�zVV��:R�9B�h��X��ꘐ���'՚��)�
L��O�Xy�}۵�dH'G�;F��b�ϗw������<�Q�q;�K��W�_k6~�[���z�a��o�g u�S��� ��9q��.�R7i����!�r�r j�~�s<��4|�SF�����4:Ӵ���|u��d�E-�o��;Ѝ��nq�qOTPXEj���6x�C�ŏ;��C��G0�<jm���z��z�oM�Fd�ΐ��n�b�ux�U���fΕR��T{8��p��!c)��w��.5����j��"z��p��S|o��̤���wi�.b}�9Y��u��`���u����фD;Zu7��"�4S=�y�`��~�u��Y�D�Ex3�c��(qa�+�ih�V<�j���h��7�/_��)���d)��|�S8��߆Eǉ���S���	�g�R�\zN���h�L;�
9u��%�߰�y̧Kx�������ܷ�ȷ*�%��w�&��F��wOҥ+�y���Ƶ��s�@yMH�N�q��ǭz1���2�̿�UO��K��B$�"y�J����sc���Յ���9L�����Y����M0��8m^�+Þ�X.�����BƢ��
��\�0��i#ޥ��g��d-��/F����Lb;#O"H���Ʃ|:��G�Vd��F6��/���Z�/k̼��/���ex�8��@��D�'�Q�
���mc�����5�X�1��{+W�F)�zi�q�Cfʡ"��4'�?}.:F4��4��S��� Y_e>Y�}�2�f��e�u�%�ꛦak1������G~���#u���g��$\Ǟ2��~����K��	w� �K���M���w��6Hr�©���}�r���"�s�Kd_*iy,7�Y���DZH}*�/4�᳭�+��
"���z?8�1�&ul���~2�g�ah�Ɵ ��[��}`豐[�lT"�`K#���i�@�Vz�O�v+T7�E�ʔ]�K�0�翕R�DZ�K%��61)�����=��6G:��[J�[#��NB��3�;v�LT��A�NM���Z96����������~��-uIy���Wʒ�@��+KT]i�8�ڍ��a�0�G�w�PZ&9L�٢���P�)�]R����g�C<���ӱ�W\�=����į�1I���Q�uFv0]O�O��/�OƊ#��t�M��E4^X��+j�ݼ"�s{��h��������7��&��b�w�%�����9�ۆz�դ�."��/��R/l07��z+�N5C�j��u�l$,B�
AT�Jˑ|忌1/%�LWh-�뚝��-��\Y���^�'�"2#ʟbޓ�Yݠ6�V'ۅ�e�u��o\Uh���u��o3uZ���߅`�\h�X�>�4P;��neg[o�ϰR�m+�T�l&��{�b� 8��2�>j3�] Y�Rif��}k��9\^<� ��
(�t-\A-v}k�	��/��8���p�C�6\-�~)�ndP, ��f_�
:��(/�OΆ���9�`��9;b8{t���v�X�����?|E5 2�kb�]!CRȕ"�wh�� q�sb����J{��ôx�t�>_Ċy�]���J��גcl_��NS��\&�v#�v��;���"��7'm64��S2zE׏��9E���g���.21�e��D��^���qkm��6���D�` Lvzf�9T����/���7��P<�*��u�>��NG)LW^w�+�0��	���4Z7OMʶ��<ױe��UR��Y״�g�c�����w"�LH8EVS'�'ϔ8q�X�<'��,���~��}�	~-llo�4�j�*�2S)��#��~SA;��-$v�
s��w���&�*�k�iɂ�C�̈F�&8ȫ,^��9���@�ûw���R��.g9Nv}~~��R�AY"��[c�	�f�������ڈ����a��ڧ	��M~��*�awV?�AT�oX�ix7qƕ�&��X��O��=���ׄyJ�����}��W�9?�ӡ�A�vrM��D����*RBM�o���\9�1)C3f]=0W�:�¶t|�y7�N�ީ�s�W	�خx��r)cU~|��(6�Ȫl�LiT ��n3��KFy�����"�4��m")�W7�l>�*��2v���Ǉŉ=9I���3oK �
�Gr�Cv8�A���-�,C�a�W��4 ���g�sb��+��!����|]K^"�P�����X�\O�}��O��������vk�������G8t�#�*S1�O��e,@˱I5��J�I����!2�J�(��}r���G��ю� 0^���C���.���5�bb�*x>i��o	����z�H���8�Č�O;�e	�'�������V��཈��eZ�y1�w��E1��*���=a�Y}M��ޖs�~�@F~��XV
f�[�On/���u��f���33�Z��7�2����������8���\Ѧ��V�8�w�H�՚߭�qm��T)�ު��x`�>3K���5�a��}{7�u7��[�o�@S���d(��K*1��_Hsv�汤�$mws�G-�(�1������RH��5�B�1�S�B��)��ݕ[W5Z�ܕ��V)����ANXtPYr̛9����@Qh��e�I52A�S�4b��y~�#�.`��_m���
b5�F��Xo��Oe�R�F���a5���5PWs�����&��pܪ5���O��CH�f�+N�=��y�OԿ2[�Z5���C�k7a��v5�WƸ.�ցeh?��M�^*�6�?����o���Q��WS�]����}$}�<�^����j�:�0ˬ���Jr��0/m
(2�٤�J���)_�fS�<�ܸ�YA���}�U�L=��D?�.�z^%���]���� ��n7ES�����w�_^�)��c��W.�O�z�;��p��,_��'H��ܽFY㨞���r��z"�e�R� ĹC���І�7��D�Ov�F�tO�oD��N"�f@٨�0,�ۓ�&�|�=g�m���&K���1��Y�ff�Ǳ�զ7B0!����%��P�&(��ғ���@Ywk�$V����r�F�?!��D�<m&,Ù�Sr����q�pG�*�߸J�6\��>�y�&^����<�k4ô�۩��O�٧��Ձ����{֑�f2w\ͬB���S�u�b"�b��=J�]n���0bI�ɽm4�:��߁���~Uj\�Y�0���`F�I�'�q�R��(�W{ڸ�s��ab��	^[+�$�х�dFC��🎕��A���0Y�4kzYm/3FE��������\lLڬ�0g��I���@��D>��e�/��]�@,�[Ő{}�/�g����c�z���*4�P��Xحdw��D�#�H*b��p����&\(ſ� ��2V�jG��u��٤�Ɛ^�a�X�s@�>Dx��+�r�M�*����ěG=7M5�@Ha��(7�qm��2��nY�M�}n���,NRt?6;0��?��̠���������B�����٬D��h�D��:����{|�#���ę�R������au���+{S�Q��y7]�k�^�5*�+�_J���n�)�V����S�Z6&��[�&]���!�\�G&1�;��@��d�F!Xh��o�#�Vv���˄Q�H�[���y�tzo��'�;�I�G��!Y5#5�
�WI�a���*#��k�B��Sie�jM����I"�d.��?���;�8�Vh��n�FR�ֺ�+&�p����V;�oa<�r�^~�bB��'���f����%����c�U 9���ȝ)A����ģ/%|�������z%�\a������2I/L�#�(>z9c^T3(�y}H,�����;�j��Р)��������ab~r�+O�����ҼF��}��1��
R{�g�Y�k�M�Z�)eQ@RT�s�N����	&�֠>b��/������Cj�1���:<��f�Bd��I��4��?4yoY;Ӯ�3hp�h1vq��7�G����j��� ��b`�H��\;�(m�]��f.Y<��xS)�-�	��G��5\	��Nn�G���+|���$O� ۢ�Ѱ�D����I~U�?,x�U��h�� ��	��3�\�Lz��Q�)�K�_� i5��vI���`wjI�� 7��s95��}��2,����p�!HT(��z-N�VIrl��ޕּtɣA�,E`FD�7W%�@��3#���P����\�>���+��5�9.m�������8��Q�zRJ ����J�P"���S���ƚ�Ɩ����[N�QII�� %�u�4,�GO\$V?�RJ�Vh����� O��	o��WE}�l�ۤ�EG����h�!�����WX4�h� �C8ɍG��E��̫eK�|z�CJ�����Ahe�Pu
n�P�����ҡ����%{��N���RZW�c]����t���~�P�9�!�)Ov	��ʫ�Tr��{�x���mG��=��4�%ɤ�	��;��s������'0!�R��� �Y�QH�x���wm)��-�y��\&j��[���%�J���>̎g�]K:9�x�O47�v��|�@�o�\mCg��/�r��_�R�^|�1���������k>���^ �o1R�!ڒ{8v~��`}��gx��fK$�C��t�}��ݷMqۊ�.DZ�=���,C��[�ўζ�mJ�O�o�4�`",�یL�ӆ��.�\��t*�ml���L���6 ��/�
]�tR�R�����'�4Q]�C���P�>gW[�^^��+s������K�3kmsM&�ha��[�L��T�Oܱ�Y_���ݫH��@�@V�.�B~^�;1���}��?6����D����ϵ�pi8Kn�q�" ��~��[Ћ@D�7zP�X��?գ��0�!)g䰫��-�š��6@9P�C_����y��)��ކ���t|��9�Q�װ]gҘ�e�:I=J$���ѫT�i����X L�{x@̓��Y�xe���>������/��X�)<�ܞY6����ٌ�[�G�&�d����A:-�=X�e�:Ȥ����{�����[�z{���U�X�X�nL<B�먭��x�m�r>eR���_���|��'j��ZɪXrN�񡄿�oM�A��/RƂ�e�h�⍳g�Y1V�	3�g&��E
Uڪ3����݈Q}��W��ƘnBB��$�'�9�ho
ǝ�,)}haĈ)u����:�ȅVˢ9�B�Z�%�:��T�~�������T�#��;�""��w�����L{�b��F�Cz��/�m���� �jB#��I�d"�a��X�F4���Ck�h2/���7�qVm�ӽ�����r4R[c��:�;)tj�*Qp�kO�(��=�{~4��
O�훺Y��V�R�3�[1�=����.f��BY<9�RNf�XVR��2����Α�4�>��)�Qv� ���𢧱�f8�x΂��aM���ݼf��$ㅬ+��e�%�ht,?�mrj��ڜ������~���'��C`�j�>���Uzu��J=@�й����$��0��d4:�1��ۋ�A�<�(L]��2�C��o��|�4������.���fנ��]/�b�ښϋ1��_�s˞	*<U�B�+�p���"���h�⸁6�<f����}��+�[�ړ0��E26>l�l��a��
L�c��gd���`��#w1��)M'���0���t��(���b'�2-e-�_[�b���VL(L:	$ࣲ�� �Ⱥ���H;H�Ԟ6�{� v���B����ch���hN�s2��g��,(`�Ɏa�9��ԷEb7N����}ĨeP��+�]�⢵�][ma̱�>�}Ar��)m������8��)T�T�B�����ܓ�A��yC�^x"���eg�'ܳ�І��?I�qZ�ހz�1vX/WZk3��5��D=�ob/�	^;qKx׳�Ќ��q����F���_�{� YcQ���d�b�)�:�1*rj*��Y	��z��+�-4��&=H&�g��ou��qj��D3� �|Ch��Z�}���e�a/�E�3s�>���i�gc�r*��]O�4�ජ�楜���_��ݕ�%8@?�~"��r�Վ������]&��EO_ܼ�T�Y���&rx�̶��v�.��I�fN��m|5-��"^啁D�a�6w�{m���,W�8��e�������-O�� 9��+�,�̹j�2N|�L҆���G��p��r�YF�j�蔜-WӮ2�&zX�c�j볂NdS���Q!�������g3GQT)GΔ5?��6�h�s���)�[K �M^;M��'s�K�bQ���O�l���t�aR��hB�J^�bdg�=6��]�����w��?���3�2E;Jb���\L����؋���a�ը�ّ��Q�P����E�ˢ��y������
�� xU��X94����C�k�P��ϻ��A�F.i��#�����-��
���"����G�!#���˼�CpSo�&�{Zޓ�O(k�ۊ��4��/�Dѻ���,PZi���t�.BЪ�.���*:h&��1n��R�9Y8����E�X�#j�L��x{O��Fj�����O�6��� ���1P�2�\?7Lc��!s���6��$�v6�Q�4ڬ��l{��N��d���m���k�e��V��z�f�(ࡵ;W���~��Y ��v;l�y��tP��3�[�#��EN�\���C�S�g�_�?��Nۈ �dJ�(�Ǌ�����G��%{p��+y�߾�m���1���t@��DbN�{��ϛ[��
M]�A�士��ڏ�!��r���8�+���ğ�#���e��MY	(�O��*������+�0,�p޾�K�>����2�)��e��f~
�0�1D�,�V �*��&����|���v�r����8}����7&�
�}���-��X��Z�1��g��$��;	]Zd�1 ���ON�C�!��.W���H���O�:�]�	�_�o����6w}��VG4:.��|��42h���9yaF��
��ܬ�y��$��l3 ,�1X��MC�ۅ����/Q:b�8�/(M�����|�gN$���
eþ����ǊYѸ��r?��O.�U:�VV�?�N��_E_�����V���ίv�|,�HM�5%T�,���� B3P��C!t�Ly��'ް�c�h/q}u-x�]�9�y����J��$VFǲ�~�jJ�t�Ry�^#�}�z����/_�魏ͭ{wF���b0���n�V���:_t��ʬ܄�N�x&]2�,3�f��и�j�3�F��ԕ�~ڢ���WA%�b�Z/ܪp'�Ln�O�Aߝ���{�`�N�i���M[�^&wK���R�"/����g�>@����,t��˃��O9�V���������q�8_�r�'��#f�N���kd����Y�txgM��߁쮣G����MF���NjyM���^�3��֏�G� �l����@W �`�T�Y,�M�5���pm�Ǥe]iF�7�äE�e
؝~���ތ򉯛��@���|A������Rz#������F��g��ɥ{z����>���O9��JT���k����EfV;�M��)Aߠea�Lu�z��901�$*j��s��؞8����'����C
O6�vS�Z��S�y^���J�.���0��c��cmߡF�C��F�R�E�Cs˅�6��a~� �z�^5(aЍV��z3jm<J\s�m�$�>F�VfH�Ϩ-]|}#ջ��I�N.s���t׹��[zO�0�J���=w�������W�WFt�*�m�����yo�U���j?�O�W���.W00ꇞO��H�Q�&0��N@F���=���qvv�L᫙�[]�2�=M�)�mN��@A����aH���zf���M��=��IK+ʊ3$}��D��ߏ�&:xN�Ŵ�F��Ɩ�@!ִ4^-��˒��G������o�l}�fp�&h��ؠ��}Jc5gΤ$Zip�';��[����G��Μ�&�Ƈ�%k��Q=��^�<�-��.qy`:h�vv��	�<c�lғ%��)˴�\h(j�֛o��Y�G���o<D�qh�<[�W�����"�<YQ����%��,eݡ�(�E^�B��p��'�q�0Okގ��ZMԑE��ٓI�c��5�����i��	��U<"��}�Rj %��2�n7�R%h ���rV��=ݿ���0��$z�z7��~�L�җk���h`�����_���e$���S�
4w	�j�8�U<uA��cj�y��1�BT)g��b�������Y�c��%��D���ސ�����ҩGi����m�Ώ;CS�^��&��\�5)�U25wsT�&���B�?ͲI*l���[{��l3��5�/uk���ȝg
���7���ɺ����s/[�Y�\���8�Y��iC����6?{��y�]�poW�����^h��sR�mlƪ��A����eHL��E�S���X$5p��G����,E��N�#��b�(��^2s �5!��}��Gg������u�r=~�A|��Ey�%� E/=���o�h��^t|��#Aue��ʶ��&r�@��7�$ٵ���:�?�"f��h�������Gw�`�6�`P|"�H��0�� �ac�C����h@�؃Tۍ��2���_s*�[��(��y�
�a��VK�~�X�NU����Ta�Ti6<�J~��e�qubA��c�m�g���tc�T���O^j��婻�t�6���H��y��!3%�ha����K�xE�~���[���i����j��EX-��_Q��$cI��z�\/�����.���'��{�Z10jS�u�i�\�E����ޞ�B]h�H�	M��EF�2�Cc�Ŵ��0�T�XW�b5�滺����2q��b��4,%�E����}R�DE��������}�����	�.�Vj�̜��l��f`�ٹ�6��`�����*N{<�dGS��>�&��87��e꽸��T�Ku
?��7����вN����7{�-�w�o����h�*ʨ��+�|�c&
�m!����,;|ݾf��h�y6f�z������G�DR��bb�˶�gc��4�n��bh�<�� YخSad���`0��eF:�J�ݨi��42E6>��JMĒhM�����9���!��Nd�k��2������-G��oW��J�]��cO�C����y��JG�ˆ���QtEg�p]�T��w}�<:��r�g�P� ����QL�z��[9��6�&Ͽ4�2#�"X�±���22����Q����!h�Y!��&�{�[�C̈�_h�d��K�҆���es��)H�����5�D���oa���Y�BF7���^��uz7e\m��LR����r�k�B�I�h�����(�=#�t�`���6�gC������o��pV'f��L��܍��"oWm]P3�H[гK~O�la9���6SGdI�1�BdY\��ٴs�%�"�1�J�U�{�%�T�
}^�9�ȹ����iK������LF�?����e�dJ�Ү��\B����9�NP&7�~��,9�E��U�%�].���W̯6Qp��Fb^5��\��y���r����lg�%���HՌC�;_�@K��Z�d�z)��"O�|�>�R3̓�N��d����l��)Xo0�!6�S��\L4�k1u	�^`�<�?o��惡A\���ǎ���4��{A ��;ק�=[Z1�l�]�]���il񅲼�:�F=��߆�Y�,��=���+� 2�7�ZL�V%xvLWBJZ����Q�͢��F�33LƎџ;�Lz���I/���ħ	ʊ�c8Z���:�<��m�cV�r��r��u2�Te �Rdw�qu�}�R8�x��iR��̃$�K��.T�ȷGU��^��(�|�=�)9���+3��4���.ٰ�	���7D��w�0 ͼM�Uk�=�A�em�w�M�����F���A򛼡�F��;x	wx��z�R�|�J�;���9�8�r�J=�1�-s�L��9���?���p8
��������K�xLj塸�8�u)�����A��>��*yd�0B�6,��� �g�+�%�E39�_銵�=C��V0d8�Ƅ$���<��%�C�Y_�!.D�|D��������|{�����*/ծ?����H��'0����fF�TPOx����6�UA�7:=�D�숕.(�������%�뷫�}��+o ��e�f��ڃ>di]KI
�឵��i�[ɻ��9��U����'�����u�Vo�R6?����ߝ�ɸ<Wnȏ�]k(�Rh@9q��h�����c  ��u��`�Yw1`AJ�<<���tj�mvh�C}�h�5mC�fJFO�[��%͗A�^@䭣9f*�?y4��	|3�i�%�Y[����.Qc0*N~����!j�T�o�E[Op�z��bS��Ƽn����g|Xm�a����ר:���ܧ�| ]����
X�I[�co��c+T�PԺ(ЛB$��������h�kH�}�a�jt��G�E�K͊�4��8�x���{���hS�|grf���@.%��Uy�C��m����BIң&+����M����w+֭��{襟���qu9H7���s5k|������Й��+e����i�;���%'�Z�!�t< �_���B�"�}�����`�Nio�M�.)�^z��=N�W���%�Q��oe�R\������L�E_(��*�ě@� �����	U�#��r�����,�$ȣb��C1���n��jg��:!��6HB��I=�.����tPv�8)P��X�~&���Fĝ�u�Yݐ���E�B�b-���.wY�L:z�ĵ��u�U���	�,*���@�@�[�B@�VC>'v3Xw��������n+3��52ˋ|ȝ鿾�$�,�Ο��v�s&��t�O� �Hリ�E�B��9�u!���N���4iB���:���������1r���PZ�1��g'��ߗ���J�#�ec�4ǰ�A�|�Dyh����d	��$�������^�|�U~V�[���l'��4�����-c1f�4W����'���r����8WBV��(��x���o�{.<{�gقm��@f��H\&��յ$�|��d�E~�뙑U���Y۴�a��M�Ԯ�@
H���� sk���P�+`�]��H��hb��A������⁻3�mE��T��gh�W�7��=����KxB
�N�k�t���j��c-2Uħ���Cq��yS�"��c���ms���FJp�����E!k�N���,P��z�T[�4��-�8���u�;�&����W<���"vMEm��蚍b~S7��$��ݰ�K8ҹQ�!�����D� 0�\�����A�g�����|�r�'4�ֆ�.a1�e����^΢E���% :9p���5�K�^d�VM�/o�F4�Rx�Nj[��VǏ���5��.��D��XId3������C�������:)Y)\�g�g>i)�&~� �ʒ ��4��H�pԴ��D�>Զ]5ɱd*q�*�mVS���&�M�m/m��襥���J�xqiCE8�pf����jW[�1��!���:���EVeS�6��F��}��V>��
˧��� �u��:ȫN0�������1��/�qb�J���<������A��t�p��t�c�9�-�F�C	m�cL�#X@��USIh�8'�K<G���9�+?^A�7���y�Ą�_����_���O���5փ�A.�P��w�0|��㍁)[��
Еh�c�&k�:�D*��{a����-�XW�Tj��h����0�U�&_Z��f��[����i�]d�f�"��\ځgr�/,	�R��I���Ӹ�����z�t�	N��s��8V�􉤩_Tɞ��.hΪᚥ.�?2�I:b	͝U���J���Q��e�z����p%��o�N��5�F�!"|GB�L�����'G�,�7��]a���q�g��C{�W�C(�\Y��&�'�"�����j��M�5P8��ޥ��L�M��r��h0Q!-���j���7 ����om�z���R��s-�>�����J尃
#��@O��Q��YT�IV6��c0k��7�+�:�(�@ �O��s�}pL\�Vi��X?����D�&YNƷ���v��FT��)����9���|`��c����qg60bo���`j�S��K#oHn�uK�B�m�y�;G"�����C����=c8.�Ubq��ִ�����d�t�(u�^F��#ZY_��ӹ3cX2ą���ȯ���B�_��(�� ��@EMp؁q�
�|f�h���a�f�!��z�cED������+b�!�$nRC��q�C)��/$��;9ؙ��q����`��8U�Ϛi���7߽;A��/ �3��Fk���#���:�?�}6G�M0|�@f�?A�g;�-l���lK�v���x�˕���#�x/i�i!���t��	�И=���D�k���pI�-/��| c�����aIM��d/�Q���ZC0�)e��^��V�Q�/�Sܤ�"9�y�D�	7d�a�d�����l�WDt���-ʑ(�j�1�5_U�����ρ��J#	�d�Ё���	�r�̻�6@����4��۫x��}��X������x͹�;2�3�6�uG�y�����0���<���0 sEB/�W�I��f�˼�֨��VūHۥi���G���H�(A��,�n�?�$RNҼ~����E
Iɳ[k�=(��]~}!T�,t�_`#��%�I=������$ɣ�ر��1�Z��m@�� ĕ@���Ϭ��P��o/,�x�����`�N}���i���m���[��O���X�>�|����S��J�3�P
�W~��z�+�֊����Y�H/1����u@��t�6��w()�l`�s�d�E��t[�S�����hskjD�@4�����}҂$Mb�{�7���vM�U�]Zd�[a�e~W�$y��`@��;SY-JR(���B���S�u�r�^bC�bܥ�2�h��Y��,��`� ��hb=5��c�?�$5K�e��NLt�Zr��Q��t�y��-7��	i4eko�7�"N���X��V�,Վ�3�j�Fa %"5�#�N	
e��Ґ��i�6[��Uh����2�7���%rT#?�6`7�̔Ь��{�6��Ўz��*[���.{xU!yā	L�m�L[�ч'��E�0_5����W���r���@ ��ńz���2��a-~����a}\Y\?^D6v"_�V�S�?���FݗDф&	��|� �\#�z�FG����e�e�6��_� �H-XF@��F��P/�W�Bhg.��-1�x�~�-Ӥ��Ah��Q#��� ����C�d�c�+L�*�i?����L&�I r�K��@����U\��sj�{�W*^��9G�{~:>.c�����Gx�"�����E��[d��m�Q�+�{}�Q��y�7R�.8�C����({��`S�����n��=?]yp�P�$�POWT�V��nh���������o�cW�:ZK*S�����<C�ȓU}��a�p��{ktǱ��y���e	���U�Zy��,����O�i��
��j�<J��:�G'�7"i�S��KD�����-v�����Mھ��{�����a�+G�K�5=���Rb��T����c�^�� �T>e�ǯ�Z[��,��ʉ�C����1�$��M|�(��{��_�f�� Dn���n�_�p���C�41ِI8 ��Q��;�J��2Cc]N�ǘ�?���*�ϸ��7�مu6��w�G���_�V��H�����_*Ϛԗ\�p��WZk~�K	ܖl�\_HF`&���]���|A�Ş�P�s��`��h�r�$����@�.x��:���bҰ{�F�� l�7�Ӝ(���1j
���/2E\ k]��� +�<�w������y& ��4����8=�or"�ܕ�gE��c�-�B��ߊGd�u��2Wd�� 7��T��\���9�~y�|� 9��	�U��N^�l��ʠ��*W� S�&���r�@�q՚T�;7������Z�^�N!Ұ��>�=���'ݾ���}]�W������
�m(�D]���:�J�z����%����֬��tn�V�N���O|1��T�E��2Ϻ�g�IױkӶwP�{���n4��� =���F�|&�����I�vo�NW�@
��!�fߎ�x�KbP����UI<��S���k����pqs�yZh�S���0񪢝���݀�_�h���V1��. ն� �@�L3d2����V�����H�mf�=��аgo��P�n�Q�np�7��Q���/`���%�c�����\���±:?9s�ty��TDʻx#��(��^�6F�%f����GH(|�v��i��;�6�̌��v�_��#Rp���e?+f�<��&�X�Xf��V�����G��;�m�j^�8��C���C����/+%<U�sh�i��n�*3��:V�w��Z����]��u���s��L����_=����4�GRu��\KA_�C60[��p��a3���j�w|� G�,Ut��� �������*�WgN2i+��i2���ל�{ ���'�B /၍~-z	)M�^���e˶�*����)ur풙�OX�Y}0�wmT�!L�* ����m�;Lu���7��{�=�E�d�O�)�'�R4��2E����-^˯[�%Qq�Y�y�}{��A�����?Jm��m�{z��[�����cyb���H�&�M�_��?��R���,�R�Ⱥ�ְ�����J�w�K��Y�I�Νj�R�,���:�qџdk��K�5���L�$��8�w�������(��Fg]}�����Y\F�ه�k��ڃ�*��i�;��Ȭ �����PIDK�r�)��J�`RFF�f����]@!eCs�1*o�c��`�������B��䯨��J��=B��f7���f���RpN��F�Jvo���AqZ7��x&]Ve�I�f��$����5��n�vjj�T���@������,��.�CW	w��!"��m��+lD2��e�3��6��֚�6Jր�ƾ�ã��M�pJ�2�6l��5D������V�9&�T�(����1��n\A�d�Ů!Stѽ��⯛�����'��W�z�e�"iC�QX�����$���v�*ʜ�k2:W>ʟRiT�~�[fu��۱%�2�^I�Q��qnb��Z?��Ǯ���!U:D�6�Sxe���e�E�Y�#�� (�>�N<���=�H�2F�'X0������]1g �J��ɪ�k"u�}%�|!\W#��A7�u��P���:�4����]�)�;�]���u;��&Z�����2<���^�B�?<�Ô�R��J[���U+�b�,��T\JT�I9߬�`�J�z�oM���(�cPˉC���.�aa:8:���¥�9�܂������*���0��T���G�i�}��o��B�oҡ��9BA�Bf���FV�RnKধ�Zp]{$��u�8j�e����.���@g�7p$���$�� ���/V��T)њd��S���Z�4i��,d0n�yÚF�$��r�Y��<���?6�|YF�|	r�I*���AS.�݄�'<�۬�ͱ~�;O<i�9t
�=~	
Y��!����� ��
�Of=���%����
ޤ� �`�]9��ð1�������Q��+�h��ڏ�'8��&��M䀜�O���)F-�h���S�J�d%�xf�U���4\��2>L��6��L{� v.Y�O{�9߄l�@6t�V�_�!��g��D*l�إ$�aZ�K�i�ýB����!J���tq�I}_?u���㋌"!Tx�7/���*83��"�P�ao�X����o�m�`Բ���|]�^(s�Q��מ�m���]l�=�@hR?g�،*���4Ce��ȘWv��J��بc�Y�m�cd$(�<W���1�8&}c��􀓧a�8�)����9���R`͵���W0NG��߻����s%���8(�I~�
8۱f�f$�o��[�f�~����w��k��N��������ep��#�@���(�{չ*�3ڜ�=�@�����\Z��,� �SG�9CM�6�X����?��S���7m}��އ��s�1!='�}�9(��*.�)�#11�I���ѯX��TP����y��%Q�嘣��ݍF#_�e�.�vWtϪrR��$��Gn�O,8n�����鳅]���_��Ľ�}��璞�G�VLZ�Ahu�Ӓ��{?�#R�5�'u
��ޒ 4��K�H͒����'��8֐���B7nJ��?�d)��[�:_M��[� �NK��
z�)���[_���"6:o�d��g�]2���.ȿ�B2~��H��3�7S���ȯ�<=��/q���2e�Ib~�B�![�h��`��S����Ȋ<���J���C�+��|BNc��E�z�����5&��%��K X�����[\�W�k�]������2��Lu�~��K�ѡ4�i��p+�s�1�0$T��؍�'�b��~�=	�'F���S�o�7%֋$O}��c�E�,����5�3a.�$��wXD������|$Ʃ��4b~ŏ/fM&���cJ%�<lB�?r�8,�aT|$DA���#C���L�ވ��S��zQ�171�3S^�f�7�䒼�^έ,rS�;�at�L�W&;<�)����yW4���'Jz�&���q��f�h��{G�U��3�+SC��e�X�85Wܾ��r�S�Gw�ZjÑTqFD$��Z�Y�Q�jCX�r33�rJw��
�5XNV��jE��YKt
�}>��(wdx�RA"+��zj<1HlS{�[�N�L3O�s=�0gfe�I3uhY��_��蕜o�j[����r@����:x�0�A�����d� 'j�80��C臕S���0|��q�,�w.��!�,#C�)Z���'\��x��5T"X���9 �]����^���5�^]�y�h��?	'qCռNT�Lc���1�N�f�O�Gb��cU��?���^Ly�pfR���<�eV��A5S��Y�;��JK��� �*���")��I9�'����V�S�q�"����Ѽ��gD��#1�5�*؄3�&Z�]��!�7E䜟$�A�|ec�_6���,���9�>�d���%��g�8�Z
1���I���54���Z��� ��(�)��kd̩�4���U�+Q�䢊���3��mZi��axjxY����5�EG�*�ɧ�`���?@�2*�����?ɚ(A�)�o��c�a��~ץ�����'S`8������.�u2ũ̪�&��0U�ȃ��JL��� �с0B���<]�Q��� ���=��O����Z�Ӗy-�	5�>a�"7����tn�.���8k�V���X2�fUрr]�#�A�K���3XA����N�#�\�:�sHL$.\qwp5rt��:D=N\"ݝ�~��	�#�!Wn����ړ��$ª��H�"��r(�(�d�6DU^�vtу(.��b����%�ZR=�����saD���z@N����E<�/4d>N !��r�CY*|��u����Z�
�(pOc�����,�6�d�!��w���ӲhOܓ)ꮚ�ՁUR/dQ��g���q��"`Ƶ���ء%@�R^i��6�A1���8�W��{}���$�9~��G�mм�j����S?�A{�8�t�"B+(L�n9d,���l���l���$r��� ��z��Q�Q���lW�zQ�&r��J[��3��C��H[ j��AB�ۅ ��ڪ4G�+Y��jD�l�ǝN c,�j{�)�Ni���@}��"M���<A�P~�`+�h4�a�Elʨfz��2��"�� >��bv6���G?���M��JBےtƘw��.�)87� �i�bIѪ�$����Z}n�QQ#�2�x��d.�lC��>�֥`2�v�Y��ө��}x�?���C�sm�I��/)v��`�o�e)N�gw���Q;�S�r�)�j����b������wE�);CF��)���s
��qe�Q+W:.����[Z��h_m=���J4��Zѭ*ږ�&$�C���(u�c�&SeB�/�3S�+�R?_�N��j�W�=�W��A¿�~@�������n���I���[>c7(��aO�]��yӟ��؁t������w9�3{�K	Z��(?��p��E7t'r�3����b�br�N�Y�zFl�_#�j��UE��B��{R������)��}Q	h+�s���l��I\^����j�aŲ��#��������9���3�̡J�tm���}}ĸ6�|W���\B���kq/=�� NUƾ����j�Bszd�e ���Rw�|�'�[���b�Ϋ_�11� ��b�0L�]�g�T��4w��Ƴ�Y��c7(�t(�`�*~�% �v~��Y�B{G�?�pޓ�*.I��ڎ1�A��Ć�]8�/M�$,�il��7k�MT>�R5z�E�O�e�QW�Q���?ί�EuN!�=~�O���1�⋌��^"�}w���^�M���-��[ܜ�����v���<F�9�q�����7��p�n���'N����a8!�����(�]׭[��u��a��2FR\|���h̛&��\"Wq��J˦�s|��&Mٕ�F��įw,<��cC�,�ƙgYðhP�����1��jH��|O���4e *>8q��:�ӧ~�PPj+1]Tڋ�8�BN�"fݛ�;(͛ߠ������:P�����m]�ziQ�".�w�
N�J.2.�7�ξ_���ǭl��&\r��@U�!��}�q�\&���~���ΑBlA�٫'c�	9�O!��p�\�F\��R��s��;���R��9^9g�O0f{?B��<�X�3[�o��%��_�vAҩ �x�o�^z�
�S�m�UJ����X���/�=`C-"�g)��O�l�>#�	�gry"�w2�F�O\gC$;gƺPy7tc�"�;�!g��1��������H�_�1���-��<��gQ!�]g>� U�"w�}���P��S0h�sV
���F�S?J���?Z�">!��������.c�Y��H.�)o)A���rۏĶ��=7���{MZ1@�]��Ԗ⮰�)o����6S���/h���������,��U���QO��brICv��S���'1��9W���)���S<�b�ڼ6@V��P�uw�	�����雭�wu�ׇ�-|�s��<��-Z�s��"�e�Ըk9�1g��yb�Tgk^����E*�[�DU��ߖ�/�V�_;�XM�p�Mj:i�Z���_{cЛ���¾F�=)~:�X��N�q���G�-7!̽X�~��옪���rF�ӖN�\G�l�� ����*]
�0�b(��E�c�7�<���,r_H�?x�m�*H2��=�>�Ն�F�r���퍼mEW2�֭*ە�/��	��5�k���<��8��� u�`7� {�1�J�]3aVw��{]���'��M�7v1|G�\#Jό���$� RW��`e��ڸ�az��d�H$e�<=񞯆�h6���I/�����<9#J��,�βye7�s�m]�nB
ٵ�M�?O:y�_o����Ah8��rL~��4��㑔��VD��W��2>�س�m��\6���wK�Pϯ��� ��k[Ӈ4:"�
�c�N�!����s�k]ѵ�w}���ƣ�w^$HaZ<��8���N�1:X `=��)��8��Z��V+��10n��o����:�ɷ�X�o9���b�g��y#m3�`�i�c�uHє�+����O�%�]>���@9�_����{F�ƨW�0Y�Mј���#.�~N!ڜ)Я	1G�CF�<S
iAI>r)d��]K���+�{�T��,�%T�d�`W��_��E��9��﫼�2𗺿�v�����=��\���Ө��v~ffn\�]�d�r���@N��g�o�(Y8TS������m�O!$�:��%�5=��e�r�#���C�]����u�ٯ��q�K�nS��oba+��Y]����%t+�p����1�������E���)��Op������ww?���k���<v{�6�v㕫,k�Ƣu�z\����7������ѥbv��f��ӓ"�-�C�KK!ٰ�+K�D�e�:�T.���E9	W-�������'�����+��O���!7YL��e����(�?th��m�,B�*��C2&1�	�� 2M���4��f�^~6����ܺ&��
6�=�ʋ')'�����3^����᳭VO�e7z[\��QU����	{>f!-g������xa�k�G�y��ez�)ⷐ��?M�W�a�A,Vu�졥�غˇ
$��T���� M�zf?��9 C����r���<�Q꠹^zx�y@�?�z]�����i)��$=)�"�]���	<qD��Nf���n�[� qk�u1������8X$3O黂q���ڴBm���B�I@p��=R�n0"ī�UiD��=G��[����",�ܙ�fM\��scz��{:��o�HO�,�y\_H�-m.P U�A�	w�τ�/���HT�5O1 q��[���<z��R�|��Jz��/��������������X���F���V�[p=�X.�3�� �NR]���}؏��HC�i��/¦����c�#�|Bi?,�/g�~W5�{BD��er���j���]WW����Y���D)��JA�����i�C">��-G$!$U]����z�c{�ME��DI?�R�u�^�T���j����9����UgHyq�A�k9��[���P�5�Q��z��&�)�k;Mp��;���&>��s��Hw�,n(e�s�w�ד@��=��#��-��G����(�9;�pu��d�@y}�P����}�w���E�+�i-gZ��*��/�%Y2�\�a� .�@�]٨���تbM���p?_�(���v�:�K�x,�k�{��S5���e%+2&m=C�`��	���Yy��Z���
jUl���n�)�+U�5z_0ß����s�A4�B�Q�����&�^Y�~�ň�Vo�	�S:�he��s�������L�^�o�[S��$o��엙q~A��f�� �8�;��ʑtD�*��8G��{�h0t�M���GU����������WI"���Y�4��$������˻��0Ν�����:*����I�ͦ�'F��P�\H5�-Q��t�����.'�ja��V+��}u^����<�{�zv��e�(��ғ�p�eu�`q�;zFѰ��7��u�w�yO��ΰ��H��08i�p�k��լ�P���OlYۆZ�}�:��Ih��L�o��}�|�ĳ����
a}���)Rw��$�-�� ��L��!@`Z_��F�����~���RO7.e�X�QYH��͏�n�Y�O1���t�X�Ӏ��1�����R�Y֏jWyOZA�����	��of6Y�(F���m=�X�n����i�^�^���g���T��1�H$N�H�~;�Lf��p_��*���:c�k�7��y�R8��	���	b�߃}J}�jTĒ��T$H���]�t��8�CKUQ�y���Y�Ol�|�I�8�R��
"+�lh{wS��^��0R]U㳬�,}�+���쮬��R&���������F� G_ ̂0V[:�w��B�`����ȵ)���d�_��C�u71��p�o JqH��+˘8�S�Q7,�E��!����N��ߊ����E}�����V��ģ���B���J=�������E[�d��/�%_Ä��Ұ��a�0�]��p��	�t���ҿ�z�g��=X�i��s&:	19�hr4;��O����g?����~jM� ҋ�
e�l6�gM���<�cb��?�Sޡ�
X-���W�h�=�\̚Ⲥ3���|��u�7sB���d!�z��!�����Ŏ��{^���I/1!�O��P�fM"��a��H�BN����S�"�r�����ϲ裐��p$� BB�^�Cw������GD�mT(��!�w��W���B�%��yk��qI)���&]�?�ٖ��f_$��\j�!�X��H-��m�����Ƅ�R���8O"�+�p�?g	�����^�p����^�XznD)qjtSE� �C.��݂T�����kP���B<m�x��kM ��-Q��J����&m��8C率0��A�^�S���4�>�'Y-���N��9@�y�u��A�x�!}���vw:�u1���*�D�2C��z���8,Ԍ���A:G�ws��/�Wݷ-�����'�d�G�z�������de���ڕ
E.�J���Pc���2e�[�
��゠��Oˤ�R���t4u&�F���A����O)rۊs?Kf�q�|�	��$�>������)�a]�[��S��l�=�v'�Sq�U�� ��P�D���q)���$��[��k��(gvæ�dy�q�iw���H,�+;qF�:�5�cA�fp�D�g4�%�H��)�a��_��|	D��q.�fq���ӷ�N-��&1��vB����{�����c�	
��#�l7�<��HZ�(�)��\s�|�f�ӣ�iCY�wZE�e��/Y��<2��T~z�	�YRa �yR"[ǷXD��6j�S7���rL�SDP=!��fɬ��0pd�@51V��"���P���ҋNɥY����Y]��!�b����i���(pt�?Q� ���+V��bFb$ ����������ms�3 {{��������0��S�p�e��=r��"+��QA����J#g.���� m�x>%y��i�F�Ίk�6���~�wJ�lߑc{�;�����L��U+�!.�}d+񹺒Y��9El��̶�^�N���_ye�v@�-��>�2xoʎj���̙���J{�]"Ԭ۶+4���D�³��nsO `�)�~)3��"�6Lcq���	סM%ٱ�Su�j��7�{}[����udΈ��<�	B��Q�\[[	���~*��<�p�E�����m ��òK�0�P]�UA#���I�u�J��-ɏd���pv:��:��[��3!2�SPǊ�p��#A�gj�u`��H�}�l)�ֵ� ���nd�U׿�[��x3�&�&�z݂Փ�.�xΊ�U�5q/f�t;��:�3�yxI�̬iŋ�]3����깄�.H������Ơk��,�ˉdu[G��K�{}_/�e��
�i+�-��r����D/����zD���ݨ݀� �.�"~�Uxy.Gu�C��"���U�9md#�^;�d"Ր�2g��D�3=�>�`g���9��I�U{9�ec"m!���4�~� �"��:�j�]�=��	#e���ܖ@�՜z�x�H2W\]���~Ǜ�QQN��X����N��aK�>���C�xs�6$8�=�,�*H�W�4%s�"��xH��z|�_^�ذ{��J��k�3N9zz�H�d�8U6��ª4e�7��G�\�K��N��4��@4��2)w����@��qb�`�&�j�h�������1ٞKP#N�Ϊ.;&	��E����j`>�)r�J8dw�j��Ѭ<0"R��|�	t�9U�����S����}^�,#���57�?����@��ٿx.�]{�(�TC�z�aWr�ۻT�X��~��Kf|�t;�3�Ҩ��)'�%�C��8X���7�c�/�W��@��l5qW��lqӱq�F�xT�\��&��
�❁��x �eё�J
���`h�WBK(@;��wn�V��R���}j9~
V��8 O���aL�~?�ˤ'B��"4Tۊ�e7=�e���I6AyM{NX,���I�]n��U^W"�����]�3�j�u����U繯�m��s^������/爞s���cЅO ����!����*��袯L�п%�A-���z�J>
x#ߺ����[;��rfk��rhug6�pA����"��H�	uY$�Ci��ro��5xW�R�6c�^5�K�𤊆���������|�����Z��b�v�)f�5���s�"}��� �	�^,=���Ŋ�-E�q��M����-��D{؛}�M'�8��۵��_����O�;3u4VG(�bYzŨĕ�q��R��0>v,�|٧��U��G6y����O����Z�!�^k97�qYm �]z��$�F���r��z��� �px�0�:���w#����H��/�ɪm2K�
~ּk�	!�A�����x	��Tt5!^�����Ӡn��ZH�T	6$�D��@I<���1\�v�H���G�/cq\P�'�mJ�_8�t�0T���'�,�w��x�B�sT4�E�7}����7]y�b�\%^��V���)XH�\�?~��x�<\��r;�^����t�f��أʌN���W�=�	�ɴ�^�� ����,�W�H��"^j��>�[�m��5-I�����os�B���>��M&p��BIR��\��F�0���m��.3^_0����d������\	��[��|�o|��y�B�� �MBWNAD�I^�ҙ1��r{��y!C�C2��9�Y�y�g�*E�HI�9�����{��w���怛��e���\!a/��,�-�qha|��:��!m.�sV� ��<\��[D��T���≬0p|�_�-�~Iq���{�uk�y ����R3�e����y0j��ڿ��(��!�;�O��V�M)2t�]�rt��psӚ=`*�᠌u�)���x)���m⯒�<�kU�!K�,�t�;��C.u2��/��84닣}�����:i�7ͤ ����J���@��]ӠN�U���Hr��S;X����C��GӉ���d
�0FAI�(i��t�����-��z�FC�-�/U�.#��w�R�7涼[ ��3�j����8�'��_Pex:�'= �-��:+K���}���\="�d�v�wF�j!��J~qsCb~-C��dw��?kcv�TdaF-e-�?)£�Icg�􅕑�-����J�0��$(U���a�c�y�#*:����ƭj�����OC�
E�EK� �4�ksx�y�[C���.�����>*����_\@N ��o�cϑ���� ���l�=����V΅�?g=pR�$++��NͰ�FH�j��ܾ�����'�9H��$�Q����=;�<,7lAh�DJ/e�4#�����L���p�E�W>ZL��m�L�*L(���e����/� �L"hϕ�&,�N�4S��#1VeN�;V�O���}ru3�X�M�*�����{�i`P���$i�Mף{�*�?��n�������ݥ㕷5��_x �����{�B���'=
ӑV�3kҩ�m�-$p ���3k.u�p�,�����`v���������o���VƤ�qN���7�a�@�>�s���s�Η�\P���1�J�g
Y ����j=ȡ5x�%]�^ã���U��_�)��Q�f�	fy?�=�DR��2�I�ۮ�ʷ�]�{��\��smW^�V�;_Y�[D3�w��jubY�qHWg�Y�5��PIT�`uEw���њ�T_}n�彺�н7�.�ӟ�'�Cy�7�Y6[tw0�P�I�������1�z���:8���gl������� ܮy	�	M_@-�I%���2��P�@q��j�3�| �	;���|���_y��p1�
��\Ș��-Nru��,x�o���u�Y*�j./��s�Z��W*6:5ݼ�t.e�&�N>���ǔ��c8p�v=�a�_�kpX~�S�~,C�v�b�1�+A�&��l�芒�Ȯ�/��Uq��{>��o"T2��\�U[`������y�#�O��yffݛg1����!)� b�'�m-iP��B�[$�^/�3P%��Fu��fm���$|#�T���I6=�{��z#�#I+(f�������:/ȇ��;�|�A�!Q���� ���<`�+�U���'aN��nSL�;��t�T����E�y���%Dj+ΐ�Cy������,��K���3Z�P����T�.͓l���A�T�HՋ+�yq�wL?#�
t'㭠�&�$����P�j�����g�����25~1c����2�NGgwn�J���_B�&�x�W���/|��yzT�/�q���L:���J
(����!�s3 ��@� ��T��W�R�?�d2��D;�1wk����h4C�7W�݂~ ^4֡EM��V�y�@· �09���VP�j���P:����Zu�-%$�����*��$�@��tj�&~$ẛZ9�~f,،��Aftv��]� �K�t�&��b/�7WD��n��"�%��At�Ư���j��H� �HxMD��� 
��A�9Z����R�M��R��t�`<���m�3�cm4�!�;E�Gȹ醴Q2ŀ��n��Y���=o��0���i
�2�O��K�NG���9і�l���N
�'!��4�4.��&�W��y0<�v��
2θ���dH�D�[��難;T�_�}G�$���I�Ĵ�J{��c��@Z8����1��Bldo�O���ݞ��N���FL����]�B}'�;����AG7�1\�
0�Sڊz,Nm~�pe<vu�cn|=�]>c)ɳE�r�	_RU��M��H跸a��JB��7Ud��5	L���Y�c>��+}{��Y����&��|YI�) �� ks��r]�WfyrL�2jzuz�0c�KqFxs2.�W��J��s7Or���y��]k;&�8�
}y�����Ǆ h��m���fɟ|Ą�)����R;OcH1u�����߆@���&����7U�!ob"�^�i�����E��J՗�(����o�l�{d�!Ȱ)H��E#��W���}��|g��=�Q���R�A���ᨐ�`Ec#ӏ���7F�p���Tg�a��xy���T� ��@"	�w��
��=�hl�l_J�r*�9�
}��E�H5]��	�[ѐ��,�e}Ǫ������pP�bru����܆���!dZ����ҙK�� �]�?��И�Y�����̣��*a��w�k�����5/4���N��3B\��L���6��ܲeT�i'���8Έ��������0^&*��ӃP���cS�+�k�	�{M_��aU��Vʚ��}�{-�ۣ>�1��6 	Fy�ֲ����l_�ch��潞���g*����#_W9�(/����qFڏ(������8�gEE8��䪒��G��f������=,F��~?p���Ҍ�B��9��1��r��bS4��`���c��7)h� ��ϒ�s
˾kAV0��eC8��2��:!��-��M���* ��s��#e*KLL�3j�M�9���=L�i�l�h�H�m)��e���:2;q>e�:�qU�������1<k��b^��wZ\ön��3}
����Õ9Ӳ��� ����Lcu&P9'�GcY��ם�
��띅�	�l�8�$��9"}l�Qt��@.�����^��K+E�!���ݩ��
&kcF�K��Ǔ`����\�G>�Q	"6�L��i�b��B6���2b��m�L"��������*�����N8�������uҎa�Ů��2	�A���&�v���Wz����W &�1~����n+&%�ˀ��4�2@~�l��k����E�H>�D9��;�U�S�݀B=D�+�$o^�~�s̍GX�=�u!��2��^X��yF̻#؍xLGڗ�w�J1��B�a�7�s�tmW����w��GV�����`����ܖ������t�յ�j��3	��W�^4��O}����8�G��7OV��iǖ�U��ºo����1w"u�z��%$z���~
�~�r���q8��\��'���m ���Tqh��,U�)u�dz�� �آ7(!�H�,�9���LG�,"7K�DE��
K�#m������:O<5��)9��2ť"�|�G=����N�ߠCB��f;�@Ǿm��>S��	�/FQ6��y��F�iA�uRn���.�_���AH���D�� $"hcǌ�ՙ�I��We���I4�?���W;���Z�!��Am~��o�_�F1���-�;bn�tw���8�N��4��],��^���3�ŧ�-m??��MC]�\��2��͛�C���5�P�'�7&���R�a��=�@�8����P��AH?Eϊ�����^vj���ӿ�{����c�-���w�tex8�>u�#��X0���v\<�A�#�4����EOS�*ҕ���z�C%�Oۙ�8ԑ�
AY=�(N<L��'a�س{���R�#����d�ԩ����P(T�����q8�c�؄�@l=)2I��2p厩�:�f��&R?��x��jJ{�U�c�8k�.�Ȓ����Goo�Q�X�dbdR^�7쒂�5D��y4.63z��R��mCT<�Y!	��[`�/~���� G�>v�B����v�̐?��k�n[!���2��(g�QJA�R����CJA�Q�:C�p�S���C��Q��krZ�F�6� �=�/�	x�0��ny����V�T\�3|�>���M��0RgZsZ�)��ӀG)�|Ho�4�/X�ט�&l7?d��F�4=�ɕ�b�
�vc��O[�����L��\�٫��94v	���ƶ	��7�yQ�뺌� Vl����Ojc���A��j�{�o� ��� o�����~;s^��"�*S��@)�����^�h�,�Q_�8>�k��/���O�HjR����T��q֭!�\P�q��Kهl}�5�U�1�Lو��~)Ba�=�9:�|@|���e�E�J?z'����{a#�dą�0_=l�����D_&���z��T`V����I�w�?����`v��ɣ�!`O_���� ���(bi��I���V�����zwY�����*�VjY�� Q&�ww|����R�d;[NV&�b���寄�X#zǯ<���[ʽ[ըlìWO���)������%C�|�ዷpY��7&?-��PE�vȹH�|�G D�@FFX?\%y�u��g2Y��O�Z�7i�C��y�k@�o����7�ũR��*��=�&#��� �o��GG�:J�6�NQV���%���ZJ���3�:���h���eL��͈����W���5*�!�����9�TT��~��Ľi�'�<���/�C�@ˌ΢G�]�CG��	����rzx�l���\��t����T��Q�]3c����v�l^ѱ_�������G�񈟥J-w��x����bA�u�ھ�k��`�:�ZfI�tV�U��_Β UNG��!N�B)Ֆ9�s:$&B'���٣�M�l��<���bc�rsHc��e5~�g�.�E}=�jK�=�����r�Ӯ��
�.=x�|��<��&`n���Ȩ��)��'0�ͥ����\[�X~M+	�+J��p���@q$Q;�����"r������H�|��(A?����u��w�Gc�D�ڧ�A��:i����z^�B#!X"3Ă߽��8��y��]p�`
�Z�izI�Kfq��-p�TRj�6��]��
��5�1���q�]�oe��@���$���Rp �9���3]�`�x�ҵrr���9ςh����iE5�yRP�բ��{�4�����P���Б�v���FD����K�-`�X�)��Eg���I R�`	�ӳ s�T�OS�*2CZ0�Q�'��1�zC�Ꮆ7���k|��
�-�ۦ�;�%ׅd�sҥz7i��tγ�?S�ϫ?����As꾌u.ZBC���%�	Р�7�����{�Lr��]du
�~fv
��t��=�+r�-�+�`�s���Ѵ�Hg�}��Ȋ��sE�N'������(P�3d>;V�*�I$;M���Wں5�iX���J�ȃ�e��ݙ�0��6�"�`��EøtQ�J%�]�.��;�G>�� �4sbO,v�!��d � ���>º�
���Ҩ*�E���Ŝ��'�1�?���Gc�V�1������=
24�&WP3��+c^^"��&��|Sxw2(�lͧ~#�B=���_�@�2�2f@�͖G`�J���f����%,��P%#*�����"ˎ�a��s�9����eae&c*���o<Cj��6�P	+2σ�dWt«�x0�n��ݜ�PrTEpi�B�Z�{�v�m��xoӺ�r�\WI�(��g�*� ����t/.�kYҼ�1#���w=Cc�s��mݬ�&Q��A���}R�s��p�w=����l��#�C���/M�@�r�^"�+dHH�"�.��w�������̓�*��e:��M-��8.$�w'zm��U4cpE<��.'�]�j��.���`ǀO��V�N��ݜ�#�HU��QjD�r(`{��+�T@�N�?τ@�2�HM�9�R7-<��	-�Bi�9�4�
CY���/��}��o�����cl����c�'�-!#�����KG?Ajq`����T�ǝb6gK��҇��"ޞ��=
V� o(�)}⤫�Qe	��8�LC���Z�C�;���c���#\�a"���R��^Ǥ'W�V���a��ܠ��lv8�Y:Xq#1O9k��;-��U����^T��u�E8�|V�+C�/d�T�&F�e;K���N�v4p8}��p����d�����@�<�1��	җ�!. W����w�����Bр<،1��]	�jI�����huc�}3mk0�]��_gɠ�߳��0R�]�|Z��G<�K��W��T�%yaM+{U�@@T̪tC���@����N"��3��v��}@���*+m{���N�D���à[V���Z �e;a�S.S�K��<o]ܣDS�W�A�s(�O0��<A��R�X��K2�-�\j ,��~W]��SI������E�r��)M<
\�-8�h�`u�\Rc?��O���\3N�j���s�������[��l�j_��k�gQ4�["m���k$Is�����C�lc�KM�C����Gxd���X���e�&}��WH��60�!I�3
��@+I��nP*d�5#w�oL��W��C�"��X頏����l��-��ђ��%o8T��ㅡ�ɨv]�Q=�'xPO����+0�E�Y�n�#�q�/�0ݔb���|�ݬ�!z0�"�?CR��H�;l���5.�/�"ص��]o!��s�$���|3y�8��Z����S�<� �ĉ7n)1e�P�i��?U��h|��In�s�����t������e>���-9ok�&��,d�a��nKdlC�����1	�'�D+�辻\:��w��/$?d�������ph�� 9��>�̎gYZ����v-&Uy��3��8CR��9��;9�9q!SŪ�!)"��_ܼ��go)l۟�g���p���y'�	 f��:��b��NU[���F]��v\i��7�Y��-`�Nr|���
*�/��� ?6�ɫ�bxl����p'�ǽ�H}���B
H�$&l�����i�}�J���AT��[��ư���[��%5�Q�W�� d��t@��rT��c�nu���຾�_��93�L�_crE'�ښX��sNkK�?�J6M�_a߆��`r�����w��Ld��CvC�4��U�2Vp�ڧ��Ch���J#��tָX=���4(κ�(�~8ݙ/�ؔaw�-<����aZU�K1ʏogq�9�eJ�P\��Jq]�"�T��*M�ְeN�"���hA�(Rl~*#��Vp��*�
���ؠ�T�Y�:5���;4܌x\I ��?Z�_�0.{#j�Ml�$��=2�!ۙ�I��e.b�#Pv��H�AfvN?S��������؈�+*��>X5�ٞ�c��\�t��]�*�X��r@��γ�"�#E>>/�}E@���nc&��]Iᶾ�fy�<lʠ|U�7���T&Ofd��u|��$�`�!�_I�^آ6$����N4Y0�.�>fR��4X��X6��~ @P�5�YM�z�}�A�n#�d$�Q��3��$J�h�!C���H�2iMXe[_�;X?uÏ��=���p^t�&D����D�{��
Y�%��M����P�9��x$�OD�ʀð�g�H��!#d�7�Z❮����29��ˮy��3#T���Q8;�~Ű���F�WK��A�bvl���y`�ݸ��%-�`Z�[^}P-Y�K����3��k�~���i��ӈ���mS�Zʵ�(�s��t��1ˌ�E3R���[Y�;���'S���ow�_��]�*op *Gq�Ƽ ��J�d�{Vyd�z���d䂚.�߆_�@"q̚ὅ0__���!�#a��2a����$��G^���	;WC�:����E�_F}�����*(8��[�<�.D�����|2��<ܸ�p��}'V��A�����x/j�A��.I��Y$]��t
�;��()m�q�=ʋ�J0�[>��׉�N���k؁r8bt\��Z���#wp����T�� ^QZ��Ѡg��r�}�:6?mmdƶ�r�4�� �Cr���!ɉj�`f��԰ޢ��$����s-���팥Θƍ�^.�5}!ec���zn�|"m35?�D��b#�٪qXǀȒb���	w�ټo]}������&r��;�h����¸��ly0���xc���VCr��1Zۉ�PT�bۑ��7{������P(��Zd�E��z�g.��%��i��B����s2h�/_�!�v��<����_q!�ƝgC�[oݨ7��#���i/*/�-v�#�hyB�S�)�83�y?$x����̵~�/'(���DHo�Z���6wB��'���$�XT9b�N��q�X-���8*-ޗ�=�mX�P9��u�N�T�L~�b?�?��_���.��~�W���8k��ײ�Lzb�	���$r�����/�l�_,�<дs�t6�����4���+�i@�	,z�Gq�ӸR�/���Xf�0;=k�ӓ�T����^ߎY��F�'J�DDɗ�6���<�h^>շ�Z�L���&ϓhۅף�&�S=��ω��zS�R.��l�|���B/�{�L< :�V�6J�6?S��L�w:�^�H�hG��D�83<�[�3�cjȆ|'�ОXb;H��;�dyT�?;�:
�6	��ԗH|L��8h���ȇq�sMG�����kR�|����n�{+C~�Ө��;xw���������ʔۧ5t飼�����0��.Y{�2h9y��vX319�C�ܢ��IN��,�v�as��m���.S�@�8���~����{ ����n�B#ʾ�A���ӓR���s���C��?6�jZ�a�������I�N/Y�,+�Y�ڧ��B٧C��mu̓N�W0]'>�_�z����C�!�ҋ��Г�Ew�`��Vߛ1>A�t ��>(<H��X���0�1kgD �Ǐ!;/�\����.��^�@��E��}cb������F�B3����yXt�O��Jvv>E�]w�MY�����6:GLw3�4�Nc���>��/�3K	;]~O��ĞWCH���%Y5�Ō��
�?����{���`2�X�SD�����Q�1��0AR�/��V�.˞�����㩑�ӎ�� @t�j)ѯXS�a0i����s�K���iV ;�Q9�"���O�d�q���L�ʔlD�)��U�5]���c�\�h!�E~r}יEN��B-�8O3�������#v����[�:�S8��t�֢���^�O(_��	P ���3�9DR^�L�����}���[gQO�ձN��� ҵ]�i[m���q
O��X6*���ڠ�<�./,JY��U@fU¾�}��.�c(�g�G��c6(� =�P@��~��j�9��Z5�K9o8�$��)��+@N+g��}>h�@o���Z�x�SK��;�36��+��]�£ѿ����sF������FG�NmsM<�*Q�Ctj��@�V�N�l\��w�Í�0���m4f=~��7C�6�E�Ձ�23m��S�]H.>p���B�4�Щ��d�X_�;��5O�>a�=B~k���J����"��� ��o~6Җ;��xN�s ]�C�U&�7ɦ@@Y݌@��m�'=pm�ˊ���3��uɷ�Z�@��ҢV�x��ny74�طN�X�o�dק�<����B�:���K��JP����������ߞR�����p�U�<�#5V���M��lv�q�e���� ð'��PK���k$��+��f1ef�d�/>l���
�Q�5b2�b���]��0��(�6�^�l����Y�	Y�>�Ł�Tk��|�7���b<���O�\+h��2j;n�aC���3�Wz&�����v���B����067�'�;ь\NI����������Z�������-t���Ȧ����b_@L ��]<�v�D��n�&����9A�_(0��+R�/��>Lc]��`>�e�
�Qef�έ���j(v��۟@V��X�!8�Ƣ|ن�l����'��w�KѸ�!�4�6ARI F?�y��m�t����|(\0�W/E%�lD�mB��s��H���H%�aW����{6�O�k,�Vf�m�VP�>R;7K�kO2a	���b�K��� o`X+�Khq��<i�b��������K��[tl���F��E"�X�P [k�q��� ��1�RO�XA{�sm�BW,�� B$�I:�a�w�v�4].2_�i��I�L\Gl)�'�&�9:ե�IUp$	"�޶r��ق� �����P1h���~�]6Nd�3�^#�$a[��D���ɍ΃3��N�	G�)g<`(a��6B{����I�����p�]�:�IR!�܊e�&�����A��LA��8�髳(VR4����L��P�G'��l>|�G�$�"���[P>£���G�,�SgT()���<ɽ�}����$y�+@a,�}��
mHc�/~��;S��1�%UP��SqaF����u�Ɨ���a�s��0�����|���ݝ-<q���j��d�c��nj�V�Gl�9{��%Oe����3���+O`�ÚT��0WI��m<<� �۰�� ����xO��$�nx��ԤY"�v��h�ݳB9Aws^��8���1�n[Pnj��M�d����j��@A��nLDwĴu�֋?�گ�ω3�s�;.��ۣ1b��6[�� JDf߱�PqcM�����0�0	'=���\3�����ɅA�=��A��xy�����e��0��}xwva�ԅ2�{k�4�w���O�c�"L3�D���4Ȣ�x_(5)��3���-,��U�>��^��}��E��P#>��` ܷ��#\�X���ľ�#\�̘l�8� m�(�Ru��o����c\�Av9pC����>�J@�S��;��sV�Q�6�$�W�d72p���>Y:0���s�ik�
��FN3�bLX<r��������n~�[�KM�B�(X۩.( ��|p~(F���f�@������~����k]{�Ӧue�E�����64L��Y��C��o�{XĹ$uӍH������؜������Aaîz�6mO|������WH"i}��>�W]�Ibѹ�e�h�dj��#�!oH�L�oXG%�u������}wB��=F��%�/��0����W0ąpl�G⬸<s�#�����,O�*"��
�l���.N�ɱ���a��Al���)�"�m\�zkܙ%�׋��f�AˀR�<�J����@�X���Ηʛ�݊l}����;<�a�Kww3+|������jJ>��-ܮ���_�Q��m,k�u���s4g_��#8�Y�μ΃9�4$'Ҷ�'��;y��c�9U��V �co�I�)��^	��i�250�9bHq��� "�/�>ݾ�C��7���A��f�Ҏ�˕��ǃ��EM��	��4�,Ք��=�c;�=M4�9�'/��}3�s��Z��|R�8���A9#~o����3k�M�֓��P�!��,ή��æ�"��9[9��B����� ������ ��r7:*�l9�ށeЈ��#ź�	Eq� 8�mw/9�(�9�_?Hb�g��Q�6TN�]e�-��(���[R�mO7��������hw�)e4(|b���Ii��F��yi�[Sc��~;�CxvF�����	�m����d������X��k���rg�=��gv��_j��n���t�����X�� {
C��$�S�i��@1)�-�-!�d-d�.�FU�/�R��H*
t1mS����5�	������NY��K��Z���Va͑P�4_t���CeB�!���	�� y9�݂ٵ���ޛ����^5�6�e����Trh�$Bg��E�
�N{����&��F/uΏq�)T�����{X����G��bC�a8�R�o�!{�i�4�/�v��*��)�.�Y�����ֺ�Dmk�����M�
���(u���:��1 ��y�2��y�Q�}dI��Tf؝d�x�,I��ڝ��>�"�>��č0|�"Χ40c!�o���:7��~�1�5Ӓ�J��Aꈳp]��3 �H<���<���T��j�9��X�w�`~��y�9�r��T?� ��S��& �_= o��U���K�ŇWv�z�v(ä��o/_�+���+�׷��M�q���7��w�(z)3�����%���\xQi���L,��d[�=��([�:l��\��B���z!����!�ZR��3�>�}S���N����]���w�AeH��7Oa�海�~��ZB�#봞�n&�:H6^�bL}a��b@��z��	E��<��X�Q��(����q�Dx0Ȱ�L����c��;�")�(���lhm��6%�I�vغ���ה�O�q���f�#{S�jC��/(��CEdcĊॠ&k#�wp��z�1���4GX�x�Ti�tVY����l���HA�G�pOʟ�[��I��%�?'����zlc�/m���P�>�4�Tr�!oo��ls�M��N��k����,��p�&���1qa,�0�GwA����P�]Mm���I����f��C���K��:z]|�*�Y�a�DrL���Ӳ��Ef�gtU�ɪ������-C�K�Iq�"5�gz����#OAb8�I���U/Hٴ�w���z�bZ�z
qD\A{�\�5w��%㒄�N$����-��q:�Q��D�������\����]$���i^��;e|=�H����l��뒞H;MS�#��c5 ��.���'����,<�##a�[W!�7�&Wkݘ�X���2n2)�=`�%��;W��\���,���(W4y�m,ybr7�l���"Y`K!�-&`F^��u ��
&Y+�n�Z�w�j��e�K?AB�=m1��':?���[Ě]k��������D{aK��WL�� �p��R���<�����v��N��@0��TL� �?%�r7G `ZqL"��J䚞Έ��HKA�����������i5�9�(ߪ���V�|�vȂ�E(��zo�/�*��LO¢[ɐ踋������um�L���#e:��G۷7޺�hbV���j6!r�y�W�</���Z��f��+����W(دH��um&�n�٠G���A��cJU�����/"
�88�e�]���` ���-s(�r�!�k�Pl�o���^�M�� ���n/Y��S�>��4��?�nl~Z	����"=���뙇�"{~T��0�f ~����#]�@:0�"49����=
�P}&�h�H��]B�Js�ߵw�V�f�BI,Oܧ!ŀ��Տ��!$�n��2U�+2B��a���U[��Z��t�;ՆM6mւ0ō��8��ئ)��*$x+e)Ёd)vE/K��t6��#,�"���͘�"ZL����o9��3ů�l�!�<�"���%er����Y}x�_C�S ?Hb ����L�U���������%�0�\�ؾlC}��|g�@H��Wπy����'	y��G����fKl
�Yj���NT~�3�6�	0��I�Ni��l�.}��n�K�����B�a^�6;`��t��[�SL�9�1��$Iն2��q�b~��&�A�3|듮hS�����������a�M����a�i����і]2��>_	��ٞ��5�!O	PS�^qtZ����G�N��X�A�^�7�4�#�hv�-��+��^��J� L8Os��;��%_=7� _��`�������THf;������yI��#�-�B�����ċQ�e:���Ri^h芆ș���A�ҡ���B]���=�ug�9��(��Q�����Ж�'��6�H�K[U��l�0$`	�+�!������W���Xh�s�fjBE�P.6�>����B#n�~��a�udq�)
�\�X��FKqp;����6?7HN�1^���+ @���4%,�y���-f�l�C�QSKVK_��|�*�)������H<��~��c�u�p�H��Ĵ�v�I,-z��͋P��@����Z�h�qS�!ԅG�"�L�vW�z��.�������_���`��/�_�����x���'��jc�6��`֨��T%&�//�`!�쨽�[���>IS�8	���u��6Մ��b�ɦ�����U�'�����m�h�j�/n�C �����LC��%bR������3��>p�3]?F��nu2�C� [AE�륄��总Q��H��8oJ�0.G�1�)f��I(��Tw�ܘ���+�e�n�NX��9%R���㕷y���BQ�c�(�-4�u�+8�2��C��Eb�M9�:�&��HΘ4�_]� 4��Fpl�ˑ�9T�,!�ߑXk��7ط'��
-3%g�O�n����[g�vb��(?�̍�����i�9!�]_�Aڢ�϶�z/����E/ӟ��ݽ��X�׆����e�sk��di���a8Yb��%#�k�-7�7�l8	��Q�����V��b<��1��p�:P�B?��25r�в憣�l٦��[�1p���ii��ZK|з[,�8��R^
�k}0���v�$�/�<c�r|�X:&yz�s�C��Π�L��e@祙>�Nz�1f��N9yu�!�
��dH�\S�h��{�dB�'�X+����R�V��P3�����ڬ�b�+G���~�׽�"=)T��2�|��\�XL>�;�|cf3�i,�f����>O�����T:�=M�Q׫�H���"]GU��8�:�&@����j*錋���%��������+%g0�{!|p�4!}�a�Qq@�S>�^fDC�d܅���PTC�h9ii���D�y�49�^��,����3��)+�����bA�͎<1k[��.ލ��K]�ѕg���F�o�o���TѠ?�]B��xY���E�e�E�.Dqi�������V�$,0ѧ�%8�����_f����~:���&��-��N\�9�l��zl��=k>N-����c����r%��7�v}���� ���k['�<듕X����� ������iZd�:z�z#�]��TEB�	�v�s��a��!.E��{ ɑ3&�k%�u� ��D��~/��Z����!�v�����Iͺ+��*�zB��x�k��5g�[�W�:�/��~�p�G�.yf�A�]ˇ��W���j>x�&A����b֜��5�ޤ� �EU\	��PPp�,�X��M�+�f�2o�J̺]��-I�l��r�$�k_<z�*����ˎV��n[�";Цo:n�N��Y����Ϭ�BP�}B]j,
@�V�jD'����ar�^��༭�4J �ǈ��EdC��[�2��V����_�96���%B�����t�Y�hFy�Q�^����(͌O�a�� ���?�|����c4"��1	��30{��!�ȫ�40MZ�4(B���>�3=$Q�S�c���u`2�l��Һ, +/�[�H�=��	o)��JfLڧ����j�e
�J����Q��sי�ǻ�3V�9nvʎk� S�(ͣ�AG��n�{�>��U���V'B>zc:\v��6�[ǭ��qTN��^Ucм �-ٌ���� Yz�l�{����~����{A�3S�.�1��r5�w2jl�����]������t�z c��F���gmV[AkBŀ������G��
���s�XS�<\�W�֧��vtcȎI*X��e�=�����Y�9�9s������B��@�i���nO�8�Y?�:ﱀ�k2������7�Ͱ4U"ס5L��$6 ���]ܖ�D��@n���?���G���L����pkmi���;�? <.��Lx�ȏ��H�Ι*�`�j���_#��"+ ��f������hO���4�t	l�!�?�N�Z ��A<��l��8V6�z�;�y[��Y�\�I�[DA*�4d��9F�Ky཈ ��m�8�1qt��@j	!]��sQ<ۡ�ؾ��.N�bkfɍ>���ʹ';#{]��z�;�=g=���t��B:uξD������>g��p��2��6|����Ӧ4$���9 ��L�'�K���Kg�e����?�􌏤_��蹇hd#��0a�/���J��.c�R��У�Ȼx�����X2��Q�0��������Z���i,f���n2���굸4+DC��G7����K�/���&�A��ޕs }���������L��۷9Z*��2�^�
��Ǖ����M2n�<E��
x�t�@L��Q�8�l�U ,�R�~q6����A�0!���� ����r���(��t����5�J(���X��Ω;8q��� 1����#�D���TJo�O�l�uGsͧB!��1���-����p�D֨�E�<2�]X��ok�&�����#9d������1{B^q���ڽl�M�V��H��Y�0��l�h�F�;���ș\��r�1�s�V��6o�����1�"�T�튜�C�-��$q�\V� 0l�+c�Ѐ���1�ܤH���d��j�h�jx���:��m�?�^Liޖ@[���w��	T�ROM�3K}�@���}�O�e2S�6QC����*kԬZ���n>��??)����}�S_u�,ދX�Ƀ��K�g*z18� �� ww�Sj �/(��H�9�^	��Xξ�?�O�~���G��ǖ���0� R^2x��y��;j�!�i��Ӏt��5y�@p�T���Y�J�_�Cz��m_=�~(�_�r����O8��n��RD��0C^�~��fu�P���$��p�G��j:�v���z�l�3wyڕP�~�߀��j�X���&׀PP��r3WDыZ�v2߶�̯XpP�������*��߶�k��b��n:=~˗w9C��߱T�A��/5so!�8���L���=i�$���A����}�{�#�N�@�;c��O��_�ʈʎ�r>�8�8Y޸	f�-N�G�MׄP\�,�<0�b)��J����6�+�N',��s���'�r���˻e��.���
�+���i*����o��n��S�:l4Lp�9�!#~]�x�����:��]u?���Es"E���ް��m�6ihfz��x���qў]��=M��'iO�@�T���&�<B �N3�^���x��v^���4c߱��t>���e�3�����.�	: N�f�� �x�k�%��l���-	~(��$�Ɨ�+X���l��'ptB�Zf1�=��z�=U��[�uǒ9��`�1F��d�e{::s�<�=�������?Gk�w4���KgPk�4R���Z0x��V]��2 ] ����@��J��(�H���L!��V�VS U/�����Ԉ%�r��B��t�{�i�I��!N�H��M��^>!d�I�aUԲ�q��@9�䜖������ʣKS�L3��(q���<��OkM�M�Hh.M���8:�t:d8�$���W&Ӏ�^#*�OMa�މ�<h7m�`Ƚ��V�/�E����l���R���ҡUS�~�\���y��a����h���P~8�n�=� ���%�Kg�<���Wz�$N�S m����EU�C����ɏ�V� ~.=��!21�©j�n~�������a0��M?�Y�$�Z�p"��`��ޚ]�>&���( pH��,_)yl����d�e[��@־;6�?R}�&�6���YɊ���^"��Ը����v:�t������m�`�=�15��P`(7�6�e����:!7�sQ�v;Է�Q����v �`|A_Tur5��꒥��Ƥ��v�3Pk+�&��{�	��j��ʾa�;b����#�8g*�3G�g�VS�\� CG��O�W��Y*������;� ��0�r.?FCj��il�#�3"��w�Ϡ�el����YU�}���`�kb�[n�A�$�/v�_���@�)���D�ǋ��^���&����Mx{�/�8	��KK�M�4�g�sS���u я�LU�S��PNf�I����q�!N���{�O����4s=,.�����,1j�`���8ϓ��N�sYo�Z�;\��=���݃�K��:�Eʭ��%�eA�\pRG/r|�3��+�ƏT���&���Ihh�q�;��S�EQrk�/��?!��	)y���k��[T��+<������9�Y14|Pŋ- t�T\�������XV�$��Q(�#�p�f��R"%�B �m�&#�`r���n�J��S.��+���f�ؐR�<vp0l�,��b��'������#��.l\>>�+ʼIӞ� E�\�8��)$�l#�OyUT�U������+k%�E����Ǉ�O1�`C�n��Ij�6�Fk[�a�?ǘ����G^�.s򤤖����W$Ӡ"��& �Z�G'�Ne���p�P��t��2�������&#M,Z��w �x�����{2�(����D������M�8Bt⹖�����d!L����X#qL�f�����+��Cr_���������Ԏi�U�M��1{�~ ���(_L�4w�S��[ˈ�2�DD�g8#���V�vB����zT�i��h�w�?��Rٳb���v�0�yt�z`Q���ćӸ�Ċr�V,��4�����˿�D(�_�'����Z����sJt&��gp��ִ�� ��E��m�N�T��=���V��k��Rfy�&C}|N@�����<HL��'GK�A�V��;��T�Wie��!
�Nn��kP��-������R�(:s��t�ghʃ��/����$�L|��
	�1R�i�[�@��e�+ �-z4��(."f�:���J�	����:F��A7���'a�0�k�yNe=�Б��xC2C�=א�Qn����勼؁�H�A���^��л:���kQ��Tt����2c�5nm�h
K�JPYM�L3��� �S\�7�K����`V��'Mv���˘�'�X̛��Һ���}{���+�="���L�͙}�+��$m
>@N�8�O�#�:��P>�m�_.Vߍ�Q"����Ѯ�+'���>=U?f�\�b��4�L] M��m1Š� d!�pf�5ԤƴaPy�`DX*����`�L����-��g�?���E��6au���PV�|rE�𤏜*z��N�^е�=��`^�ecs>�&��Ď���� ��P���	r[L뇒4q%p�ɐ�C�A��(�/����%�O�dG�9V�
m�x���� E�c�Q�arQ�AB����г�߲7�o=du��D"z���v�H:	� ��=]�i��4,���ڸ�ao�-�͊����?���&7g�x�I��V��F;\��)K'U�E3n�W��l�N�7_����Ñ��b���3�ˌ��1��GVG&(�J; L�s�^���Ф`�8�Ԩ�~'�A�?���Գ˱'0V�H_���	�F1�hÑ�*���OOC�tX��E$=:$��	LϸqeK)�إh��i�$k�&��z!��AJ5�x*�t! ��1�	>���1Z�&2f���H(���=9baua��+0�<ĲNE�_�N����G�Q��ҭꢓ�f�Q� �;�W��� �"5fL���'#/|�x�"6IY�D�>����,����!�u2_kh��_P��S
O_��M��3N2�|��Q�\�K��ʮ��p�}�C��"���b�s�r�gp�j�eq*.Pm�Ț�B�(��!�<Ȉ�!y䤢�����N�g�y&�t����)T��Uz��¼�g9��,J�,7b@&o���H��́|E)x>8�u�:E����kӖ����=1q�]�\��Vф�W "�W�qLA�}X����rנ��4���y?sN�`�&T7%��+�|M1} "}q��T"��^�i�f!�����r��e��#��i�85�����ѩ�U�<�tAdON�������rL����C��G�k�7�Q��,��*����|�9���;�>��IQ�<3����a.<�ɜVH���w��������יA9ih�v׎��/n|�l�������{�a�������l4����¼�gi����_�>�(�<�F(.��3��k��E�A'�Kt��C-����^'z'��@�I8/�'��@+�_�7����5�S�iL%ou;B���
TX�����r.�_P>�}����?Hy.�&�,���^���-j�()F����d�$ת��dP�@��8�5XF�q��Q02��.��HC,y%Qww�`����kd����=��B��?�v8�%�W}�f�M��S��iW(ťHWJ����>m{�g��{l9�L�O��̨Wm��wƃ��h�M���:L� �R2�xHm�_�O�+��5[F*k �q����sS�ۿ�J6�E�\3�2|�%F�WH{8��w�7.E�ɦ|�q��=� �׈�?�p���8Ĝ�B��W��Q;Hsb��U�]��y���p���a6��>��.�t\���#����ƕ�Y�Z�ŕ�~U��`Q1����\��t���TA�1�f�Zn#��*�����_�x�]2������,���˞��E���i0i��m�m�ߧ�e�"�N�:��@��`� r�R���Gh�K��x5u)��8DaUrR�����
�fRyC�g*��H��E�@��PD�Kz��	���l���허�G���A�P'f�,��jd�Q�G�M��t#�s�N�Lx�b��؈�G���_�ugQ�|�[n=��;�qpߓ�ձ����2t� V��@�頚o�.ào��WM��3$|-�Z�� ��.��?R�V�]ɧ3p�Si��*�YW��ʘ���;�;\�2X����Q��B�O+̭OA
�[����E���UP?��P��Wl۴�\�q~�.�ȑ�j��H���v��B�@#�i�A(�P��3>��(s�N�(�S���0e���0�k�����C���[��i��`�Y����U���:�c�:�,��F1���%�wYIr�����/���Í�J[�%j�C!���U�4��M{xi��$j{ޡN��d�zo���DB�&9��c�e�ZW�;�(���[��GkN�I�]�v��(�J�p��"Gc��%ɇ\�����_�����6{�p�+ډ4���אD�y0�c ��0� �W.F �����S��_�w����f7�J����A���ѝ�o�������/�Ӝ��]���0o�i������,V�f _~���l�?���֥��B�ջf�>v��S�ԧ��ʞ��2(�u�/�dr��QE1ک6u0.|��]2�.Xu9� �Kq)�L/�`'F���떦�.Q����K(�[&Y&�Xh>�Qw3���̽X�2
�BkO��u!	�C�/V��q��&y��-9jq�޺C( '~���!F�2i���;�{Y�g��䃪O��ݓנ��%��?nxՐ���(��|y���;��[��x���X�|�*��+��습~�i���e7W�I?�0�T���p��v��8�<�w���H�$���l:R�2H����KQ�MH~���T~~�\O��`�u�i\����$���%�%�QuYK�=�>�w8�,�qJY�9�b�9�<%���-~�dF���%�s�z�f�õ�@��GY�u��x���&fQ���47�!�'�p4JVx���{X�ރ�pA�����{�]��R.��T �f+
{�/ɧ�p��k�k�B���8��D
S� %z<��p²�L�Q0J�7�x�����}��Alm�ǵ�����:���1��&A�,I���dQ\�L���]6uc��=�4i3� \����
���ozc�7���*̽'��״>܉#;KuU��fa/���T-�	�D��� �ҫ�"���D�륒{��&��3͸'���.�� �`�EG�D0�P�PN�sEU��2�&�$�������� ZX�l��s��ǽXČj�8=�E�����{�8m"�,F[pb\A!'bI�U|0	(�R4�����[�8�p�ʜu����Z{�_6/��n�>��ZG���y���%7κ�'�=v�D��z�3]c���$�]�D6m�Y�|����VTr��oB,�n6]R�Fssae�q�NC�]��mr�]G� �ҝN�ר��	�i˕^g�'���$��g��AX>ۗ��V�G���e�)}'��N�R�������۴��q��2�����Cl2�Y<-��2`��u�_xJ�Y�(�-���휹x��vƑ#7�� �j=�����+���ϔ�I�ۨI���ª�͕�N���7��FlS����e�i�[�2���g`tI�Cqg�Ƴ���(ڐ���P����`�5�f���B�Y�:���6*�W���HU4�\HC��Ta�'d�Up �Mx2��?:�?�X/B��G�-k@-s�)8uV*�Ι:�f&�*��c��c\G�;F!����Bf�������\ v�����UDu�b+�ޯdY���YL����u�+�vU��Bp0�I��V�+��nnU΀� ���_1<�Jp����'̕S`��8#�K �]�t�g�ݺ3ˡ榩on����k��c�m"�3o	H08��"��#� ���[��3;}��X���y�]�3'19F!�L�����|��e-�HI����[qz@>����
)]���F��=�~�]<�;�� ���K��._���S3����
]
�ܻ8:��B��1��7��x�ֿ��i��5h�D[ 4�CwǕ�����)5��B�des)n��(�����1�.��- '��6�@,��KS�U1a:9�Ǯ Sfhw?�f[!���M�g2t��9�}=�79Kf�&�ڪ�"��TXV��`�5xNmmFu�[�R{���q���4�&P]���&v�h�AK9|����o��M�5?&���iB}{�9O����x���]m[��S���at^I0`1��g|��\��q�>nb��S�ĭ�+K��M���
�#������~/,-^�e�s~���K4%Ewr$YYL"�a�j����C������4����˶[�	 ��.�FV�	&�ߑNK��ݳrY��W��e�."�t:黥�A$ߚ������;��=���vsW�Ғ��H������yO�nv�b�n���5�,��M����b%�m�� iT��ߒ�a�͸&S��ܔ�u@�֪_����LZ�z��i���,�,���21�E���v�r
�ֿ"wB��@�\����*s�nR�ۻ���0�9�S����ʿ�c2�/ç.m}�Q����$��x���%��x��c��F7?4=E�r9�!�}1	aP�]8�)���W�W�"�pa
�fo��hq�K��Z�걡�������;ީP�"Z��2�ٓ��{!([f���p������Ov8ȡ���u|���q�86�(��V��`{���}��˽�q�7��ʘ�����dH�Ǌ��+T�X<dI�~�q�,iɶq���Z��2^yM�����}�V���5If4�Х?�Yt������"��> vVX�ބp؍!��O19��?:��3"�*$F����/3�N.���π�FW�����6��ˎ�sS�ݟ/.���~N�����D@E �Z���hN�A�,�+�i_[��!H�Z�\Z�ɉ��D1յv:23�"#C�t���и�E*������y�D3����h�;�jpqךּRU �� ��v˲���y9�����Q����@�J-A8���> T�k�
0�F���!�c�"G�6!SM jQ��rO�
ʖ��+��^��)���?<3�R�v*���ai5�Li╏��	#),DdfG��k88�)G�R�!�N�/ Ms�+2R�$0���JQ��a�=��xn�筘�1�c��5)J��f$\G'�w��wjb��[��l��kr�?�%���'^����7��ΖxW��(7Oc ��P��H(� �n�6P3u 576r�9�3���U7GhtZR�(���=ƌa6	S���ѽי�_�\2�j-�u�|Jw�Lє�F�����]1���0��V잉X���6t�������U�3���PH���8�Ǡ�Ԡc����w�b4��� -ۖ�B%��� ��9jr����� 'ϸ>�f��Kd;Q}�Ct�qv�=��}.-�_�����g�Z�}��߂����R��%~�k?�פ�?&��`-!k�*��g�����4�T&e��^ы��ٽ�K���m��*	����:Scx-|��(�s��.~�*Y����k�����MuY#"S�KT=>h<:r��=
*7>K��'C��K_=��]����ԝ�!@��Y���U{R�������^ �f`�͵����ueR5�?���������6� ���3q�T��/� �����#����^�H��g9Ĵ�d���>�������|n=��;����H�n��~yC��o��Fr���^g�s뻞a�;�A��h%�YYM����`ި����J�]h\�O=B[{�~>�N�/wNį�qW1Y�GI#U}�����@��x֔�=�������ȋ��?�3#����IT�\߹��PYbq]+D�
������IHl�8�)t�9j�
�Aw$�0�ǌI?2�vu�{�����<��z�l�}f�!_tX�^|yB�mÀ��	��@�����8a;ڋ� ��,6wU��1��I�0E�����OdR��ח�5�i�C�%:pޚ&����GaYh{D�+37�ces�[���-�����0Än��I5];�Đ@֣Z#A[�߮�����Gsu��v���V�#�����5`��$�ۣ��� �6`vr�V���2>�%���Z]���@ղ>�&�1A�I �w�ѷy��^�w�V ��2_�dӷF�$�|���A#f8�?��ß�0�ڀ#@��ȯ\����6)��'T� �o�����qn|�|M�2������<�@���{j��-IS��l9{12JO�S�Jx�]��،�����x�r^����
V���vF���Z]2E�&�ڄ�Y˫9��{w��}t#*���
��Ń
4�>���P��� �5`N%�<BHS�:���aėR�U�F�P��.Xv#�8��!�
cn��"e_�@�b��*5���υ(����~m�"�E��X.�UA�Jb�Q��J�풉<�ά�&2�|+:�(��--H� ���9��)�}L!2؋7�;� �e��z�Z����渼�"7�''5D�1�ke�n�]Fx쌎��f�Q[˞RX�i>��<M�}��Ni�Ҵ#L��z��Nt�����#M�3��T�bhՆkb"=��5s����h߿��c��Μ�ąj��=qdH�N�%�l�x�A��Dϳ�4��?r	�����z�(�|�[���l ���<c�>�,F�jȰT�=ҁ��٪��t�S'1+{ϼҴ��T��hc\��܅`�ր�7�K}��*�t��g?�S�+��"���dS��L��⃧�� �_��zX>�W0���3���<~>�ڥ����#�4�ִ����shQ�6b��$-��������V�ʰ�a1��q9Ž2g	�ЖMŀ��ep8�ғK%LZ}�lX��l8�&�B�ܧ�%Y.�����L1\#w�_�k���zK�Bl�[�k�|dT�+�a0�ˀUfv���E0N~��D!�eT(��(9#��z�$V�S�3d�n�_��E(�ۗ����+�B���|O�5'�K-�;��g4�ړ�U�c� %a3��a�'B��`f������0\��C��x#�]}D�C'���qb��C��2�m��
H�5t}d�6���W�cH��Oە��\ؕiG���N�����+|$2�+�"5L9�$D[�a��:x(d.84D{�wew����I5�����#���2f�u����A��\I���,x����A=I��mp^Q��G�}�1����Џ�,h��.W�9rf�u���>A����� Ǉ��?�xB��'�}fl���)�9�JV#�Ak�sp�ƣ��U����y���C�0��E�d�[��
�YKT��p�i�.��҅�"�����'B���*v�V&�x_OeY^�N��}v$..*::�GN7��EO����q����ةPѲ����7�{��LKC�4*�1�h�̗�����\'�s�aU_���xA&��īdkr�Ld8��]0��"�(�]r��K��a�`�� ��S�)F9JS�B�b�1$8� L�%��}�Q�'h2G�qۤ�[{����I?Vs����{<i�֒�42�WC�2h#V+<Q��H�7y�=ܹǢ�M�N������l��L�A"�o���\+���0�n&F��vDN�!�2��g�6M4������wO�D}Ӣ�s4w��A��F�?�,i��I��7�
�9ÍH���K�cb+?.?��Z0�vk�g�����*k�-f�oWhw��i�_,q���H��j؀�`&P�/jCy�w�\?�d�B���@�q�������J7�SP���e����v	�J[�FK�>A׌�2�cwY>P������n+#����d�� �h�e��s�ֲ�{rʺ`e�ed�ͣ�GN��u���:Q���c�)�(�}df�	��+e�	S��H&���X�.�}kԤD��RA�\̃��X��D6ۡ>0�Q��w�E��6#E)���]��[�%}�J�n�QRڥ1~�E4�=�1��6z��&�b΃ב<:�� �S4�g4a�GV�m$IN^V�`�!����_�n�{�=Ʃ��#��vz�v�In�����VI�	١^4�!��9?K��%��b#c�yQ�T>�b����������?YᣣI�MUZ5!�v[3������3�]wJ��|���S��(���N�
T<���ۏynYT�`�O�/���a�$�K���8��t+��#g~A��!�$B��wO�Ӷo&��7Q�~K�dX6+�¾��jD_��5���'>ʓۀ;�@_K[0"g��Fn��(����0b�b83�[�v3<����-�砃t��G~��QQR]*���J>��hԀ�\yQ��`[��K���F����<�8c���M�%�{����O�&�ex��Q�Ԉ]�ӴoG/Yg�aIL��!(��tV^Cu���F�n~�5�SK<CT�D����2�HHJZ�Wn?�vּ��� �^�����iI�n|���wߕ��,�/�:W�-��zM}��_YAxC��5���h���;y���@�����{V`K�4��Ni��5G�������ɖKrAd�|�X�꟬��a�C�����u�EkPmt�jZv�� �F�_��������DI����<����-
�ɭ�J�n
EV���tW�V�^�Aw>��pfk��-���E
��J�Ǭ��@���3b����B�6��밟^�P=��_��`'��k���\�-.��j�&v5Un���ȱ���XJ�e�p�E�Ͳ�s��~�B��!����QL'2�e��nT����ε��M��Ե���b��mUW��FI'!�H�dk͌$���*a�hT�4E.M<�7*����qH��L~����o� �I��q�	��D�z_��g1��^�$H�VWU/l?�� Q�}ᜋ@�S�����B���q7�D���b�|� �^4wv@��I<?RN% �8E�\����P�9�.�@�hr�$ݫD��'�t�B:��Mh�ͣT�ʾ���=t�9]q�sᒓ�|��j!8gA�>�)]P�j�>���X�~����x�ͥ�(_�fڃ�z��
��8*7�a���8��jՂ��,c�wY���$���ber��F�C�c]����MƸ�oI���L�o+�<X�Q{���(ڹ�u��]���>�4ә;�o?&<{�)VVr��M��t��2R�t*vS�w�5m{ P�Ϋ�b��xcJ3P#����1S;�c�ү�#�5W�����xeo0ʲ��l���ӊ����w��$#
ț㐄5�B�3h%���
<Y]]�a�vHg�D�^�kB��͕۸RZu��C]�!��HL9��?��2 �P���\E�j� ��~�sM�,Q������^�{d�D��M�D�]B�/q��E����P'�z�����e:�#4C��JO�ӊH� @Y[Q��%x�c4T�.G�C�&�m�M<��*ǒ���h�;�:�Z���h������Tc)р�����ڍ]���2	Yrf*fN�{m$�O��8��{�}
���+��j�
�:�a�P��~ֿ����v�rZ�F�t�:����D��f}b�:�����|���{�nS�f�Q�̣xW+
E~{`��ć���RD�� �z���k�$g�W��-,�c�V��n������	;�m7�LwJ+I�z,9Z �^�~�Z��v�o*ƜS�sܕ֚�b�Cxif����j1Ep��I��t�B���Wy=��ږ�]�=@iH�ū�4*I�2ص�n�
�1�� JSm��b��XM!bn��h]��V5d�?�\d;]Ńj�ml�$U��z���Đ�7A�,�<�̅Vzr���gV�IgR�:�� $n<��F/¶����ڶh/�]02�T����U�w�StǨ�<I煺���*�KOӿ�������Mڸ�e&؛�0�	�|MQpc㾕�(�e�4�P�֋(��B���q������T�nj�@l���R�5��EV�r�`�4ID{��?+��[oɛo�EX�codǉ�����ph���Ĩ+Z/���D~���;�R�0�/��v��@J���9�vU����W�/�Oel!uY��"������ؽ�m�� �����vFXR{2�܋��<Ӽ����dw����G:�)('��f���\6�-������4�^�����Z�4�#.<���(�xG��Z��G_�V�<��=��rJ+�'K/=�t�,(��r[Q0�gH�׺�@�r:�x�������G/��u�8�V+p��Q�c���UR1}*�:�Q�	2.�r\O�̴]5��O��YI�!��oI	����M(zJލ
��۱��M�S�>��Fy�QFr�4��S�'��?��P� $+�Ɂ��מ,.�b��~J��\W'%�D0�խT��"s�'��P��R�c����@y�xF��-�#1�n�(GI�d\l�{+Б$����*VO�*��f�9u�%�$� XGw�?\"��a�ZN3���62&��W��V^C��s^�Q)���#o;_��L��Ԟ/M�?��nQ8Zit�p�R�wkHǽ���Ώ�%�1����p�|o�4S��K��t��j�Ŷ�S����Ѥ�����A����p
�\Dq&!-�i���ݡi�a2OE��W�b������ZM�
�ෂlG�"5[��M�,jX��S������a+��l��qH���ᒰVM˒��R��g�5K��nH�/�u]G��6d�*��'Ɋ��+#�۸t�4���p���҆��q������T�;|���l���>w:�a���R�v��]���>|�rI,a&�͠��]�&1ݫ�l��,�t���z�k�@_$�t��V�\*��ح�}rÑ��w�wJ�]!����)���v��G[� �/�떲R @S���iO}��ڹv]"�b|+�<�k8s|s�Ui�H���ߕ=�c���ZB����@5,E;��H�Q���i(U9	,ž<=�	�6��s� x��D>�T,��J<ӆ2ɠ�P���6�C���� 2L���Ab��J���Sͅ�r�!�����V�.�ov�����q�7�W'���ʀ����}N]R�l����y��kQa�uG8�n�n�l��>)����\�|�'��b����2��� 4���>����^�##�T�$K����	�h�OkC<�br�h�Áu�$��"����3P���24��n�do6�K��?��	���J�
JG�)�ec�V�,G"�Mы�WiF5�.~�];{�c%t����G�#W����u�[��s��}>��B�����^#"�g_�w~c���1u��|/�f�HdO�EWd��Am��MIТkK���z�L�w�6ҔQ�M C���A$�O�hh���
S�Ϛތ�����*�d���U>�C�Wj��ܩL��Ny%z}*?@�܈��d�#��T.�gCq� Ps�	#��?��(A}�0h�]]}��������s�,�bU0Y}S�xV��f���:��	�fK6K�G�ԑf�s(���%gÅ�f�ZO���y��*��r��+���^�%~6!���z��D�B����㌘�'��K��ϲl�=�x}�\N����t���݇�0�D��naA�h�o��[O������y�\ ��^ہ��"$���/�����Z�p��j��܇��j�D�bJs��If���B�vK�B���]���;��m`3VK����R$�V m�J���d?7����~��W����Z:3FX�Tk��a���/�e|�1g�K�Za��@�D�n���V��ު����1�a�\�X��SQ��� �I�=��OlޡŬ�p��W�g1}qF}¬ұ�k����o�W�z���br��^��U˱cǌnf$�v�������$�`Dh�+3oPʬ/��e��z-��.����Ǹg�ԽY���n��~)��� ੼<˙�hӶ��D@��fT��R'�"�8�Kщ:JM���KG�Q�� �-��ُ�Q�J>�:8�k��xn� #령(����P�Ǥl�XI��
���ܒ'O���<�I��e<G�)�P!��.��9���~��뒵u��rP�]���������[)�K_��H�ly���?:6���8f�r��9.�;��S�M�:�h�R&�����(��v$l���5S����P	��_|]��ѕ���"�M�:��'�E�b{�J�?�Э2�ŭ+*[�*��ێOs|�|��ʱ31�ƚ�\���s ��
�f%���`�y�!<^HW]�㽬U�C�0~�1VݰV@aGI��୙iȁ@t��G)��jr$%�H�n�W 8�u��l)Q ������2責�y%(^� ���L.[b��Z�kn��3�b�4���#�̸�B,.��dFRNG9��s4[�W�hdϵ�d�X�[Jx�����q��cǛ6�[��%=�j�-�M	�?�� E;��Y���$x=i(3��,������$����������{���SGU�[*?���x����m�3��M㬹+I�d+�09�z�k�'���}bbf�6Β��y���
#��\˘rC���"��sӕ�n��L��3��I��J�k����#��M�!x[Ssb�,n��x�)����*���b�+�����(J�E�.O/wG5���,E��Kgd9�,��������vj�Z�H�\I�	�̠�d�$�X>��_���h�}���<|^���s�6�ve�^�7#��YOe�d\b�L�K�H#\0�� �Ҵ�w c߅�eN�A��PxP�Κ�ԟ�Z��ɂ0̺1]ƛ���kFN�
#��'0iu�&!�����	�W����V�e���-��be]VŲ`���S=�m�m�H'�f4[�����,Y���|}5%W�â�B���Vd�;�%ܚD!C�p��E���&w��O�t ��"~� �*�Rg^�do���ʓrG�IRh<4����9�ߌ���4��%U��RT�@a{�%M�Ee/��`���ȝ���t�d��WC뫪W��U�Q��j#ў�6X_��|^�]�t�0Y�^@�V F*�DK׾L��)m�I�k�4j�B�
�������(��~҉�9��t\��������R�r
:s�e U$^A��8�owҧ��2���#os�}�|��6�v�Ş%J��M��ͺw�j��s��"�J��qF��������38"Ƚ���8,P�r�]��H���03�[)��'e�,�<��Q�3�:��	L�y���`r���z�?)U��@U��>�
�׹ ��J���V��
��1n�M�9i���YGF�~�<I���& �V6V��
�6��,�p��X���".c=�$��t�d\O��h�tW�S��<�>'c������x=�� �����Sd���/ժڛաy�E�f����U�;J�W仄6ԇ$f/����\(�\�pՇV_T�a�Ɵ��K;(�Ws�g6P�
�:�Qn��v��X�-���A��<���\C��_~�l��-�X������Y�һzu<q>�9�P� ��p����{�y�z��:z��bX�n@_Z��2��Ev���W�F�Z �F"��*��7�/�w��W�M�����)�R���[M23�d��xe�.S�bI��8*�:�4�V!���kf����g]N������y���c����.MGiU�M5#G}����t��ֽ���ZK��a���usp�(�Z�eu�GmL5v0�]�(206{���I7��sZ�x�z�Щk�y��A��l.��
e��i���G��z�᜖���'	�1Z�U{�ݻ����*�.b��
1\��廐���T�QDB�V;��*a?�Ue�26c�14�L��`�[Y#w��m���7�S���=�l'��'d\�`Hyݼ��H��"ќb(:�>��tv�0i}1��qS60"��o��ߜR?��ƵE��ʼ�Tgq�,��p�Bxu�f-�+Y�n�qo{�o��zo��]R�U\{x��ΚxY�~�����)�Ә�Z�<E,a�9���7Ɋ�β� �M.���zQ?Ң}<(���7�&,c�!��(���5�CZ �����x1����O�q�?���ŚF�Y�eɂ�����bSο`n�w@�|�,�M+ #��_�Jݲk탄F)�]� ���uy�F��de��?|�l �����Q������E3R!���]A�1��%ى!��2^��+oݦ�W��w��(�qtf��EZp�Ϊ���C&�ꄆ�O|��9\�:�}�7�tA�^e3��[�wV���w��$�ԑͭ�q���FU�a���Ste ��8$�.�#�<a;}�-4���ųy�Ɲ�YR����:ܢ���~�2��'}�Z8�IW�y�BA샥�Ɯ�?mY�A��Aę��,��D/ils��N��5f5RP0-
K��;�"���˂p�Y��@$��4�p}\nV��Ú߿�F9To�槰�Th���G����V`:�&9o�0�a�E�[�����P)��u����E^��w�����
z>�:>��`-ݩ�-~˴]`p����j�?�=��ptx*&���b�r�*�����ݔ�{G�_a�	܎������ ��M�>$>��Ӫl����$�y)>��w=��l�XB����0[ˠ����=�ݬ6����i���RQ�]�\q��=ǡ<�"�����hhR~���P,tkd�ȚY��IF���d{1���O��'̷3]^���[���~���		� ��S�s�PE��`e<+fu!dy&Z�A��E�L񍔷���pp��|��܃���8�!~��7�S�? ��j�[��N3+��L��:@�4z�;$
w�5s�ٳ��dˍ�
Qf.WD��D\��<�11e"�0G@W��c�A�P����͹�h�8.���T����bZ��訿����&¼��ۦ��6��k�BNd��3��[n�����D&I{s�����î��ߋp�Z.�
��`�۲�߬����=#?���L�N��k���
��5WS�;��u4O�y��8���I!E���<����`y�l�G���+p��4;X��=��ܩI��\�TP����8��ۙX���al�%,Ʋ��{��I� C�\=�3;��+�crm�e^����{QQΒ�����Γ���)U�K
OL��L �f3������ƥ+�S
���<�)�hq���~,�1��Co�&��3QI��ye�?�;�V���#�8m2$�<��{��?a�NT����,x��³�
�熃�?	rS���J��/"��t���u�GP ��v��
�A�{�|LX�FE3����vi�m��ڪ��������`%��p�ɛ��0N�v�Y��%�'��Ie�GB��m���;�8�=���I�\1����;�GU��M��k=7�����s�J؈�j�ǥ0��R�'i���븪\�%�Z��c-y�	ۏ�0�F����f�,�&�o��s����D�&��40~�y����#{�#�RD�8""��
�>8Ց�Yҡ����R���<����R�-�w�1ꮭ�}K���dC��k�'��a��s�ll�8�E&�}��'넺�v�����l�<U�]�6قo�K�(�Fjz�	z����S�upöo�1�m�Z؄'��n�YV�ɒ̕��#G|(�$���Ti �(�I�t���J���1��=@�Ee��[���BwKb(��}>�x��g�9n��X��i�����2�N6��`����*���o�$5*f'��/�e߰,D����mG�6�Ϩ �B^·��bb�hdt��e���e���d��C����I������w��B�E2dz	B�ݯF>rG���ⷣ`�3���%ib4P� PR�z���ʯ6U���b�Ps���oU�l��yd ,3����g�7���ݳ��GHd�RÎ�%nZ����{:P��:殭۩P�pQ��u#��lc!���#��oP>{>��#�ώ%�qS#ݨ�!�k�o��s/Ч_7�9P�3|y#��Ѷ\��CA��f��'���-����*,����ivb����E��j���C`�,��J���K.���N��>Dj}� �"��fmP��\o^SI����m9�}-�,�����Ơ������3���4�8��~�F�6�$��&DnF^�������*��y�b�ޡA
��-��ذ5&��3�<����i_�����j�LE �&����i����R�U�'���ρݱ3?�Is+���[=�m�k�ئ��8a��'�^NTd�~R��.)F.��:[�@�����Q�Q>�f�qY<������#�+���W�������[v]̵R�ih<��k�+^���m�ձ��ߚ��G*y=@\f}���:�K}��z7���E$XQ��J�]�M7��ze<����C��ѯL_L����[��/��/4`2�2�M��@�o_�P����0�k�na.9���j�U���nZf�} =*�d/�v��ͨ�T4�3�d%��w�J_���+�Ζ~��H��HA"�(���n�-FZ�w"�?}����C���⌅6QlG�x��1��q�{5J[ڕ�AځNIh\��r�
r�>o\���at7�"I=���2ɜ�z�
'�������E�I
c�$e% ɉ��ʲ�Ϸ�,d�F2����iB=��<Sek��#H��d�7?g����lUe��!����"�pTS[��!L���s�\��޻u7�� �{���+��ԯ�M ��Do�|$�KZ�ֵ��P��Ѽ�dyj� O�B�}?m;�l	 �`k��b���F��3;����S�vMl�V0���8�vdg".��K�e#���('��I7���݆]X�3�?	�vt����o,_�k;7�Ј�n�Wic����O*��L�����S i9����t��W��I�UR���5e8������dY]��	�k�u5��5�oWY$��*y]�+wm�]'&�Oe�o���bu\����������+b�>yQs��;��]��N��=��6t*V��ඝ��Ҩ���6�l��;A0��#/����,��Ψm=j���1���D�A�RP5�qhsbVCm�_�zn~��sU޻ ��-a�{D�5~���%�B|ﷵڏ!a�:�Tic<2����K�D�H�ΫT��8ޒP�4�1�1y\��S�5O08�WYNL"#��Y)�������J�������d|/\^�����7l����v 7�X�w���������s\���ke0��.�QeX����	5���4,�+y��ѷ�I;�9�Ν�4���v��)�|���T�Œ�Gt��;&���yGO0E���f�R�O�zS�Դ����c����T���=�����R&����Y�O����$�VT_I+�Ԫ���b.	��=!c�0'r�7e��_3��R�c#@�(�rmc��`���4N�����v2y*�* ��l�C�\^괳���n�<!��}����h��v"9�љ�<1o�t1��)qj&r���F�}A������
h�)�)����+�S�H��a����gc���zpHi���.@�J���lgI���`��z�b\>��~Y �2��̖a�H��I���T����LO��{�<<*ړ��5�>b��Լ̯0�̤)�v�bCW�"�B���+]O }8�H-Y�֨�K�X��j�h�IS=ቓ��)�V!��wf.�dqt�/����e V���������n��ɡ�C��ųn�<mFK�a
�<z�	z�0+`cTN%���z:��'�ª>��Ij��QJ�B@��ю�2.��i��]���$O&
�д���N�ė�r���)�u�C����1>@��y��)?�b*��ʍ���e�~hM?|�F,@RE1n�лgA���ͳO53�L�Q�1��9�~�f�꬘�B@��/�Ƙ��M��kUҼ�T�kƼ��j݅)�1&�����V�����`����n�E�P����ZA����N����L��p��`���c��Db�]q7�U�?l�+S��^ƼSIIn��i���rb��6,����7��ȳ)?> c�Gr��&�l��6oQ�rչ�l��^e
�Y �ֱ��3�g�U}u�b)�}u
T�e��~k <����a�D+Νj�+t!��$=J�e���7ɀ�A⮱��;�Iq�~h���w���4�;��ܧ��Hz��������6-o)o�=
�Q����� ��×�'�iG�4��йmHb�?F� ]�Z�[;<��ʰ�L���UBg6T�ϛ�TX×��
5^Ցm�	zt��
/u�*�m�v�2����ų�`�k
��L��k��-뗱ǯ#���4a��w�e^�g�@$��|hlUH�
g��$������P+��{�		��~���b<B��M�d���j!eq�86=���!ɂ?��X���v����o�!�/q��msλ���{�`g�UH�fGI옵�~M�>	S��D�Uq�.h@)z���?U�n���,������oЁG�pR%��k��YM�[�����|�X���T2�ݝ� ������M53n|��K�.f�
ڱδK��ȶ����s���q��r�@�x�x�9[�TV=�SW\����U��!�시�{|��\�(��F�%)��2�U�]r&�.��pR4-L�"�S�� ���n�\��^���~QBC����hV�ҿ�\�>$k���Tu���K�τr=D����\��o{:��#�x1v����!����%�9u���������9�n����$F��_i��
����(gߨ9���6�ho�j��)�Ǿv��0���a���q�j�Z��a�@��\|Y����z���ԓ���W�J'��F�-���d^V�А1D{1���&m���=9BNe��`�{�7gs7"�d���D\UX�݄_p�X�!�������e@!V�t�n�@#W84�_����?�8ldc{H�e,L6Wuz����x��Ũ��K�c!/�"J��� z���*ϐ"##�e�.�0��*@u*7��LR~q6(�ʸ�|*�O�;��}j��!�����D'��1�T��'�|.ڣ[ �����XǤ�����<T |o�m �+��"�n:�$�N{���]�����x�o&T�V�G�� ��U�c�I�̔꾬֧��� ڳ	:N��e���'��� �b�
��'��C(��Ȩܞ(} �;D�7iaIO���s�;�3�	ST�s��,H��.D<f)e0G$!��zL��4���[��l*͆����St��аw��o����m�x�����["�)�a��~��5����`߿EmN�,b�.W%�=xQ���� �X���$YX���p��!�H����N���3���$}��#���o�0Q~0LN.�0���뻗ۍ��n����S���]�㱾�qVu5�<׈K�C��-S)�#�{�'z ��!�I�$�D���籖7*�h���@Ƴ�GYE3�Z�ӱy�
w�ooO$Љ���xa�c�@�]?郆��=7lF1��"��3�J��޽�G��o:�C�L���Y��d� '�uX3��eW�����q�d��Q���;��ɳ����p�4��њr���#`|�(�� ���L���k��g�G�1����{���^=��n"�0�e���ܨ���yb��d(����Y����v�׹2�:���
"k�h�n���Ғ�&:��W$J��t��6՛��߬�\m��5�_ΐ�R��u@��{�n�C]<h����dN���^���Q^��[�>&�*�r��~^ɽ*��g��,��@�Wu�8�θ��j�4,O5�a�����:bsxb��C�,�}(!(X������Z[����Ҥ�oO���K+��!���W��At��|ȇ�-��Ūfw�o,@��T����3��.�����O�I����:^�U�a�H�ꨙ��
��u~�OO��YC��Ƞ�*���h@}�y��?��ښ%�.��ʈ�1r����6P�j՜����[�̧��C�ũǶu�dx�S���]��]�QÊ:$c����Nv���L`JE�s�L_��?䧟�%�~��5s�[NW�od��\z�GU�&E\bpk\�*�$K�xF�d3�(�TK#���<ѹ����na1���-�h��Ly���Hk��23�'q��Pa�Q_7�X>�C
o��Wt�����YO1:#�{MHa�}r�������n�0t�>��k^[�8��L����_��Cߩ"`#���tƻ 0������
oY�%�;��*jAF��>�@ ռ9�K!�O�7��1�~ä�%O)��'	Z�ù�}B�k�<����@�h>����J�-�pSm<>��#�C�a�R������|���jP]��<�gU*�\T3K�8qX���Nyǹ���ŜD6YGDCm�sCIKhmB�T��TD@��֐�h�����N�[��%�9�֐�r�o-��~% mAԵ�*���p�E����p@P�[�kX�P��g����9,S͝��P^u��#�R����>�
�:m���}?-�v�@��2� u�i��s��� ��~\;���K!����*�ߦ�V�4���w>��#|�QȊ��`UG*7:�zaӶu�^���P�!�RX�Q�����@J�yH��TN���X�yF�ln��'�n\���L��u�o�
q4��Nl�+��9��������ZD��w��h�'\I�G_�G��h���̩������6_+#�p�l�΅3�M���8�sP���Q�}&�+7O��i���~����N�ƣB����znLce��U^Q5�Q��yH�w�u����Lj���J8G�WM��;R�}?�z-�O|Q��n����}��6�P��;�y���:�+���[E�=�e
n�D�����ut����*5��w����v