��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�!��
��%Y l�׾����|R�bD�E���y"���7�cZ��T�1��I���̲4
 �����h����N�b7�{P��B-ş�y��jҹj���p�&�x4��r��~�������>�.�����d����H2��(�{�At�8��D>\�?}���*�~+�䣡M1�����)H�+�҅6T�����В���^F~k�W>1Z�fzi\�+��IQ�d�i��F�1[��GH8θ�1��2����lq~�������G)߲.�����zև�b
2�몫���W7�m+V+���4�$j��@3̗��"%�Z=�dY�Ή�|�'
�x����9�n������n�0�y�$�����p���z��:� S���2J��؀b��5pt��{�	�\U�Fn�,�x�1��sE7gZ)�t"�ΗUE��F��ޛ��bQg,�~c&$ ��_����
�}4<+h*U��BqG���hK�;N�_'7g������\�(� �OJ'�`Ƃ�S�U��P�XO������O�F�I��>p���}�7���j>[S�=]����=vK�ڲ�f=fп�B�Gg�-T���4�G�,;��i�F�Q���?�bv�X/�׊\���Y;�j���Rd����l #�	!������3�f�s�'�Lx��l��N��m���z�)Ѭq��4�d���%�S��y!�������9ٜĆ�N��fV��n/^����u���Ԣ|����ig�����w���\�`��,�|]� o[��Cd�-N;{�:�3�[
�v[��o86vj�>d!�"���]a26i}��'�m@�W��#��2s�r��W�%����ֵ@�*�����;�u�����״G^�]��E7qK���f��'GN���TI9j���n���*\����XGK��9�/v��?HS,���W�U���R���@�j�jM���?��X��W�&KD�Od�V:O���Z8a��}`
��
��vñ@jS��%"�=˪kw��Y�`AU,;/D��Q��w�X���1y�+R+^��o/m��n�$m������[#C}
�o�m=�9�\�U�nɗ���;�Z�����I��_����l���!�J����޳�[�����nT�9(%\-�D�p_��1���h�ā���U!~���SS���ԠPs1��ոw�o�[m%���0~LG��,NL�ow�� A�E�8�T�� h��	�2Il�/�a������_ӱ~��γ�ʃp���C�7�T��k#7uP�醐nTGmV��8_d4�Hd����ԃ"E��"5��w�R$�7B:6��{O�ς������kF=Z�N�B�@��+�a���b��\������R�����n<�O��7A�%%��#3��"��D�S�
����+ƹm���@K��w�r�񫓔���Dpg猑�DK<U�����_������Ѹ6��ണev����9��	��_����Uĕu���T���;kxŕ��!�D!T.�CD:J�F�)��!t1U��Y�`c�2�l�	1��?��: �;�%d�A���;'��,"�����[�,<��k�aؤވc�����bIc��=��p�7m�<���7)��4łL��OY�tdF���p��lTe79B��o/���������&e�xU��[���`�~©�,F��#��M��ODӅ����hڳ��F�T���7�!b��d��n:�~%���N�'ѪFKS�����|#��.����y�)�a�.�������P��.�K=�0�!/ڨB��H̳l�Xz�`���N��P�����sB&��]��/b��ܘb8���,`�_��p�^q}X"����?%x�͌-�i�"���'h�ֹ�+}��YpK�� q_\���g�@%4=ʃ`�^NY"�C ����`#������-�M4�e�����K��:6�����	�G2�y� S��i��'��~r\T\JӀ0�d_rIq0�lN7u�G��m7���f*�>!k��p~���?��m��U���y$S�8��'T�1����g�!�:Z[[f7*0J���!�|��H��U#�*��_	ڛ#b[z�Xw�#����������r���L^�6�(q4TWf�9�YV�0p������\�un`��6$B�ĩ��wO%�D���|��ao��L��nW^���ɲ���q�,U$��6�;o����|J.��D���=[o��.�ٻ`r�'o
�ݙ�=����R�u� ��5�%Sψ� �2fܲ�rw�k;7%v2�-R&�?k�&P��K�:C΍>�	����d������f��'�{���$k�iE�:!Sb�1l<��>J0���2�B�k�_�Y�D$׈WG|��_O_�^���j���*&�t�Nk/:?,�+d��P�;Wd��<���|�ɒzB����Wok���q�QF k�X������S/ԥ���LUԹӼ�:��Y�VS<~������'K�Md�!x�*�Cf�\�[J��X�7�ּ��S
3�t����~J�/���C�����0�����!_�+c�:��5�2�r����0��Iޜ�G���!�������m�KN^M#�!F�'�΄��Y�m�pj�̮f�7e������on�c/[��`�b�m�yZ��i�-f!�E�tN�b$z���EY� |��1�N�[��L��O|3�t�x�h(��K4���g�i�h��j��1���L.(���89ϲ��CW�g����y�����G-L TX���y�ۭ��4)�uƋc�e�
��T���a]��M������4^ing������#��y���t�Mo�h1����]���Y;����+���O6.�A�'�:}�#j�h\{�Lt�O!i��W�W��xD<7��ܩ� ��ew�ta�������He	�<h�E��2��kHl����+<$x�\u�����vt�">,(|�y�3̚�:	��6�� � '�҄�%�^��GWe�7��e��C{��Z(�(�a��PA���5xv��� гι���-��Щh�u_����-����i���Ȳ�(�|�W��X�EM��cq����䈏Fa�1uT�+���� ��Q�J�N����[<L�8��%%���V�[������p]=!�ܿ�Eˤ���)o�ad�K^�a5;jre6���u�('o�� ��Z�*�[�E�2k�&Ǯ�{�ήCu��[��ˀ���U�����O�0�"K�D�\��cx�(��t��I�{�RE��dK���L�Z^�8��[�&0PW