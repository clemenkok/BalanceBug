��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�!��
��%Y l�׾�m�F��������2�p0�:��%��uV�%i�~<���~��ϫ?Ys��E���A%�����6vzbf��f�e�tK>3�]�hȭc�60XF�ǈ )��i���=2��4�R�����y'��&����?���	�g%����R;��Ԋ�r�=�.Df*ȿ���{��B��7��J��P2t9���yD=��5��v�\���9*����{4��%f���O{��P��l��o��)��ͣ�<�=�uj];�E[���&UIe�9|w��B�� d�vD��1�����C�}y��RLM/��c�8�$�[�2F��^� ��|~������ �jm-�j��EA;���"w�q�hX���}�ꈬ��ܞ(Ϙ�ipF�S0���3.f��T��֐N�3nS<�Zh	З:2W��=�0�̥��JH���5����Uǫ_�S�)�2O!�vW�<{�+"d9�:?�T͵6�y#�����)�\�^S0q?6�u����ӕ~
�b���c
<�x���7 ��h�	""���T8E������Gv�L3�%�a0z_�T�XK��Z&~�b0�.�F/��|�6"�Ȋͷi}�;A����b�uژ��M��orE���r�^��1�{a�`7$�\W7��AttЄ(m���7�4W7�@�qV�����b�$�-Kt�u��A�5�q䍅��N��0�����M.ˢ�O3�&uqv�^��46Tn�F��>(��ʲ��D��vY/�91 [��e�G���,�ꉋ�Ϊ*q A��b:����<pթ3�F!'���ΐ/5C�o�&�m��;zL8�4��A����}�_t^kd	�H=2X`^�J��"��6���|i/���k�Ռd��$��>�o��Ў�3���NQ�3�x�)��<������=7E�mۂ���[�$
��H����(�×r�1?��e��O��@-,��@��hO�힄5��߮�6j�Z-d9 yuVVb�Q��9}"H!��4Z(�h��;mnB�A��E8�l���#���\�: ���n� �)��Ӡ$5�����X�&�Z����qi��N����{�%KS��/e��=6��в�X\v�Q͚1����e�Šj�5`�)����:^z��N��ǵ�;��ڴ9e:��P����c�d��ܫ �އ���%Ǭ�<M��?+�ڂ��"�ո�z�rW�\����fCWep�h��4�0���Z~O����;���X��z
<�O��޾[�/$p�{�RY��Į���yq�5��,���^=�J�~�owk��[����-��m{28,��Y\�{>��1�`��|��u���������_���'�Ҙ��O�#'�&�o펳Uė�:�8=G3��_GZ��-я���#��ZS&1��2�_�o(S0�����o6��z�8�4~Ѱ��
�YT)c�\�oϢ�''��)�������#�c�&QS�U��v�ҵ2���&J�+�u$�*��	Q�� S�Xf�)�]n�\�c����\eN�p��˦7^���N�.��Фv8Ɔa�j���Vh�)O��e��m�(�[�[)lfA*�m�u倳.0���Y�=�5��0�5eNA<����!��>�vxEf�-A��{}�k��_�M��%b���;RэNM���![�o)mϖ�B��L Jz;P0�@G�*Է�p��ʺy��2�.zZ�G{4~��?)�:�#�|�N7���!�0C��#F�*��!�f�y3�6vك�ȍ�]��&�w�O!t�k�:���x�[�l���(��]���n����=��E�\iW%Ǖ7����x��p)�4W}q1Z�C�~<y�L}8в/9s���O�ɢ�?����eUI4��@�<�� �� ���a8��c�T�t�}��c3����ʙ'ª@3�S7�:(!��\ODǚ2��Z@`C�����^:M�ڷ�� ���4B�v�4;(����+);����u~��N�3R��U�Ss���e�6Yq2�D��AH���b�+����E�[�R-�I�C�ۭ%���5d��AN8�u��)�i.8��ǖ�T}
��OE�@l	,L�GqQ,
a}��1�C�y�ͼ2�t+��D��K�q����X�_Ѓ�ݚ4���ҵ�cj�+�o+e�Y�Lת���\/��JÇ�7_m���L��Fǧ��>���hꁠ����T�.M���T�4���a�lA�Z�&���7F�8�d
��Y�R�V�:i�#�>�$`�i���i�Q���'��ҟ�$,~�t}R����'?���ğ����!����$�+nd��.��� SPS2��M��]�ר�����zƫ�����[5U`��kаC��~v�d�<��땚}n������r'à��b����lH9�t��D��*�ǚK�g���r]�`��A.�|�"Gr'߆_[�P��;9��b9�J']�eč�W��%u��
����i�B&u������
��g���;C���p��Z�ĺ����S�w�?ŎF��T�L�.)3�#��P��ۥE�m�<�I} �8(�C��-���:a����0��*V~@\�$
`.�i9*�6�{�x��Z5�t%<�K�۴D�b�����/15�e���\�W����L1���a���H?Wn��_̟4�@����(�}Ր	���/uB��_�zj�����3y��%T��N����F�9x��R\<Z�k�䥆#ɮ��w��2��'����C�ǫ	��"��54ӷ�t9UC��*��Cb�p}E:��X�؜�e�cU�-:86%��R�����H@Uv��Z�.'������s��*��C�`�bֱ1�F��ͧ�Q�oo,�疻{���	���-���ް�ME�J��B���&�!1�[M��3�����:ۨ�c�Ӯ�.�f/�w3���׊�/�A:�1y��gWl)�IU��B����PN7lB'k^7�ʿ`��I}�g�U��jm�|���g���k�'}���k�".RUh���B�i�w�߉d��$��t�)7v��&��I˶ޛ�;Ho
�����L�|�4�axG��C����S�|#�'�DĠx9�˃���EɌ�<4�ί��xMrȇa������Ji�]S��~�dBQ37�7���/q<�)UY���є�d�����+�ʼ���͉Wx�e��A�w\�Ð� �2J-�J�f��dW��P���j��������+$�\gx;�L��y=�C �B�*�P���EӅ_\���S��9U����
��&��x�#���u�6և�$ɿcTlt�������'�ƛ�]������X9�W��g��x�,q@(7�����&���[=.,��p���!��.K�/C�� ҄]@_0Mh;P�j̫��P�7��O�E�p��nVb�UJ��O&�_ �H��شUM�b;=�l�Dx�e��(����mZ`N�U�cGYE��xf�� ;����!����abϖ�RI��d�0ݦ{%r����c�� ��q8������p�.疄�a��.}�����~�=�p)L��Ђ63�}��Y�	�
Sz{3�4�3 �Sk���B���R|ډu���p�n:'k/�F�.��� ;��n}����aת6��oA�`�T���[0n#5�~Z�kV��7�e��@�|�F�3<���ko�n�~&h�3t("Mt]qT�1�:�O}�W�^�z�����&�a��j�9-�
�\���	;3��z�;��G܎���}�X����dv���c���W�\�����H�����
r��;^�-�:4��<�X�j A\��12����c��:�P������"�����ʍ����y�,�6loS�Ml� �A�_T>��F���V�(��WP�6�θ��5������nYM��"U!��XN�Z�����S�q/r�)8�i��s#�	��p��wm������t�]��$@�8LUX�9#]�$��p��ⅱ2��܍%������K�C��	�c������,)R�z�FJ_+Ӣ��o��q{f�����t�>}[~7?,,ޑA~�A�����4 ����w��>F�����쒱ϕb��l�\Bˁx-Ĵ3Y>�����MZ��딟z�qmY������m��V���d�d�t�{Lk8��ou�7s��Q+�6��p�@;��O���"u �_	�z�goC��߆ΒeS��}wj!�p��?j�q%�t��VJ��[�k�p\�f�j ��Vnu����:��y���Z63�M;][gE�b�8�f���v2�2�K�)9�C�$�X�<	��
vZOZ��O�����g�n��6F$��5�	�	��|a�����0;MD��u�Ǽ����}-�0��,�;d���Pa4�"���Q��ka?����'~~�X8�)#�vq��X�h���9:��*C]��
�������9���>ԯ�Gj�@�fT���?�Nߵ`vf���5����H�o��g��XK��ɗ�oLx�B����"���<b�Si�����ѐ̝��@�Wq	W�xǥ	�hv�ߎܡz��+8��_�@,L��G�xe�Y��3az�?�H]�U} ��|m�a[$E4�U!��N�������8���+.qՐx Q{��E9��MO]xz�W2bD����#����8B��[�,��2�r��@A�kxi�0X%�f��d��#�D ��ؙ-`�8i%�a��<�E���gZ6cz��6�,q Ve��@�y�Fe�w��=���^�r?�� Ո���2�J/1rĄ7'�`b9L6����}'P�Y��c��4��t����a��G����;��?)`,����@ޱ�X�m%�0e�gs$��>����t��[*���fh3���#�-[��#e��n�7!��%�KM/Ff��emV3���T�Y��G���)o�xS�G�]MB8(b�j�?"!��4�}�.��H�X,��4�0*l�+P������