��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�!��
��%Y l�׾����|R�b�@�n�?���i��%)��3��M` /A<DVg��?):�<�>
�Ҩ��>\'.��[�].OM����{���yzR��eלҥ��?��8I�j�_�Yw��
�U/����*^��	^��ן����������'₝�����g���G��jＲu����e'��^H���nC�1�-��5�
�k�'�r�g�fw���T��S;!��a�X|"��D �*�h��/b���k�?��qٝP.����(}�D�u��i�Om�|��E��,��������}�2P^�Nï�k�D�<b�(� )�9���^YQ�ߦળL��&<_���@�R����E�n��_�j,|�M_�Ɏ�b��Qn����5�	ER4ޟ��0��qtX;�R�8��2�y.��=��_54�dc���׊�^Z����lӧ��I�m��R�*�?I���0,W�Ue���FH)�Yc�^xk5��<�W��d&;��A���P�PZh�.y[ � ?��m@�x�`0c���\�f�g����߾�A��lĽ�X2�ʑ<�gƼƆ���>���|�Ӿ�`k� �b�܆����	DggR(��#��-\<��mr��"S���b�v���쉼�;Q�US#��d���k����rG�q�Ӷ5�u�'��jȮD|ڥ����iX�xE0��Z5I��펼�_��H�Nt	-����Õ�/��b ��e��0��p
62�T�[��>��o&�
\��"�cG�\�(6b��N��b�Rp�y�h���8U���1�L�D����[~��l���SM:�Gd/�{	�=G�=��բU�͟�<#`�w���8���?���j�����9�Wmh�Dr���dg�{'�~�X,&�Q���>��ɽu�ȷ,D���3h��(�*�?^�����r��UE��wߊ��Ԝ�1.S�|mRt�\�_�9�に�����Y"�o-��m=ۢ�	��й�<x��p����<��k�t��a�'�M7S ����J1��V��%n��O�+&}��_���� 9���0�
[~�n���i�i|l��Pd���M�_�p-Ï�K�B���%(\�eT�2VE?��;~Fb�|	�ۻ�"�҅�{E[��m��7���BD����7׽�z��MX72����v���:��Y6�f��g��'���8[�Z�U}��d�ll�3\�v)7����3��m����F�Y=��)(��(���NOzL�.PR|� e��Ʋ��޷hE�kŰs1�L�0����zb�AW�?�����=c�[/�G��F+
�~v!|I��$�J�?����P(p�_��1��*�M��,��۬����ܫR��n��[S�*B � ^y�#v �9>%͖b��a4w��`ض�I�}�`�~�J�t�J�8Pf�\{ܜ��h&�o�Ui�fw[P�\�r�$�
�Q��R�񥛱W#��b�����S�-R��>8�٭V��^����C��K�7-�]u�Kl�Fx��EW�Y�U����J��=���X�zB��=��������(hx�($u8���xx�TK|�H?�Rms��o�>��@�<���I������F���l���_P�S��F����+��o��4j�V��sΉ��.-�\��I�5��q����s����'u�W]����Ĥb�e�H��/Ę~�%�K��uvr�����u�n>o�Ӊn����:�w�P-�x?���Y#�8��K�CJ�Y��ha�Sm��B?|���'z]��w�^����T�HV��t��������~���.���b��+�4be�{=y���q��R"�P}��f������Hq����f˞_K0��3ޒIW�b�=��QKb��O�R��pָK�U���pQ͝�w�ǹ��!j.�v%��W(���P[���+C0��_3��-�8�NCYD�]��vv ���G�p����ާ�p�8X	�hhz=9!Q����͘� 	���� �d���dq��S�@{�
e}9�ƴ:)����4����M�2�g�z�ZL�������eGH�����@ƳG��\6��������U؋�"Nd]���Eɣ�(�� ��4b�ʌ�9K�ahC`��h�]���v�(�b(��J�T<��ϩ�=�����l�,ŔA�L'zv4���ɤ�OA���-��ZL\��^�K��`d5R��X�E-��0�\�Ia�!�����\��I{�b����V���N/X�%X,����5�c�mf�n_Eˉhw�:0�;�@��4wxR�z����?b�
�a�U��	ӑ\��p��@}���l�
_�F�~8���d�;�u}᜴��7�l�xgh#ywk�W�&:��ݾDQQK/��)i%	���@�B>I�5�]f����*�e.<���ZSWÏ��|�4�F�8���C�7&%�x�����#�:�n
7;���Ui>�R%�=�kR�,��\�lG)��a��10��؞]WnA�fl�ξpۖ���@��Y�LH;~����#�i+h�>�APJ����^Ƶ1�����ȍnJ��h���?G��2��?sQ_W5�D��Ժ���9��_�Zτ7J\�Mu�knB�^��e�a��	�|Ք���N�6Q�j��F<�U����f#eӱϕ���i��$�eWl[_�3Mf�5G��ё��� � ���4(��燌����p�6��2��\ O��iR$/�]S���������C}��%e5���d�����<���[̉�̶�A�������s��c���BL��[�&��5ߜ�����x��@�L|���L	�ä�Ɯ�wOqj�D	��7-]����T� ?�㐉��y�tBF���/��>N�@��n��	�Z���5�	QFrʺ�zv����8�ሞ�+�����	\���L&3�L7�z��ي:����@�3�YrS�� ����ĺ���v��:��
֏�S#U?F������,�+�ɕ���߷(�?��s�ԯ��PE��:�b�}&{�A%
Y� ��}'����w4�o��Cj��+Y~qu�+���^�"8Z\B�+"7��;�S�;Mec%pg�@_�|' �.�gŒd'3����_�E�]�B�.м-ΰ8�E���M�VT
���� ��7��I�҄�Nbg�#�]�IbB�����2'��'��L�GH3���nZw�?���0�v^�6�I�OM�Q���C1�ę9��.s�3ʝ�{��L�=�{��v��ז/+�eR4%��d2���b��<� ���q�'��0�q��5�'&[D}Rj�z9�r ��؎%�[��aU���K��=�A�.Vy���H�(���iF���-2/��n`�W���L�>L���^�A��/�\�)@��%�Y�C�q��!��|���^�DwD��aU��c3K1&���:�`��տ�3�M�0�;Ʒ�5������Μ$ANz$e`?=X�xF�+
g��2f��ٰ��	?~f俈?�N9��Iu)N�N j�%#'-�V�"9�)_�d�m�b��ă�@����2)�����i�J��峎��ZNw�~�)��C��=Y���*�=L�܉9��\�^8����T�.DQ䋆rProE;.�S_�k��`���rKc=;�ɯ(� pI�x9��ٷ��,k~[��YK;S03 1���JRv�x8�j��U�pc�\�Z���iF�4G��v�Li«����z�j�us@s�4�����1K�X#�GG�O~"mK��U�i�Sf��5YɡD6T���n��lN3��j�Bi�����Y/]�L���M�Fхk<}eb��ϞE�H �f�e{�H�-��(�M�y���+�i���3Дz���;L0�.�|���ߑ�+5���q��h&��ĎH�h��gEc�p����7*`�ԗV#�cD����~���$k�yP~��L��h;�G�{I����^�&>�q��p�ƞW�������@�c�q�Ǿ-QϳNb_V�oM����\�(E��퉷b|?z�@d)v����������r�~8����GL�3	l��E"nؼ������=1�ט<jQ!���	sp&=��^`[;�� ��F�;�-4�I�&��j�����+�/(d�c0�2SPs��q�Z�_��IˍV��ghh��@��gI���"r�s����$���Uj��ў�h���8-#L/�w�w�%��Y�[k���$�����ԉv�G?֙�g��r��=���g��#k��`/etFzP&i���Yo���al���^�̒���	W�?>�/�����X��爅��ʃ2a���z���E0l��266��N�ӄ�Q���-����-�J�a5&H�[O��f:��@EE���y8��I#:���������"I��L��1۝m��xF�N3��D�Q#W �F	��0��D�n�v����
Z`���B�
��3Y��� v���i��PF����5�o�����}��Q�Oc�֥6v	/L�%Zhn���T��h�
�]�y7d���'����P=�Z¥5���̚�ٿ�-��pWG�4�nu4����7��Q��������K&���[:��+��'d�sO�_�Z!��(��΢m����j�p �8�z�
����0|D�����՘h�쯺�}�F.s#��W��,���7�
ۗ�pR��O�r)�xADV8��u6*�����d�;=��ݽ��ƈ?�봽,�����$T��.cK>�n)'�cIޠޏ���_El��"@L��I�|�ȩ�(��{��S����#�������޾F��ɳR:E�r�u�V���ֿ 4������bٗ�pa��;P��a�Ǖ�b�4l�8�D0���W��,������%�c�12($�|1��m���!f$��.!�� 6�������8���a�W�U��?L{��w%��=h �����d@G�B�Z�B�X�+�
�W�P�G��7)�D�8`���\��8�����Fo!�=��a���I<
x��j;���(�j��kI�?��e��Q�C#���W�����<H�өHF'� �C.�҃���8F��5�C�C#���������9G �����5E}�ԟT�WI�U���؂��v������I���ɟ�������XW�
G�&�2͗�TKHef}h>:��w�?Y!��.D.oy��v�._*:"/F�ٜ=�BGn���E�Oj��y��|s�y��P ?_f�"�I�n�ɟ�2g7�_�6�Ӻԝ�"��h�5�Ԣ��^���WL)���բ�q=�t�;է�-@�4
��]��̈��\2��)! H�Fs�2	�Q���ll_��i�T�?��Ǿ�s��]� ��R�7e���=K��{�{�#hWQhX�K���nyc��~wCז�E�OZ�H(S���>QaP��ɭ�9�c)�P��q@_�Ǌ����<��nf��`Js���qYord�	u@�:��L[��X�d��z���v�ū#��k�sg�����U���1�ԭ_:�k'Zc2el7�{.~;��� X�ae��\q.�i�a>K���nԐP�U�DX#\ɏ��w �F5��܌���k]`��wc���>�118#��Z��$��r⪭�W6�Dl�wb[O	��N��C禯�>�*q���7u�ӿ+�|l���_��2�uI$k>��hz.^`(2�U>u�� �|�8s8������%ȩ�f�҂M#,����A�6`�w�j7�E�Y�R�����&�4}�2v��>�z�ї���$a[,�|��H�1f@l����
�5:��������YJ4�dk�hKҁպ?W�[�Џ9�I"C`�*;��S�819��Ż7?�k5�hw�@$�#���6I����6�+�����!=�|c�I֟Тg�[�عi�)���ݯZ�7ȇ�iYv��=۵�m�5���A����
}k����?�P��=�$y��X�&I���^M�*U�L�LI��X����S,ǆ�^3euq6,�����V!��&丹(��NI�`A���&� �:~�g	�[�>��:)>j�~�Q1:���$�Y/�Jki�L��Dp�SMF=,����N������alw��G�8���G�$Pb �^hP�U��x�e *�B��):&=yz���'����A��2�����ń�j�;��S��	�l���/��X��Aib��A���ꛠ XW#�<��|L�,�:�*���?;�āԔ��S�{�'Y�"/��uJ/Dm� ��3!6���g�K��ޗ\���6i�r}½�C�t����nn�k� Ш�E�k�+���q��j^���?0h(�T��z���6�#�w�Sz��g\m3'�����N@D�C-�!E���ן� �����W ���AU����u��0)�ÑQdfNK
����j�Ѯ����L��a�3�v��$���R���/��x��X��O��y6� �/wf8�_w�������J���v�z_tl�N5������b����E،���K:�>8�4�ȵ``{�)*eO�{ؘ�Ka|$Y�����
-�A�:�1�e���ʆ�\�I�t4\��&k��Fհjm@�
/X=w�rp�1Ͷ�Es^����RL�
v�������e��aM��ew�l�,�}� ����1@Y�c����/q9�kX��pY���������vG�=B�Ǯսr��& �v��%��l�"=�&¿d��8����M�*ϡ���3/�6#|%����oYs�~�Z�-�ތ�&�m��
hW:4����&P\Yt��oE��&IYX���4�^z&�s�N��?��|cP�q��f͎���DU%�V�f�U �bm�y(�R�~����\�m�Y�Dp�����>Ed<�]��^���^
�^(�B*�f��yIc�
S�H��W��K�9���x�7����8��1�@�mB,��/�1�2��<R�������n[2��L(���ZJ�؜qŚn��6݇c3��ޖ���/ ��j��	B�Ԟ �nN�#��"5�� ��: Ud���?�V|�4UG��Y�C�y�B��n^ihް����R4�zxv���0|e���u� D�/���]=���=����5�O�<��E��j�^%<���
˭�̄VMh�l=Jo>�D��|i1�ɩ�Ʈ��Ų�FY��5��J!�����2��#Ս�|�K�i�P�xCNj'�5)���_�`��.m���dj-����n���GU�&�)�ф�,`�l��`4�T'2{`�+�+�	�W�'�U�C��.���k�kXQT��[�Q�����s)h��g#�4T�;����5"�5��`�9P����?%�?��@��*l3N�ȟ?�;��j��8<�?�OKK^��XN,A�h`��@���EӍlp*$�SS�/�����
�t-Tp�c@��ر�T�A0
�nct���!�
ӄ���^!m��)�Q�7�C�4�?�ά�!_;��ޓ��: l�
�i����U>݄[O�ɪ����F�oB���xUV�83���ڹ��w��2"��.(5:����4z6h2�$�c%qg5߫`<Ք������pm?�Ϯ��&�է�[�-����4���D�y����)pU�hP.i&9r?y2/3�y�R�?AGk��89�����,�`���L�X�,�C[�57n�:��I��Ls�^YXއ�-���%�f����k�M���05�n)���=��۝J�� ��Ϋ�@êt�$�0f���d���ػv �#�T}*�Qj�s��8>�!Fp\1�-��`U����"��@
g4��?�l��!~;��3GO���w��ۧ��'�Lq���'<AC@�	�F�/��ߥ�,�>�V@X��*
Y��h��ى@0�~��P�X�)�-�z���!����ܲ�H���$Jz�N��e�M]�bg'�����	����u�X�NS�k��3oeOeu�9�Q�>���h�b=cR���r�Q�Nm~󥮯k�ش�΢��f��7#h��2w֘��*����~��ˈ�����/uĕ )F����$tF`J ��fxG\$x�}QHk��վ�n���y� ��n�R�5ދ�b`?�M�T��ƴ!7�Zc�Ɣb�1�E�0,���1n ;�e���-~���f#�T߼�]iMl,_���M%^5st4��=��ˉR�̂��%��9���)�c$q
C�b����b�?�v*߭��؅6쫎HU�)�(���|F5%�4�s� 2.$��չ|QY���|��������,���J��_s������~��q�`���l�DUق�Xx-E{�1C��QG���5��j<=cd�&�f���2ea�P�vψq�xw�;���x��N��U^r@8��U��S�s|Xh��RAI:I�uA��wo�������/v�yߑ����~0g,8�	�Ʌs�3��j]#����s��g������4�^�6*^���8�v�ֽb���;���&�g�nO78L����gdH���5��̉ ���JmxڭRi�p2R�9K�J{y
)� �Vd�hj�'���b�^0[�jV�(���=)���*�̪F�V���z-�ȭW3����-��K��G�/�L���Y@߭}�(��u���s�!H42(�>�
	���	�U�Q�����G�bKKX!��tJBx��X�vh��=5�h��7�e&U�%Ah�Y�.��&�����s�)w�Jpv�T��IN@�[���y�;25g���YR2����ݘ��4j��HP%Uo��@��d>L�O�u�����]�aB-�ܝV��uG�<�Iz�)nB�M���vFʺ�����tG���R,#:;�#�_���.kX}�՛J�Z�*&�8�QeȮ�U�0���@�v��#D+���cE��%;�7�o�]\�i[�ͅ���鈸e�3UU|��b�KeXaQ�'����x����"���t�\R_xk��⏆#%D']���ߚ/�����.[�jˏ�-#�+���G <���9[��1q ������j2�Y4?_��~A�ݞ�% �+�����8��l�H`�gJP�� s;�6��c�7m.�c�w[�Maټ��HTjN|@J�ـ��5�m1�Ld~aɢh����{g����������r�g�X���v#D�g�/h]�$�b�_�5�^�G�9$�d���P|.;��E껋��G�`��a����&-�ڕV|�'l8�y^9K,�fƪ�IY��H>�O�g�朤fS�(*NBDr5�D:�[���aw׊��]Ǯ^ak���.`=%J�I���Zw�EU��m_�����U�$%�XUy������X5k��|s�Ow`�(rjN�Q��?x�7���r���Q�I��0�8��ڨS�Ρ� �����W��i��҄w�r&�ց!?ڂ1��J���	d�gD��ZJ֖���m�k?;�Ŏ�ЄǶN&������9��;`h�Gw�^a����3t*j��<�C�(��:#�SK-�U�W����Zf�Ct�L� w�T1'�bfE�k>�� �L]�z���h�x\H�d<~.�
l.��)2�\rh͡K���Hw��;R5�p���Ŵ~�ۈ~�w{~�o�}̣|�y1��;����ÄH��A���b���:�K������`(�U}M�}ɓ�5$m��5�
[5�g~)绫��8��I���G�_#jp�z0��\��t��߇���+�����If���P�6�t�Pa�Uc'`%�Ώ�@�
\�2ڨ�Q;*���}_�־.x�(k5�Wϊ8O����@� �F.bNjx.J�k�,j�*���-������9A/g(�Dl�N�#�?��=��#_J��z�D8P&��ƉΗ�t���t �xUOo?0M�}ߤ<��~�`G�BM��.�G��[�$|2��t�ɗ9�4	�%��	~J���/�b>-O�ݶR���[�ӣT�3@�o��p,�֕���kT�&��	�`��W8� ��}���.=�������F�*���Ҫ�Y��,yd��������|`���,��!d�ӱ��Z2�V.�0�{�<QL��A�.�� �(ؼy�g魊q�|*��A�3s��2���g��4�'6��g�!��K}Dl��~�n�[N�)ܨ��ôԄG��)'cB�{5K��WI��'3�f��
�����{-q�>�,�����4�6e ��\i�60ވ���	r��{Z�ސ3ᒕ��c0�Z�*�'!�i�7�l�r&C�;��/�a��La�Zw��&���|L�`�;��֒�����ֱ�EP/;�����Ms=��YO��m���fWt����B_�2�d@b�[p�1q�f���H`Jh�msũ
������Ǒx��ځ}<���2��I^M�&j{�����Sw�ۤdȀ�Bs�;~ʣï�$B;�{ֹ�!����3�,<R�3~kI�O�͔�8�v���:m�˰�ذ�>N�z�6s�ߣ?�f;���W�i��s	k8�Vx���F2R����넼�aDr�X���n�ݩ� ُ��Rb�,p�1�~��Xא<ٖ��
u۠��d��,P� :� �t�姘?�Ơ@y7�>�'����A߁dKe�범���(�[DwF�%��&��>0��bђ�9c�W�K,B������B7E��إ����S#�\L�k0�D��'����=�߈��zw�m,�+��շm�ۣ6>�[\Om�]*�A!!at��g�n�C"����X��c[Oa7�8tf�� ��#�s)`�C�	q� �P��>� >�58�+����Rض�f��'���k?�q�xTJڞd�?�U��P�e�M4�Iq�ݼ�AIb5t�R�k+��[��O�X^#�2�{�8z	����٭n�s,F3e��/@����z�/m��� ��X���T�%ſP}&�l�#�<�Fe9��3TIϡX�Z�E�Q�����s��V���Iuy�ˋ�8���6��;�v���(�C�����`��JM���u����O��i{H����3ҳ	]e#d [S�2���C��'+�7�l	:R's�o]�A.�\�'<�=�l�S���\�=�����ҩgG����B�����b�Ym�.3�P�� B�#V$1q�����G��R,2�&&x��	J&A ݏe�Zt�%2�=���|| �u��g�Z�x)�J~�ݓ�Wa�OyǅwsG%w�Qλ ���uTp��n)Dr�H�5)�V�2�uM�cx�
�X��P	��1�k��� *��đp����[�b��ʎD[b&w�G���F*2iT<��(�+�^��+0���
m"��q_�d�d�k��F�@	kQy@1��'c�x�m��\K�s�@acL��ĳL*�<T��^��/N��Tp�1�g��)Y�I�L��J%�D�h���AqP�v�GI43��&W� UoZ�k�4��I&��{M�-s�H�a���8ܒ�/Jׯ�A؛�N���F�F�?,�(W��1�Ǡ�r���y�؟0R������
�ӻwu�����҇#?(�?۶~*�NT	g��]w1�%�A3��w�5[���1�[��UEG���M�!�4A�,͔t�R�!�.7�71��%�dš�A����N�I��z˂�`��4x��G�n��ߙ�q2	h,�t9d�O\��I�Nw���LNNii�9�
������$����L�wE��^t���c �X��� AiI��5E�_>�Ӈ�U~��"|�!���.�K�]4_U�i 1�IEЬ\�f9փR��*�����X��z}���g5DGe�{,�.���kqڈst�C�Y�8C����
�O�3R}�`��g9����ٕ)W���o{�����S��jB�NXx����m|�1)���l\l���C��<H�?�
r�7�y��Z󌌎1VB����gfm5��
�!l:�1:"����n� ��(����YCGd���(gQ#�R��������' ~ч﨎���1�������?w#����]Y�6��F�(D��TH��4��U����[���<�u�;�O��$" �U.����;�_���m��H���k\2�0O����^�����{��M���%y�V�����U7G`�o�U7OH5���Djyy=��Bc#�8G��;*Ο��$mB\;���	N�� ��hY�|�D�%���-36��S~�b���Y9P����j�C8���F>>�n<}�1	N��ֶj��Z��6Ų�N�_53� �!���V�©�N��`I�����ڿv�|�����z\�I=dW�T>�ًa�#rRzm��7r��(ӱ�p��=N�R Y]���������DL��4[��QR\N������A.�}Q;P[*M ���k�a��+���\�r�(���wbE���4Av�Q�4q�N4������)$D�}�I7Cc�A����ST=?��=_c�q�W�1���T�d�c�}���!��g!�.Vo�,:��*X�<���
�`�Z=�&�m��K�~��fŶ��{OXZ�Kq�eծ����k����-2��J�)xq��_#�a��R�!9n�. '�X��-5��+���(,��J-���}�T���@�Yz`W%vU86���;�dx�.��.��
�ʱa���"{5�$5W}ׯp�?�.���lAdQ�o;Ãp^k��9�L��B�)�+�c��t"�{T"!%����~!��3��2%n�DC<u\}f��B��vc���8�_�H�n|]�'V�M�@!�>�_�!�Z����b>Q�-(ۼ��M�\6�w�|��,��vYu/)Y��~v�N�c�:)�s�,�p�]��BrSq�k�ݍ�䃉�˳t�0L�u���
6Q	��5�xȠ�U��bc\;v�*��՛ R��kcѻ�{Lh���{ y�C�u�
Ҭ�?�n����!x�uD0��o�`�7v 5�&]P8�ae��',lY{z˕��kf${Bx�/�u����=�ݣN�P��3�h�J֔��_�0���X� \L�)��*P��N���g�c��o�z���+��*�;k�l�"�XK6���M�C�_�P��P�����鞛�UI�/�׸+��+��ͦ�V&O���� �P�4� !�S�"�<�!�hi�0$�5֔�e�r��� u�;�=D�?�4�[�B�Uq�E����p��tss���Ymw �wE��{A��s�\|����pp<}�X��}.3(�}�Ov�>xm:շ�?%��) ?�Pm<�R�&6�غF�\4k�&:H)+%�7U�}�͠;;x,]�pl='��;��f��(���QasuJ/�hXa��/ng�Ųf�=�?�l�b��M(Om3��\\����.��V[��ĆdԎ��@��|�	��w\�š�p��Ga?�����DV (�n�Q��b��;��3��U??w�Z��~���i{��7�� �v�������eS�+��b�g{��'�/k�]�{��dgԿ:F[hX�$�!"�F��vAn��B.�����	iRg|���	;���ڸˑ��+�BE��0N�&�Z�L�ޝ��������FY�i$b	�M���(*t�LO潶/�W�)L�8�V�, #c�oÿ<`V��Vɇ�Pr�$p�F.U_�}��N4��!�o������ ��T�͹�qR�g�������';�,A�/e¢+�����'�B���%0!\j])�_+�gv��nQx��Ss�jeU��ވ�lȰґ��[�q�7H*�q��w|_����''�HqW7q�8�,���i����y*N�������0�(.
�T�˖��W/	U�9���0	�Йȵ�k��3� .�E�����ԔrC ���]F{�@(���"���T��i:�B��d{����C�.�A(q��,M�䚸=4��AJ�,��)h;P�|�YZ�(�ՠ�
1��EE<�tw+��.��M:�UL��jۥAP������$㛆�j�TK�)��:�[�����˽H� �Mh;������&�� �c*���@]�,��{a���:<���3�o#'��,\y���~HM̴6�(Q�ß�𚰳���Ԏ�PP>�;l�>��ѻ��c�Ȥ,T�+1W����E�[�wlw#���,a��Ь�,wӉ��E1��E�$ +:����3sk�d�=�Ig!����8�DX��9GpBZL� ��SF�r�w�`������U�W;4"�$�����n��F=j�kX�@kJQ_�/u ��϶Æ�M~^^_�o���ݺ�b���r�J�X���LK��u��~�N<@n]]���[�e,�Fj��%�D�6����c����{�����f�$�BjC��x��	�aM��y�G���B�Ó?7*���؁��,^�<�ˇq� ��F3�����[�F�y���5���s��u�(�q������R�#�LCe`�Ek-�y��d�}�줘�tM��hj���EvU�Z[��u&e[�g��Y�B�uEև�*
��\�X�va&��q�t��i�p���Yu%�A����LD���u@ ����ɑ2cl��I�߲uz����Pʰ��˦PzƂ:A3PG6�F��K
��nE쳌I���Co�'�m=���{�B��!I���P�a:��,~�1B���{$o�PŽ�r���.�}c[��]���T��p���~��PrD[(�S	�э1R$�s�i�	|4����^��W�����:d0�3����=~Q_�zU��c����V �e�R��l�'�Z����Zr=Q{�i�J[qj�ġ�u^41	�8�aݐ�8���;���e�)#Mt�o>U��a�)����\�'u�i~a*��JN��@�G�����{����,�C�rH0u����0�͐��U�����z]�����D�\����h�'fU��jF��H�Zl����&�Kꞌ#*��L�����2PÃUȲ0a�{jS::SR���ZQ۳U��u'(�c����a���^A2��#t�;Yw��I�M3����~��&以�L��z����fN:���lp���>�X�;����΋tGLł���A�S��!3�萉�+��Yҝ�Xɐ!���懀d-E;���}�>�p��Ζ�l��N(�A��m��pj���Vi�>v? Ǿ;����.��M�}���;����L/hl��86��HD��9I+��Z��P�L�p�d���l@��3��b~�m��2��QxQ&%�<o;o:�{
Oؤ��5��?r+����\G(�B �� 9}w���ODs
�w�4�Ĝ?r�֜�0��Lb��g����<D���,Nu�r7�����\vb,�	_ er"�_b՘�dQ)5�:�0�k�8���\��#�7������!>� Ø��\��nҺt~�b ��!b�L}�!ZJ`ɀ�ԃrW�_ʷ�mb���O
'���jM�A�N�L�J���U�7^�~$��7Xg�)��]�:�q�
�#���a���[Buxn��Y��ņ�T�^�A�1�y�����
�lQS�R&��N"_=*q3�o������|MG2���fQ��Hގ��k����Q 3�
3������k��Z[`z��P�����h%R2_CEB4s%��
�(K�p<�)A�����>�}iI�
l�h����m������I`�ҕ���/��-xc+H=Cxe�d�/o�m �F��T�9�O��.sԧ�Q�5�l!��x��
�s�~�*vGT'9�бZ߆��E�����^�
���3ۓ~�I �d�6!gD�V5\�]�a�n4t�ʥ�1�I#�1	j�^������@�_���53���=|������M�͆�K��e���!�n�Fx������DlV\�`/U0V��`>,3[1>*o\�l
��ϰj���e~�P���x�"���1F�z/�[.v�H�6ի<��-I�b%�Ό��ې�I`̆���8�I�ߟ�^�J�fEv����t#x'�%�d*���l:�����vY�#_/Gb��ѷ����c���h���ԍ�?r��3� a~��)F��=CI#+J���J^��z�T��ݹh:�G?�[���|�[ް��6�"��2�v?��u���v�P?�����╁j�$$�)9h��O��8
�Æ��C�"����VX^i��BU;��#�{|)+�����D�*�̷f6�$ȣU� ��'C��]�S�s]��Y�'W� �,�?{���Q�p�/���N=X�=�]3J��xH��z5>�e3S��繑h�Alo���I�rNF�A�uX'�2;[x�3j +�H�e�g�|�2,��_�a��Ms1�A��9���[{W��捤)R������B���`��s����ٸ-%���n@��Ԛ��c���K&�},(!�;����s�ئ�i��v��E�V<�㩒��`i����7�'��L�k8r�a�n�y���(�7��i�)�?^ѴQY�q��W�󭜆e��5Qg������7h�_d�ӿzuiv�&9����|f�8�� �ɯ��f���)��'PRn/Z�=�s:����P���D�#���N�����2�	���(�l�p9KHp�i.�#҃����UJ�]ס,Yzk�w�,�}WW-�Q����w��8����:Y�[q�mh�T/g8F]+к��,:�)��	�}�F������X�2���eh���a�����I���T'�����Ƥ����
mOL-Z���=+�*�Fѯ��Uj��r6���H�����@ส�!�(O��q���_�'��W���MV}��Ou1��h+8�<��J�'� �C�X*ӷ4����N���E�{-P�nA�?�}	���F�Ǟ�if�T�۴�Ct�(I��V�}	���r9�|���a )o.p��d�1N���b�jc��˺����82D���-�Z-Ȁ�ʘ�kV9�֨�捹}p�s���=�\�u R�v�&xSV�����Ub�Yk{��:��2������`c� ����������Ҫ1�Pj%�I���o%�q/m�~�}T�dC�@a��@	�Ew�.C߯�rZ�Z�d�AQ�Lǜ����Qw@델�>��m�c7mC��,by��+���R긃a�I��s��e�q)�q��nnx�m:1(��G!{���M�Ќ�F�d<�Y�,�=����%eK~;��� ��T7/L"} 	c�ӜT{����~���H�Fo��Xb�}�$g�r
Zg�<��9��e��2�$��c��56�+�M����JG����� ��,��H���E���B�FrLEԭ����e�����Җ�:i�[ņ�����mڻ��ʀ.g^�n��z:3�8��X|b�U�~@ ����C&��*\�ӠR�!H���]7�r=��s���\vgs��\���Zm�n���A9Pip8k.8��.Iw�&��1����%�8����x����ơJ���%�W<��7�!�ɤ�MQ|���Epw��lGB9��I�up��M	LIMү����33�m!K\*-j�]���w�~"�x������8R�NU�Z|�8�"Y�zNQ]�"�W�;f�$j�*��[�+Uơ[� �+��}�ɡX�t��:�D�|��/��F�ߓQ�$RN,e0I_M���9�.����*0���Ii�����DD��x�_���/�;������F��ykJ�Ŏ�ԝ��*]��N��{[V�7����SQ:�H.<��i�H������}ԣ�nT�WNT��h��.�UU���忾�U�4�E)���HɲN�'J �����<;#'���E�F�[��5~{b����N��A��Bs#��j	+qS�ʀO@]�m� }S�����ن.	7	��Ӌ���#j@6b���5�,|S�^'�7)�����"(H��wv��;�׉:vY��<��Uҷ��T/���G	�Di�M��i�E�"��z�)J�y즟��u�m\���q�=K_ǹ��,��ߩ��;�ѵQѱ3��e+.���JH[��ȁ؍n��r���e9���o���d������II��ĳ���[?��#�^��>�^��(�>Z�L�1#��e��Q���(�o���X��v����%�_�Yl��w}��6�".i6T�����(/B���CC
f��X�����ቃ�֧vVp|��q�e,���m|�
�tz�.�wS�<M0h~�T� �5�k��� ߯E��n�[�nE%=߇�pR�}�\��R�gnM;NX_����V�y$��&�򄼫�+3u��F��`��������*��VqZZ����:G�{���P�ɥ�i�א��6��a~�9�}Ȝ;`�f�8Mkk�>T���}�v^�6�>�$-���gF)��@'"1`i����� ��S���_�t�����/��5&���~{0�U�^��'G�S���C :���}jn
O,�1���մO��υ���l��U��*&�7v��QLki"^��)6��z�{�u�����WԬ2ҳ�D��; ��/��.sM���s�N�CRD��f�<g؈�5:3Fr#�N8B!�q|5M�`�ù2d�W�s3�?%�5�Q�J�����fI>�G����zԂ%���6F��rN9�_ˁ�|��@)������"����^<Qga~�k=�Cuפ�@�(Eh*1qj�^���K/	�Fu;?��	��g������Y�&�v�O���>3�UH���uT�����H1�]E�Q;`�jTo�P�Sb�������AU��^s����:�i��	v��c��g���_�q�nX��@[���v]p��QX�'w7�s`7-����M�w8�S��%��^pft��{�Ǧ���6�&�����I��f_��T��cP�Kz-|��ճ,-����`& 8���g��vEk�˿F	^��r,������$>�~#��Z��/|z8(��i�g|�B���34�C�9��Q�̤&�R�`Ze�?�f��uP��p��/L�HN�Q�W�7"Ӵ�\I^���yj�1)�vy�]kV���#�	������(hJΎ���b;�&t�AM����� M��Z6nm[dG�ߴ^!�s�sj��h�2��;�y5�.�l��K�� �ԚL
A㺳֦���WL}����I�Vl�����hw'#�$���f��X|b=�/k.yr:�؛�Ė��P�ďZF�]����Z-��=ۨ7����^,�78Z�t�T�+*�h�]$��]��Y6I(u3J�j��,�1�ш�"ߵ�+ddh��C_�H�)6��8�O5 :��ٰ�v|q-���u�#O��Q FH}< x�6ĵ�ܒ̜�5-��yR�ڢ!/T%�+��ϵF�%b�����{��m���Qݎ���v�Y$�8 �g/�+ ��A�CH���d�,#�(�k%���n�Dl��y���{�&�/�Q�S�"z���;Ct٣U��lRGb\a`�Fu����2$�^���[}�XMl��7�G[���u���EW�An�]���ۯ�j~R]�3��aH�(��4�Qs�$p�<fn��Z�8�o��{�%�����}���M�]�/���g���U������g�P��,�o��n/d����Si;���Q�VbbC?�ռl`d��lB�����p~���{�s>	�eb�)�M<�L�32�@.�� �(����58MT�Pe��%!�>����x�M�K�	BDo��4e�G��}����$K�"^/����0�1�Q�C�����sqmm�u�a�9�n!nN���a�o򏺧���+-kX���
�f����h|��)O��#\�(�m�qSB���,��0 Pɡ��{ħ{�i��F�#�q )� �3)Ll<P�H��8g%������3��r_����A�$E0Kj'H�x�A8�����V�Ns,�k�@ӵ��IK�/��G�bbZ�/����j0?ʱiJƝ���S�8?JF�Z"����|
DRߟ����;;�M����^)��'�V��0�bǾ���q鉲��nbN�h��Ӡ���E�û�k�K?���
�i��o��������gS�/�׋��@��.��S��������3:SzfZ�jG�/[)���H/��wٻ�cbu[�,鰐2m���__�%�C|�����m�ׄ�a��K-������FsKSU�#�������Y�Ǆ���H?��"}͋yw#F�z��eI�3��j%cd�[�e�Q^B�1 ���T���P -M�t�Lѐ���^]3+����פ��B�W���{�����t]�e��>��=(�L�3�G%O,����7qVUx��-,,�5��������,Ѩ1+,��9U;����$���vy�)�~uv��F�b@FcNYĈj�^O�>�\3@�x[Զ�uzIͯ���z Z4�YD$��&L�(;8�a�#��hy*"s�^7�8�"{�=um��U�TM���k�
[�@~�H��U��}���4�{bN�eްQ�=_�eQ´Z>�_�)�C��~�F�;��1��gP5�����T ��"�$�J�����OH����=�}Qs�or0 Ȱj$E��orKɜӋ�^�SZ��^Z��qr�K�u6 Ƕ�Q����*�5��/�����nv'�UnN����^[%<���} L$�ˬ��_C}_J7�,�3��ШOF�^8X� �����ʅG�|:+� ��)�Pc�ȱ�JKYBa��@zC��c�H��뙥������+:�YDE��p^)RO-���$<�6tAwQ$ܟmצ�F���o�ʺF��G��4����o�EA�)���r����+��S�t�R_1�F;3_rZ�3e��FF��>�����j�(zt9󾮣�NSS[�S�.�ڵ���'�a�X�3�}2~[Rd��\����)�ٯ���)?@�z�]�0���[���`�V�t�݀l?+ii�T�c�V��M7���)s��ȟk\HRw/�s���Q�#�иE~q�U���������X/�8�P�~�U`���ճE7$8�U<�"�o�����T[�lHvo��\����	�Vke�o;�tu���C��2�-y6�����u:�K���.R�R����k̃�n�c���GK�!|�d�7��LQ��Nb�vL�]-?b�f�c���vq�W�໪_��yɬ���| �@��[Ч�}=$w�^
>�	�h�Ռ�"�-=��b��'�b���嵼M�e5�.�*F��@>��h����g�n##���	��ٳ�4=5��Ip���� �pȅR�����.����1Q��� X���+S�Ϳ��A��4JJ��aDl�/����Щ�����3�$�?��a�g#n� ����ʔ�L�ɩE�j�cV� �خPB���D2�yƷ�@��<������^���f�$"r������!.w���H֮���r�ǋ�1ΧvmzΑE�0/����Y9>�ؒ2mpu���#��nZ>am�Z`� /=ʚ�Gomܹ�~D�����W$�ԃ�M�ɤ���Κfח@Uit���ioԏ�">+����Wލ�D<�Q�e�O���<�PX�0^�ۍ����zaK���qАGϿJ�l��9�M�X
��$+�&Ӡj{�%V�N(�u��w�}ČC��\����ߍ�k} {�6��.𞩄��L�D��EM��V�)ǩ_{&�?��-Ƞ�~��:����K#S��*��� �!`�q��)��f\�-�ftcw��QWR�4˚��ܖCȴ���Tē-��o���������H�^�e��X�6)�	�̯�u%4]�:u��h%�W��b��iejQ��I�B}T})\@]��<R�M.ڪ����x商��:;�ɳ�"�YOWL2m{y�H���(z�g, ����
����a-0=�7����s�l�|G�m��B��jq�ٲ����v�\(�^x�|���_�h\se����~�£��y�1���q�Lp����T�	{N�Q.���Y�H�ˢ���mB��`�]�O��0]�)�;� ��n−�J�MTM���P�#K�#�W`I�Cg��I�[�ꕏ'���C
�:����b?	��N���2-3Sɰ���
��!	��r�팬���(+34�V��T�7�y��.?�B���W�5z{J]{�b$R =5v���xA�´E�_��'���ql\�rS�UiD�8)
e��.åٞd��w;F���D'{��@���4�?��MV{��Zk@煱?��-��e<;��9E偠t��'�����X���Y��P��m��q�e`���7�):v榣hf����e�^b� ��֢u5V�!<�!��,��A����/�(�;��4 �MT���WX
bq�h��)����i���	�y�*��K���\��	nԦ_&ҷ�f���q��C��q{�u�Y�C�Z���Y��'�.M�iӘ���1oN�!G���#��Q�T��	�� �IY��Iet2:��V�s�(�Qo���u��z"���B)�AqB��`�B����A��R.�+��2�~��r����u�]̇�r�8�;�r1�\cGx��lխMs���c;���^�0a/�����D0l�xj�:�I�F��v>@��h��E�Au���\����3����_(�ןV���g�x6�z2�������1��y)�3S�|NdY���s�x�Bz��L���tKQ;����s;Ba�y�mhI��e�`&��w�cq�1�B�~�ig/�9�-;87֓��݈���f'�X\'�N`Q�����w�:��qꬓPj��6�2�E�xФ����O
�l /6�P6�k�N0 y���m�Ϋv��{D���8 w��=X�o �TK�A>6֛W1�{C�����("dQ��<��]h?��ow\�Kx#o�l���O�n�eOb-.ǚ���x�Jj��*�R����K�EmO�*�LI� X��]�Ϙy���OV-Ѻ=]�F� f���ٲp��Wᾢh��������(��O��v_�;Q(������[��Q¨��~���O��\��k�#���ۼ��o} y��O�&A����Bj�	�	�Q9�a�"@J���~���D�dTÈ'�'�6�Uo��h�;OtZSC��P�?�%C��2��%2^R|�P%�o�&>�[��6u��h^��讉�(c�.��ꆅ/g��e�f�_*
*}���b�mM��@Pi'O�2"yVa�w��z_,�{�Z��ZlԖX�f-n�s�Ȭ�-����g�.<L�9o����"�m�0%e�!'ʙ�{^�Vu�_A�N�G�2�<���1�S���ᖹ�(�&��>����2{����O��,��T��S�i�f�KXǸ��n���(���u�2�#=E���^?H�O��Ȳ���;M)dN��It�3�1�O�_���02.[���WNc��]}�a [���U��\�:ެ�(H��)-����˴�_�:q<Vmu^���uq5�c�I���#���3�n��`а��F�6VI�iE�e��[=�hU����<ͩ����BKB���"n�0&o(��(��֝ʍ�������]`�I�5Q�a]�v��q��H���p����n�*4�e�	@��D�E���^IT�f�&\��O'à�E���&�x�>}��w0��M<��t���-�e���QZN�O�uT�Yd�uv@��>�?0�%PC�� ��x��b����U�Oeq �X/�xM��!�7��^K5`%MZJXU}c���@�!,)"��U{�h��kr{�E�D�j�s2 �T��2���dd��S�I01��?�)�����ifD��J�&�E͒G�J�I�k؜�'U<��������u� ;�88�x�j����������.���_�,�w:���i+7����p���_9NH��Y[y��&GU'�h�~BFrZ�R+Wҧ��X����ة/ 어�����f5ڴ{�S^K��9�Y�6#N�A��u��mÆጦ.;�2���������~P�
�4k���+�Ž����k;?��<zw���8)�07;z�RS��6���:�����%�,�٥��-L@t0����އ�ˎ���t���|���$�]����/.9�G:7��E���6o�̳�7�pZ9���x����	�c��"��R�^_ef�y�o�a��HV�F��BMDa����6Z��Q�
�0Ej�}���r�d�	�.F9��B�f�;�<��������6��SYBo���A1~<.�x@����G�2I�_,�a,���G�����BԬ�����>��i1��:��������=������U���I�Z	����"�S���u�t(��-U�?�ݑB����,����B�����6<�D�����x1��k(��'|��0��� ��u(+���ȍ���z��F����M3�r��d�]y�����RRi���^���.1��=����\X�5z �7��@��/g=�����E~'��)ۡG�2h�`�L��\Fɞ+��C�?$�>=2G2�A�s;�O�H\��g2�L&�`� �� ]��wda��͋u�=A����|����bc ��9�F�_'=58N��L�L���,K8O2�#��Z��2�C{��ƽ��0[��*�*��U��pn�K��c5���pe���ݩ)R���Ãf�e�]](U�x��xք�\�� ��bC,2$�UENSC�̘J@b��5.�N-13k_Y���?����v���VM6�)#�O�;E�HC*bH�0XEK�۹���Z��ڇ^� ����t�ieU�՞�_��-�_d�� &j����)���c����nݯ�<m�3�}~�h������Y�D���4���n��)��ͭ�zL���7���g�Ӹ�:������*6-����>�J��	{�"}'��A-�b�-���d�}?��
YS�Hz\w�� ���%V}���e�C��<.�����1^R�$U��g�p)3�@"����Zi��*'���>��X�
:��_-� �W�%p�/�xS8n�v���Leh�{���p���U��A��pȺi����7�`Bw|M%��$��+����oJI�bu�~(�E�Չ���(�x�Ҟ$�pX�I�w V+�Ҕ���ׅ���7����b���N���.��(q��rs��0U��+�����=���c��^r��H٘���'{��$Kw�8l�����x
���AH/�b{,���PU��nB�4��]�:H�-�;�!�q��Rg�j��,��갲����K����R�|õ#�`\��'�4�����t=>`��-_�b���y��u�\�NsW��x���	�r�xrH8����c\�/�xE�G��WU-��Pӎ����p��X1E	B]hO����*/�^Ĥ�_��]߮;�]��ܝ�k�z@��.��ęRF���Tʬ�w�/R;��D%&'�������~6�8,v`���TB�1��M�'�B���#���\�͈�@h�K�p�!�����f��C37\f�i0�A���8Y<ߟ -��2�DߵG��}�f�'�馿~��,�1$w�T�IUᰆ�.�Km�W��c���I�����ڛc/3t�;ub���^Մ�Z�����K�=�5sW#�ޙt����Vd~h�	vM{��) �9=
��KO&�;-�L�.,D�>�D���sh�'�Q�>�gh+�cQ��W��O�:{�H-�2���;���_��L��Ҋ2���˻�����5p�@�
H���q4��� �x;7
�԰���u��`u�ӟOA�����lޟ|B7��T��
N����	4:�+�/駢g?g�!JkH���=l�"��.[����n�e�4'��5ew$���G�\~&��������9��U?J`hj��qo;~��U�uݍu�-U�ؒ���e�����C\�\��sލ��kHF�x�d=\���gNq��ͪ0�>��,4dԮ�O備���ڲ��i���C�;���YMZB���/��U9׾�,�����wN��+1���/;>�	v<d���#���"/�U���P���Yl����q�_/�A[����i����(c(�vJU#7���t�ۉ���w礝^���yv^�'!Jq,�ǀ]�M�<��)����UL6�K�7i4���m���kR��%����hT�,��nY�`>�?�ۙ���mNl���sn_�3�}�������y#�g���[5S�*#UV��4�������������`���=�̼���cS�w�˲�_HG��(ֲ{��)���̂�gY�4��ak�q��ƴkZ우��:�F��퓪ˈ&x;�lQyc���+�4��㙲*75I�*E�Ν<����(.K�X�d�O� 8���J�
d��4��$w��^�g��j�:�7�����~���(Ԍ*je@Q�j�w�����XN��_Oڙ����y����H@�hq��h��ujAn)Ψ�lU�|�r?za��>(�����\X����rB����	.�U�hT����B����x6˛���{r{��qQ���ɭWэ� ���X�_i~���Jd>G�4m�h��,�\�wW��j�{A�o��w�A�*�)�h�r��Q(�{Ut�鵟ǓηO6 h���QdjXk�~z�G�(��]$�)B�	�J���R����Ê�A}-�j7K_uX�M��L�+)�ƹ�Xty� ڳ!pV?aL�6��X�P� �b#x��!5�g9.�1����8򌳄h�Ƅ��3�@�F�^����+IU�@�~��%����R)�0:p�W��`��!����M̦��$�Y���Zm=[m�J_� ~â9�!x����U��=��+lg	
2S'����.�f3��29T��ۈ#[l_oOh�0l�Ԟ��ky���)0\T%.s�Xt]�Ow�e����?�ˋ�����z�Y��\8
���a5=��)��hr��._j����Mэ�,����S~1B�f���6���dٸ�V*f�ݖ_�6��p�W�ҽ����>��j�:����4k�E� ğk[��/���Ό������A!��[��X�tp��Ҕfꑢ�-[N;�,�@#~�~�O��Cvu���X�:�bwB�vD(]0�� ��6��H��zc+6vnAjD��̭9�>*�f{�w�����H�{�����K|H���I�B�W�0*��E��#`�8��b�
f#�{���M&Kx:5�,~/R��X�w�I�~��h�#�6����p�.�1��_��G����υ\���y{�e��?������fQrv0#��a��SDzS���y���?섅n� ������E�1�vZF�C� 'Qx�"����w�BV�>��=�$� �n'�4��.h�Iy���0���2N�lF��p�u��9��c'l�CӪ�V��9Ғ0!l���pBn��kLZ�_<�;�و����:IFmST3��~��d��>*o\B��߁���=��d��&G�����\4~-��C��ۭ��K�Ml���<Ĉ��7�	MLEUbսk�aM��`�mDP��H��8`�a���f����azɐ��Y0���i)���y�׏s�S_��'�2�&6�q尬e��0���ɩ��`F�3�ۥTY���?��B��HE�}�������`_�������NIx.��QSW���$���2<����@���Οrd5�~�/�@�d-�\j�TF��w߅�e�9٠H
D�}(�L��?y�$1£`�p�h�(��<��@�3�CB�mUAע�;"��o����s��1�^AE+d ��l���~�Q���x|��.��/��oe2�=X����V�3���o�ϛ ����FN��5�z.��������J%�P�&4a�C[at���*KN>���oIIZ�P$�7��mDs�X�`$���!ۂ�JIŗ�����0ܝZ�w3�C����i����	���(k�j�qr�%�"�$����7��/�~M:V	���z��>�? V��g��ʿ���[���ݞ!].\[@�;2�v���Сt�\a����#�:[��;�^�󸬖�2sO��9.fj?6����1��k�7��>����r�h�O[2F�9���R�SOߜ�f�����mr3��������;��C�bP�+�PO�n/~����Dt�Z���g��8j��<u"�`˃��v,P_g=p�~4���.38f?�g��[4���֜���!��$�Ԛ�x����a�hO�,�S�=gz�2�E��.��įv���Vj�,����`|�
k������Y�� #��F�=��려�y�S@�穲أ��qa=g;%��k<D��RR�)#[���ur�N;:�&��`��*�����b�b��mp]��@�p/�G�ǺzC�э�ԲTsL�4�革�.�-fɆp?RAz }�B��Ջ�k��hᘼAN�vb���ͤ�����1|R�g�Zį�KZhR ��W	����͔gR��85��X��?3Qz�"��бU�&ÿ��+�4�@��6��f�p���N�S�@�R�,Y�e�mJۯj�o��ljd�Ж�t4��~�0�{+��#�8��gD?ȇ��F�y�F�@ǏE�bԸ�)����
��?�ӈ����Q��e�����S�7�B¯���ea)�L\�6,f�Z�׶�,���R��U0iY�+����UV�2?v/��g��(;�?��~&�n#��*L��"b�N�P?��3Đc�Z��1�a���NΔb��v�����3ͼ��@��˘�UZS�� ���	;2=cR/Ǌ��
Ft!f!����3�Uv��@#�Q���D��ЙK3�yEh���qGb��uYW��Zm;j�!S��'$����t����1�:�����?���&
����F
�H� �̠g�	X9k���Ϥ�f�3c����P$�Ľ��0쫇��V�"	M|Oʩ�$u$���)� �����p��s�X�2f3�@?I��3�o}P����lu%�1��[�97�{�Xv��$����F���D�.���Z�<�w���LVC��GS�>,��^u1���=���٨Q4F���0�u�8JzA�ɛϤ�� �ʘ�ͧ%02��e����U��!���F�Z�m*[�,ߙԔr����8�~�o�Q�?�ʳܼWb�l6�u}���ti�λ�0������+�U��up�{��I�(�l��,U0���C�ٰk�uQ<.�+hĶ��Cu��M�.m�.��@�V�qP)u?q�	�+e�[D56��ׄ�	u����) [%����U���#
Q�j6,T0Y	P3�����e	Qv���B���AM� ��ݨ���='[��{P�oW
�>���扵n�5EZ�1�����������Έ��q6��Q�$�=Σk/4�m�j�+Q��~@�^�
� r7z���&�,�(լ�l�p��H��W�/��6O/�jŁ�n�G�������r��u�A�կ�m`Fk��fy��ӷ&����}[Е�]hlբ��Q�o`ܦT	�Up}��a�ic��`��t�,qb�@�^�W��(���ET�m�r|��%w�7��䵕�HfS�!d�\6,����h�?�L�:)0Zgf_Fj��4��h'���Rs�踤R�bg��ɼ���:F�&�7��������f
z��c9��daRZB�ds�F�
�tؓ�bnC��w���#�ݬ�f΃��Ӈ�8����x����3�u����	Tg=U�ʥ!�0���2��W��m�z��t!\!���?�d-k���PQ��e�_}�>�#��,G6�ڊ�64��T�ȣ�ݮ��JO��3Hx-G6B����������d;��J�SM���������IS���>#��n�`o���"1yd��ޒ�*���f�w���h&^����=OѮ~���|h���8��d"+��X��8��2�)��ߩB��nvj����ް�� ��p��j�] }E�ڬ/�^> v������Of��78ɔ ��|Q�L�ï�3��@O��@:�~��/�K򠔑կ�,Jj:|���L�JqS��~ݗ�2�@-�E"A*��Hf��6���|�\��e�9�%�6!e R��hQ�4Xf�o=,���_�t��Q���TNTZ��n��C�3��7HxW?3/��Վcl?w巿hH1 ���J �_ͷx��pgHt;���.���x�$v��!��؎��D�Ķs_8wC������MX=�ǆ�����l?,*Qwm^n�0 ڕ�ž���la�`�,�W���<��%};)-0v]�͡l��rJ�ך�܍E��e��=3�Jw8�ܞ����2/`$���ʸ3���$��=��I.�hD���x��D���u��������n�U�WP�l'�4>L�6��81�l��Ӱ�����I�E��<�b���ҿ�ˉ",>XGw	\����#[��#kHsz5�ݪ uE�������
��r�v&ب!S��I�N�b~�'������Ko��P/*���TU�A�3�D����T��`~��sL���N�#.�6H7�M5<n����2` ��ikK>��J5.U��E��b�W�*�qh?�@�d�/Q:�xZ�3�L����ՠrr�!K��e���2������}�8�i��P*��΂B+��3,bQ�*��
+k�~tM�����'}�&V}f1�<�U�����I59��c���r��p�"-��
�2��|A��Q��*oD�D||�?|�<�&t�1M1q����S��6���@�Ȼ����=��^-"r#rp�JC�?��ʀBZ߅�7���rL0�Ц��i���CX��D��H�	��3�۬�5A;4U3��G�s\퀎��Zi'^P��2Wޛ��3[i�Fy�v������H��((�a�+g�1^C!��&�C�E���������������YТ�GYX�����"��F����j�%�主�6���4���[Q��a/2�CåBd���Nʮ�*�m�#�L��&�E�y��2*���y򭟶�!Y�����|�9���(+�v��ɫД}���L����ͦ՟����J���^������չ��gX��l���S�8���]#�5Ǘ���`C{R)�Nw����w=w�ZR����t��O��T1S�rˠ�[�%]TϚ��tJL��,U�ޙ��Ʋ������,c���T�`@��_p��ڮ	���V���o��,Gn�5�LɆr�S����^��r�-�(�ɂ�nbr�tk��U��-N�Cf*n`II����X�������|�ko�С,g1l�֭��\�)(U�yh��AIC���က[xjl���g@�0��s@��d��)���Z����ڞ9�7��S��2�d�?���<��I/��m!y���V��ۀ�5���0,C��t$h�J��u1������ rW*u9�ü�J�,�C]쓺t�S�6
�rZ�{�+���!�	)ɖ~��o��� Q��8R�{��T����u�3@H:�.Ҡ~��>v�9�̳me+�!5� �������b �b!b�p��l��o�o�H�Yˠ��~���k�VH�A��;�n�� ��2\�7>��oBa'p�*br%J����g�^���~��`�Mm����9�]�T���G<~<�7z��"�
�L�:N�\�X��~�2T���Y*�l��#Z��x�;GL��fÍ�H[�_D؟��R��,IK�Zg�Ζ�s��	F'D�P�s�"`s��egj\Aw�I������JF�@;T{@}���V�?B�a5������r��h�m���6���t(ܿ�����%�Ⱦ��U��ڈ�\�NV@�o���Y�>��ٗM����KT"j/94Z�h��7�T��� �%s�b ���f������|f�l=�A�۔��x ��t2�	��:�{.�LܛF�9��^�1������2F��3t��9�m� ]p��%�6��N�1�W�$a�A'\�����&���/�J�
�D����i3������L�H��|�B���MX�c�V��@���QD�(���+|��][�)DX��<A�70��-�Mp�!�!�=;�PlwC
�(��/8���F���x7j�n/Щ��EzJ�P�/��o�=;ܳ;��^��j,����^M8�Ԯ�o��+K㘇=�w�N��$�
ɧ�M��y�[͗_R�a9����Lݲ1ԆJ&��%3_���FM��F��;Ю���x��^�^s<H2���+hZ�2*��^�ֺy��rNf���{��p�O�_�玿^�u�O�st#������z5"���C������
�!~�hH�PqL�mJ�2��%�M��Ѭc�����̷��ZO�iL�d�W�r?�����S~��d/�~,x�m0��(,B+��y3/,�~뛙c���y[Ө�(R&O�U�ͥ�~ҡ������+V�D
��b˶�[U�������f&gF��"��"",[��d��+P�|Ŭ��+����Eװ�g6�	�%�V��� 3�)�=��*���Ť��F����t�	��C1�kw�woDm�����O���!iT���6j$��20������;ؙ#�~�Pv��� �� Hv��+ciI�t�2.�X�y;����i��|1�x��#�k�Iħ�k[���}��x���xT��T�����'�f٢���"��  ��B�F�1��|�[���>�������x��V������NSr!X0�K��7��yԜ�",����;48���37�l�P�e��l��lwYlȨQ�֍�$k�y���m�l9�Jk���Yq�s�2H���U��$���f�bT���ң��y� ���<����,�##�OVqN��R�5�C5q����n]��w�=��Q����T���"õ12����E{kLsK)`�t����5<?',�u������p��&'�Q�{5���P��D����Թ;���UQX�n�bC%0�R�붱4.H�����}���!L0���㌺��%�x��J�,��$�i��x&������NQX.|�:S����җˠ��r5�2��wꅯ��Tl�=�b�T��z�C[�%е�ݬt��AQ��ʮ����x�r������W�vA�9����	������l>]OĪ3�������Tl<p��(h��OX���+���g��)ǫw���*�y
_�Ff���+y#?*x(o{ǥ��O�3�Xq?=�3O�NJE����\�aTy�E�ֶ/\ ��z�<��Ã4V�������؝&� ч�k&B#���o�vo!O�O�,m�������.!f3��L��N�]��k�"S(��G$��GPm��eo�4�Eu`�M�*��M���@H����.�:_��Ȗf���錥?�m[�T�r���no��τ���#��q�z�uf?sY_�d#"�^��{Ųˡz��~+��/�BW�ygl�(���	Ń��!�]n��9��q��W�;�����Y�E ��#}������F�I���8�]��l[7\.�X@���I����j�+q��Ekx��{<�`3�;!7��m@�����@B#{�S�j��7��X�7����y=�v�
k�vuGl�d���F�G�p��]�_�6U���d��{v^� ��2h��ͪ/�r;� �k�i�e�,��Nk�?�=B�y$t��
��܍��J��c�o%��fvH���qhϐ�g�<���i]���2�=�4�'���
(K2Ⱥ@�8��p�ӝ���Zf�-~T��)�eh3�o����-�l@O5��wj9w�1�� ����BZ��n9r(�)����@Bg�݄��?j�U���N�1�V67��æ!��%U좚���I}/�O�z�e�,Bnf��C�CE��/y����Ci�_��Բ.�7+�]��H\hKeᄕml���r4�+a9bc�oca�y��_�X����/�'��j
D^E����!t����@Z�\t�g�pśY&6�_����AdE��S| �)�$���6(�d� ��ጓ[�����Y����N ��`�l�&Sz�ߩ��#rL�7�?�*+��c��[pT�kW��
^�;��(ԺN��Ѻ�{B�������>7��V��[�B\B�م�p ��)��s\���D��%�^΋�6L��6SWT/ZtG٘�%��_�=7�q��$��X�D2�ޮM�T�D����� z�(	(w�ucD�4#NǞj�E��\�1t�<��LTO��l�K@�1(��E(?)��� )�:�֪��ٙdO&j��Vu�`�/���Gߩ?<��������9w��P��2V/�F����&��/Mv�7�'X {W)}H ����w�
�)�F#<����z" ��d�c[��6�����6�L�u��om���'�y����(�V�/�f�([�`3�"a;U��j*�E
���(Q�)p���:ٳ�u�y��m��qT�e��z�AG���*(�ׁ՘�]D�q��N�>�y[�(��xU�=��r����u�e�S �Q@%�eZL���}��Aަ�ǎ(u��� ����N�ϻ)	+�	�a�m�P�t���K�ޥAQ�`ܡ��V�7�:owL��AsZ^�S�������х�dB��,��۔S�ۮ7���F�eѤ@!L_����G���7���"ύե4OL���R��/]'g��t��mr�̅�������fm���L��!��K)��5(B�0:���N������-jBF%��������	��%w8��s��4uDvl��̛�5K�-�<������.F<X�q	jj~{LLO��TN[��!�ܔ�7��6<A`��GK0~�3�E���?GӤ���1�zjao��p���u	��\�+zu�W�Q�k��g�%�D��&d��b�>�U)���p�Aq�?,-9\���P3��1�Ӆ�3�f��-E��.+�Rk��M'���E%�Fp�k����gܞ�����'F��MK-%	�`� �EH���!-ms 6�
�w3����z�ߺ�S����R���pd���
�;H`u�V��RŸ��=K��^7�@zu�jXZ[U:�6M�F=�݁s�>`~9�7 Ǯ�bm}���R��Sd�7�U���˃z��
��ֽd�o��R$���X����4׸�"�)R��g�^Z�D���闣�C=�c�hia�p��%o0����JՊ �p.��	�%��L���Ҕ�����^]�D�IN�e�=a�{�f�t����F[C��'��a�:�h��<��׹��unS�l�CD埌럣�Ω�ZTp���H�C��:��Ñb�L��c�j�� ������b��WJ{��l]eҟ?zU�?��ܳ��(����3�
{0(��P~�T-��y7����,��!w.и�^*�P>�S,��6�_�9=&�֏.l�	�9~�jQb��	�n�9�3=}�)/	2�\�>��3Ӕ�&8�.��e�j�[�.�v�o�IEX�3+Ý�t�T��]�J��S��X�'#w��ٿr�!���"��\n�
b�#E#��2=_���,8<}1�� �P�c��Dj�[�3|
a�as���ca0�U}Q�s����[����	�)A�25 �n��*���@~߷��Đå�eONM�4H5H;�7���g���1���΄T0-T�����߁!��X'�$�x��F�i�ځ �8��	�)WO3}/Tg<݁����	:�'ϝ�"�M�\�֫K�-��~Ɇ�u��U�T���
�@(S�v�g?*_l��b-�	���u�aE��'���`�Z�0���ӏ���L��zm��7���	�꛿u�,V;�1w@�~��_��$CX؊���"y^Ju�%�8��PX����,�u]��v�ʼÜ��W�)[�(˛�Je{{^"`e�}a����,��8˩ۂ7��)5F�x�HXMT��l�������L3�.� �Q�U)2ʛς�sؤ-��:�6��d��h7+4���\!�5�o�R�99��Ƴ��9�����n��,�Z�n4�2�ЀO�<���-%�w^3X��P_L3T!OvV{���%�#�����͟e��S�Q
��f�Lp�8���ysf�~�9�� `�#r얐;v0�b��|K��t����0�Ѝ��1TT�=���zM�Q��&��#}ǐ|ziqt��F9�s�X2����̚�ڬ�s����KxIゑ��Z��#��Ru<02�8b)��n]Ki\g'��q��L�6(��}���E
�V=V�ㄶU��U2Ѱ5�W1����67�f/"���v/�?w���������='X��L�p�K;AɊ����	��;�el�w��碣�C�`2EQ�#����g$<V��ů��ۏ���0�)oE��A���ee�3u�J��@>��pxT�L*6`����7!�/��I��8����#�l�8z��ձ�n�t"(�(�����j��RG:#��.a%݅T2x�7G�1N�G��2z$f�Lb�Ha��X�/����5�(�MLo�ũ//{bv�/EL�p��c��[�k�F4�l2���k2�D�SB�%��Cx�g=K�^�o�n<#,����)%���-t�d�9�\��G*�zT���B����v�4-u7�b���������z7����y'�����	���5L|2��'���
�}�~��1��VZ��4��=��Cw!���ܡ�Dzt�zv5���J�uډ*J�� c�(��f�p��������i-z�g��Aw5
j;/�h{�lJt�5V"�^Ti�f�O	�?������x �,rDX#����@��Y���I�<q=VN�:Y໺���뀥p]L�\�M<��X��������8x������X~`z�S��"0�-q���g`i	ļ~c�i'�S�7�]�㺗�=�T2xp���]f�E�������զ�QD_���I��@<�� �.�W��ŭ�I�D.�@����y������E'{��̾\+��g���"t��$������*���У9�R�z���A��܎=�ͤ�����|~fW�.Zc��G�Ct��n����Y�Z��=�e�V覦$(I�����{`�p@p��ZRލIrf�%�+�C�x�T���/n���gP�%��_����m2��ߘV�R���}��x�zf�x[�������$��Ŀ�<b��n�'=��6��e���mE��A�G��&v�w��S��>�t�k5��"\�Es:�j+L��J�^� �U�=2s(�,$�wv:ME��4�����Ô9��x>�F�� �-Q�7z��� �'�01�"k��P�����N�A�E@��:Ǌ�j��܇-y�o ��מ� ~?"�;�9L3�����T�(����U�����"�ؖ���i��;�OH�|�I��|��'$��;�lqJ�Eb����ت{tV��,l,�C��֏fa�k$*/2�	嫍�����=��f^�Sd�S���Xb��a֒�K����EY�%�2Q7x#|���.`Ub����̗>xq��r��P�_�e��xB��b��dC'�ZQ-�"D��k�]"#��Y��A�y'7�7���w�|�l`�6!�)nX��_��x�u>����#g�%;1�(/!y�c#��7~�I�����������(	�I�X��#���n�Y�]T�xiƱ}ڲ��+(i��U(���$m��^��h'`���)��e���[%-���+/�w[N�!@xW��2�ۥ����S��]G���տ�< �t�Z��VΘ�fV��7Q�<4	3�xP��_d*������:{xG��(�sx�VQA��LE����Qu9+�Ig�Խ0	ae�T�Y�K�ά�=k~fCS����;�
�aL.�?�]$ �����o�������!)�smNɳ�BP�L�1�A%���_�9��,����[��ՐTzp
2d���6%}=Y���x;��C%��w��S��|�v��;a���Ep<o��d����N����XO7p�?
	��-���L�M�1O}�v���"ț������D��H�D��M��	R�ޚ,Y������@8���<��xG.��.d�ҧ����[�����.�rG��u��#:�O�v*�Tu8a1�n�s����'b��
�X�y�,�iA!� ���t>1y��5-)��B=AC�/��.�(t���ng��j���@F2�*:Þ�&�%j��,��"�o�c(�y�����BQ�MXj�}1&ع�.�6��W6�d�3�7zV�.��e��0���9���:9��>2��<)�w�RD
E�F��FfWD+�u�8��~iB1�q��[�Ʀ����3#o}�?�$�W6��4���z{��oi�`(���?B�&tz)`$��3�!�F�@gM��q���4�"LDil,��<~�؀�����ȓ!�>ފYDZ��Ð"��g��+;숹��ͽ��'y�X�&7&Ʒ~V⬊zSN��z	�bi+є�9?��F�����U��
{K谳����Pm���ۧ�'�Iv�\�b`ǓP���iV�A���)6F��:D΃+0#~nZ2�����_�۩�����VK�ב���)V�Pm8Q�d>�0�1#�ĝ��<
��
��s�ãs��癃��_��8�(�ôQ�׉�ҁ��Ğ��q�M�p�@:�`���q�V����CY*f�%Q�����`j#s.O�1�)Op�ր/�=s�,յ)�S��\�>�,���N���(LA�:�_��|���b#`![6��S�a�`쑆����B!��Z��)*H A��F�$�d������ʔ8�#|Vn1VVb��:�a��P[3�Ne���o�{��H��x����D����ʢ�C`���8��[�����2����o}�����xbSZ�L��WT�Z����ʬ/�~�C��$���W�W��6�{�6���w{s�x����`��)�`^Q7AN-�.@ý~�h�eS� bhޏf�y��O%���;Wy}�:��a�����,>������cOj�{!t!�mt�e��l4�|� ��j3�V�-܌�K�y���Wu�/7�@T+,t�J�$Yx�~a��`��m�p�Z\1����������nH��L ���O��p�_J C0��� U��&�9�w�9�����^���o�sW�[�˔��- �o�*�f��P�I��y��������IϨ]��|�;dM��Re��ZPo=^�@�?�/�T@{�����c���)!�^���Q(X����lm�J��;ݳYM�	�����$dp��uײp	�/j��דt��6`�3˻�11�ch�F��������'_���)��C��.h��Ju��Y�y�*��W�T0��Ecנ��О��t<�� ��(�s����`H�H�� =��)�#����|c�O�@=���(�ۨ�U��j��)M����eZ�*��E�ŤŭY��,FSӧ�A��K�o�I�HPɦM0�,�R����妀����C�z�C�3�֤�r�� �|��;/4�=�D�o�N�=�Dm��>7X�TC����;�o9�^2Ѿq-X�$�? m�{�r�·Y���T�@l�E��B�s�z�E�l���&�e���t9�[�
���j�V��8�b�dHu�"��-��h˷z1��gmB✲���]������M������$�������W�W#�ԶU�`��CaZ���Z�y��-q
3k6���������@3�^}CfN���'x��߶<w f�G��2�@��\�=V����H��!l��8W�gxBFw7H��G�ģ<���v/�.��;� 4[���c1��
;@m���.�j�<��pIއ�5:��U8X��dZ��<-�5|ȉ���gP���
4��$Aa�C���Q4(�wg.p�4���Z�c�-%�/�x�F���ϧ���%ٽ[oz�H`7��Tb1�C���M�I�-��(�	]�:�Xa�߀�S�D� o)0���_���-i�X�3��KA�bc�Z|���Ҩ��/�(c��C��<�Rn�m.3����XӍ�2z�����~�D��,�Łb�n��:P��]l!]�Ô	N�\�`���
�'#6�m��X�c����d�銀��tG3~��+�#���k҂i(a`��؝,t�c�
�p�w��&*��V���K�8�-z�����XRN��ywQ��������SP�ߑ�IX�T����0����q_���X�}{D�Yo���g?�F0��$�17<L�[����2b���7�{C�歀�P#�	hs9,;�!@K\uX&o3'��*�GT)�֝}�,X�ڲ���$h�`�Q�3?�F��ka��$S���Ӭ�n8�eq��h8���&��3$ᚒ�Z#�n��l����.�����f�./�o�C����#|���WqG�#/���g�v�+�q�_,�0��o��^h��6�ۂ}(�������ӏ&,�u�F%yt~�-����et�挼Q��ޗY��G��9��+:´iU9� ej;�e���Q�M��#=��v�?������P^,����ȕ:k�(aM!����&5�D���.C ����#Vw���`���7��[�h0eI�k�H��a��Z(J���1�����HzB4���;ĺw��7�9͕׉ά�6�ȶM���i���w�)8�޼��Ϝ�3��C^g��~ʹY�1��n i��;��a4��"eh���}�Ǐз<�㫿��t 7t��xV1���΀����~^�5���e�����~�r�ԗ`��S o g�@����;%�J;����nS�ǔD�~k��UE|�(
i������j{z�&Z�3�J��_yɇѠ$S*���X5�Pj6��F�FZ�
R�GU,6`��^Y�D踉`>��qJח�/~M=��[�
L��K�w���y������=����N$w�d9���f�� ����\��E��2.2kJ�Չ< *�������Um��OlՃ���ɛ���!un��~'�����o��R�����\�R�d�" 1�q6��
�pZ�S�-��=| ͠5�3�i8�3�)Z#2DrI�<�H}�n�K��#���� �F�w9z�.ú� ;?dB^��,p���R�q�
�2�(��b׏�������9���`F�/��I�2eʅyD�g4K|TP����f�S�VV�C� �a�j���&�������hC,~jg������Ȓ�����ZT�5��D��S$jX%�Y_�#���`�Nj��~��#.��N��z^0��| ��r��f!���;�L�Т���F��S��9������)p���g
�ٟ��
cʫ����S����	�`lfF��m�C��EUg��,b�@���6E��&e�1n�Ǯ/n�l�+��:�7�z�������g+w��T�%���Q��z'�- �NN ::��Y�d��ω8���)�ީ�y�����J�Sm�+�8p�2���cP2�T4��D��m�u�Ne��f�h�u�o�Y�Xx♇� Y�>3��V�*�W^ac�j>+��:m�h�\nJF���h�� 5�4�D����a�7�"�8���^����q�b�35n�"�L���w��
E��㈄�j{f��^�k����p�÷@m9�Չ'8e^]�aB������-����1d�;��`r%Ơ)6�{����էu�G.8����Qz0����F���/�3�Vq%	b��hw������9ֵ�į�V�[l�%p8(*c:�[CZ�)xS�����fn�k�@Th�	{c�E�|eD�x�LA�$�BDV�Y���Ӑm�nm�����N��J~��ւ1�?u�D(x49K{��<>��z�q	��U4��? 2����GU�xbA��%!���2k�a���׽p��p	-�վԥȃᡘ��"�/%�C�!�oy�; �԰�#Mw����+��Η؀tE�73�mO~�n���H��˩����9��jy�׃��ij���ϟJ= GֺP���
y���W�B���N��C}e��!ֲǧ��I.�t�|3J{16d�GL��mտ@:�jא q�2�֩��G��6}W|��C�e�4�,J�x��t��j][1�S��?W\���f��BY����0�Op�szR�	�&�C���UD˯�'�ܳ���p�
�n�Շ;��J��L�V�� l�ϚI�m�G��
�� �	i0�q��.mg����|���m�Q-� �����5��"�t��^s]�����~N+'��E����VG$� ��qX	�P�oe��K��p��j��@wJLa}T�yY���D�Pi�ɦڟ]+��{C�
@o��V}��eĺ}=��!���	������}>._�L�D7��w�֧�+� Fϙ�y�Ի�u�T07o=��;'�8k�$��"ţ�j�Ե��4�X�i���AA?N'��%��Լ{�v(	h�QB?��	��/'y�Z��Q\�׵�����o�6ϱ^Պ�:�y��JO0	1�B;�����7��71��OzЊ�k�&�s��"[��son�3�T�˳������dZ�y�`2�#��K����&�t�Z�;Lt�ݻO�\2�F���?q6�D����,1h�Cu�Cg�%´۽�qq��-:1ls w�v���"I�Q֢�`��5�uN(�K^2(I�7H����O6k����)�����-u�f��߭ڀg=,����*r�t��
Y����:��������W�!��UNO���u�Ɏ���O�Z=9\!�;�qcK�,�!��wR�B���!���`��*$�*Ɵ"j���>�����{去�����&i�[�z��W)Jnu���<��ж�JEe*��s��+�o�J8O�jȫ����a��[��6ݿ����eTw���м��wT��ۿsrt�{�P�3ly�s��_�
�?�,����+])�d:�%\��c
 �Z��*"�(�N\���/y��<Q�B����
q0���,O�I�fN>�� �q2���v�=�ၛ�|�yJ�;�,�G��h��@D�m��Gۣ�əw�.U�ȳ���W6�6*1��0`a+
ax�nFz,�LZ��4glJҹ��s���+:��$4ZC9�єB@c��
��( �<5&�|8Y�V�m	�
!�v[���� i�ә1�����b7"d+����G��ߒi	�>���q&�/����뀜P�jQ6*�T���D����m���t�xCV�Y��JqG]IA��� ?'c~D��%��?Unh�ZI/�w��#ur$@�3ȋV4K	-�0
�s�ֲ�Q�H

�5��]�������u>WQ�)�~Ŗe��4:1����1'��i�E�N��a�G���"��gn�F��T|��5��࣢&|;�R�
�߻��F~9FM
9^� *c�0�����^xw���h!�V��ΐ�_�� ,o)aV2O����X[&��,�m)˨�3�U��]��W� �'���O){j�����`�T���5JϨ�vܽ���AK��з���GL
����51�mM�̺�7(��K�L��ZT�E��x�j����0���&n*WIN�g���<҅�6�	��y��^���Kj�n��9��8�v��m%���t����s����95f*�v*���o��i��F����H���H�/��Pf
�l5n�c BD4k�V?������z~^�LH�� D�Q�X���3kx������ZV�r۬�+�*o�����y壋w-鋺˦��Ҏb����}cE�fg/�Ӫ+sa���})pX#4�oc��ԑ�0�p��L�v���`�Q�l1�0q֎n}8)A�n��p��� %N{,�S](��T��:�����ԓ G��=�1�ri��9\��<�e��v�М#�\L�ۯ���Y�:Bh���!�Y�@���=�YZ��(MG#}b*��Z0���G.Nh)�p��p^�+��)�d��o�p�(���iԔ[��� �A�� ��� �B �$�]�7�Zb�r�Ns9�>��B$K゚ˍN���5�:T2���T���GXZ�<b����8rQ��ۑb!թQ��w�˟v��Hh����<�R���ek�|�E���9�6A�kܽ�w�Ԙ6�7f�*�C�F+��E&Vɡ�I �23K��F��Y���)ʩ�*��?㦉��jR�����#�Ε@��4HY�8o��F�h���y���92��l��@��g�1~�be��,'"㥇��qH�u���K��숔�N����r<��`���K�ɹ�ۘ⃕y��ѫ���opbgl�ap�KVϽU�~���pˌO��5����C��8f��}�qŀ�*�x�R������=7������`�3M����'o&��J@�E0e������~���΄����n8f�?Zum�3��q\[�����D������&��ٝ;q���J�(���i?��<���r�gL�2�-���Xx^�`~��4N�2�&�o艷ɼ�3? ���Lܷ��ž��_���kB.�#W�P�ƥ���|?�q%�Z,��
AVHp���m���V"|c&��c�Eq3c�Q��S{�q�ʄ+�䰎��7��{7M7<�9�������&��gGx�wVH����kƗ�c
�_�a�gQdpm�)�F$�!�z^��r#����}�
_�qGR,�k�g/�Clq�?��eG��Gx΀�$)�;�j#�������gO��|i)�hP�� ���᜿*�k&a�z��7T�N��AE&��k�L����Zp��)�Y��8�+�؍���T��;��:��Hp��� �fN�Vŀ�#����R�u�x:Ȩ���""
PgNy#wV`��9`�8���$hb��$p�0��wm� ��9vU$0�1Q�t1��Ɍ�˨W�Oϖ���66q(x5��e0�D'p���Ⱥn]�X�?���PE�,����#�$���@�l9�J��_�mz�)5e���O��*��]Hr���hYJc�\�o�Q�^��n��e���L���Gm6^��|���ߠS%{����Ğ��
�=(/���E�	��Q�0�ֳ�/%J�g�&��`� n�92L�W�7�C!Ig���Ԣ�����N���� �~:,���
RL�JI$����chz)��
��a���L�<��Wt�}cok�B�aq�,?B�A�US��ܡU��#�P�f��k5Z��I��Fz�{o�
��E˶�����9w.L�6�� �s}�rR���s7�ʍ��6k4�m}�;�i�T��GZ'�WZ�0�%7�4�=�d�m���ދߤ��z��&,v�2�8��\9�Һ���,����0�?�H�fS��	��3��~�{A����e�=�-�>�/R�������W�F����� Iۤ�'�x����Ѱ�ST��Qm ̠�bt� v��!c"br�zy�h��`�pH�>_��/;�SQ�ӯ5tE�)/y�q.�
H�8e(:�uNg;��,,+ )�@��;�?�;��ڧY)kj��3��5̄����e��GL8^�׫�����_n��R�/�W��P�(�v�,4-d�����i�W��T��\&�.�oM�b�^�;�E<�l�QCn<�C�F�.����9e�D�8���rz�L� �wF�A��D��	$o��n�y�e��^w�zs�QG���/��ߧ!��D��7�!*d�2� Q����)X�$8j�R�_b敲B[j�U/������x�ɒ�h;�K�Gɵ4�|R���>C�ެ�liMV�=ږ�E�,��o�Jv�\yĕ����BvV�8��3h�ˣ��뭶���1s��e�����<p�l蔳���ֱ=V*H��٢���q�O Az�gB&��
�ˢQK4Vf.	!b�D''�����B�=y�u�H�vS�jo<_�jf�dA���	i�c���g�3Fk^�-,���� D�p5�O;�L��h�A��G���bBuo���/��ߑ]���� �B����R�"��PA�j%��D8³��WU����XV�N2�
�#��T"�X�#/�p?t����Rz�m�E�g�g��e�~�����|�l�	�[&4�l�0����;��pŵ�[/Q�/��*�P8�$]���X��S���į\����G��f���o�v��#�L6��M������Ϻ͖Au�Q���'"s�ӭ,y����G��bꡟ������6([]u��X۔�X=�g~vnq;�L�0ӝ�q�e���$�'��r��	N��^C�n��s�D�Rq.!�`�2�;�\ԇxt� �Mg��cp�4Xb� �Bw˼�",���)���2��#���U�
����[S~�Mw"�R������bȞ*�����	f\P3�ξڼL�-�)��x]�m�G�m̕�t{����.#�i�x2z�sԃ&���`�u,���&o�F���MxX��@���6U�~^��S���D�v��ۺ��LT�� �)�@��0$�Hk���鲪�'��V�BD��=q;�Z3����Pm��÷����K�V,�U+�s#D�� �~�9���C�bZ>)�T��uY��B�j�W��"�� E��p�{Jh2<��Vw���yGBIBG�^�yg�<��a"I����0���^�ud�^��g�ҍ��&=�V��1,
��g��F�����n��$��7�^3�UB����5_�t�wV
��Oh�3���8������D ��6��'�q&���g�1����-v�&�qc�X��H� w��%�<P*���l���0>�sE�s�u����c�� �g�c� V���e���X<�ͳ��
NCA���,T��Z�S)�b��C^�3$m��WǺ�y*S5�'�	��m��`v��u��}Y�3�d;�����q�ߍ�n��Q&Jf' ˎ�����)����� �˭� �֡��������&���Y'�i��(.�� �zu�b^�R��G-�������6��3z�nX$�c^��s�K��%�E�w�'��I�</R�N�������}}#��!l���ӧ�h���uV��AI5j� 6?Vb��n�����;�Y`YDwE|�#�W�� K3g9���+�jE7G����������|F��)�i����CF@K χ t��o�)tFhEX��Y��Іy�;^8��HD�ߔY2�u
�7#!�/���౭{`�4�J�L�fͲƌ���v���ml�w9�%�[�?/�eGNg�'�{��a=Uh�ba)��}�u�Lb_l�@wS��VR��t�J�{y��0��v�5��3�%ȓ
� H>�_4�ߡM�����C��A�ǧZ�bek#U���m:�(�&���7RI�p�p�uuܗ/GP!�5W����9Α���ɴ��_���S�;q�����p@Yee^���f��6B�� y�����BhQ:��>'�&�v�v������qD�G� @�c�7��/��z��N��&M*$d�F2��*<@�-�'Fd��ajxN�\�������B�rX�#y$��>!�.����8��u��b��%~r)�"ZXYȷ
@�Xgkv�z�޼r.}M�
�K�b�:��+���n )`�u��#��14�K΅NSA|廦�/�}��a���d;��y�N�C_�f�J݌��"���������i?p<X�u�}W@s��:Q9 �s��A�DD>܌�ֺ�(Zq�
�bP�A`��~�.��Ņ�%\:��C/Xv��{�"��99���ͧ��cs@7�����6� �KvKx-�(0M>�/uz�NYu��t��7�0A����K`�����v|�ɿcǆ����>(�Xd�m@��I�뫌h ���<m���އ,�V�0�����ؐJԯ��2�RF5&�OãlsL���]�Q��o0�D�[�V�.� �2��n'ޡ�А],�=%gD[2����+�k�~&��n:����[�9�������Ia��6����R�lH���[��SU��:dnm��`'g7��ʹ��A����h5Gɋ7Ϥ�H���үˆ$�Q�&j�Px��'Ʉ>����U�A�,\�>Z��~�n��������r�U�w�'�{-�)-�'���k"Ƶh
_y�ew�pf�vu�}���2:0�l�NSǿ?S� Y��o ��^@᱕@%���5u+��L��/~�[�ι�0���fZ&��Ņ)R�����;NU�2�������=�9�ZU�t_���գ�>���#��уk�7A�,�	�C�j���\~B~C��Hg�@f���=Zɗ��es5%��}vj&�z����0ڍ�v��M�f��"�t��<��g����5l��B�@�(D頷�VsA����Y
4Y��G�EҔ���t��괄ozl
�4��lب�a��s#�XEiNq/򬋓Vov2I3#��@h�Eg�\M����o٧�C��z���j;���8���=�eM�η{��gɾ�Z�%�s6���`�#���4��^fN���i�A�Dk$٤��8����Z
��w=�~�_�eyc��]I�cn˝R�,�R�*suܡ�k:�6��0g�*���V�~k�eV�#��f�]��Y��j�C�� G3��G�e��~�<�;�>+y���a_f�{�3tG�3W�
���(a��!�!H�����f��ѧ�� 4tu�%�V����ǈ&�L1�'���xTȲ:~`��X/��L$h���k�~�A3A��e������g��e=��'בo�[�xdU�R������]5�4hp[�����r̈́�e��!�,L�*V�A4����y����z������C(�ц�����!.�ep��U*G-�&��M�����b|�1�j���c��s�b�ظ��mϽb=]�≅���5IC���.��fJ~5+s����s�q�ZhunB�	���FI�"X��;ő9лRT���e��F��6�۟��n��ke�>7Sᬈ?7n���8��&�
(O}xׅb[��vLX����f�ql,�Ioo��!�Gz�0�VX����Қ�h�u�x�Ց`�r[0g<iG0/f�t��G�^C4\�6���}$���"]����=>�n`��K�Sf8�Ap�MK�z1i{�gj ��ک[ �kU@	U�����u�n�z`��j�e���נ���8�!b�9���i��9��A�e��!��1�4�o]�Xo
4����8����H��!j���/��KZ��21�BH-�t��O��.���<)�Mz� |_�r��U��RM�������<���]�VJ#�ơU��8G)��Qc���8U�ڟB1�T�s�����1pyH�rz[���Sk��������ǟ�	�f{k�)\x�R�,0Swg��"E��|:X� o"9�M�2����@y���y���2l�z��NQ2��*�Q�,�J���Ӵ^��(F�yE#8�C(�i�w��
�s�h�W��TЕxC,}��S��e�v���4�@đ�u���f�|�ά�oG��j�I�~D@�hs~��5K���U�A��Ӛ<J;�
��g��p����W�c�Ruaq�^�_�9>+�RV�2h�g�������T��?@i��MzvZ-����(��e�K��������7 *����V��M�D�cy����y)�>���4<7I��$#����K]�(î���2��^���oBL���Ǟ%"<�Hu@��ͪ��ZG���P�z>�5��>9K�F S*<�)��v��\Jwc6�y��v+�4�'����Ϯ>望�8�5�qw�lJ��NTɗֻ�&�ӄ4F��4!l3J��J�� �)�3�ܜ|�_�o(�	\�� ��oE�5�Ď?��)�`��'�e�mx4�����Y&�i.�WF}���"At�Ă��c���E�t2&\C
��.u�:���iȹ��t�@�!�vb�'Ѓ�<��ڝd7�ϑ�WDG�3x�௵�o"����`�*.v�;����H�'�x�ړ8��+�P݂���Z�z��\4���lo��><��#֌�**���A��U�`jb�q��Wt
4z(
HV	����2�;��ӳ��F���pN�,=�Ad|�B���ygI~gAd�f�.MHq3��S_U�����3Ph�n|i��	t���f���"���]�F��}/�D�5=�R؝�� �-�'\��N>�l
xz,SǨ+�[ *G�*���AT��n-ރ��ٓǂN��78A$%�&R�w�G&^H�K!�3�n��
"���� ��f6V��xC@���ؐ ����.�u�^H�q�B�9v"v�)l�{v\�W#�{��t�ɐ�<~��pTz�;���u��uI0��E��.�.�k���Zh��M�[�}�ӣ�<O[!�|���Y(8a��0�K�"�,!�)\���"�U�ڻZE�P�}������u�m�����������|.%������a�K�2�oKs�.K�ߍ��l���Qq��>j5K��R|�c��<�����m$އ����l]нݠ���2TO!�"��@�Cz�
CB�|u�#g�a�I� <4d�qd��u�7%�G|�E�\�r�CC����T5?Ziu�.3�:�/Fg%Hv�m,.��'�I�J"��/����5����Π�ux!�>��.��/���R��W�o��=���/|��}%fQ5t'�
{n�[�-9a谗�u�ˎ`�Vo�Y�zdnK�B�Pr;��v_�ԙn�̏/h�O��qر�QX�ʂk}�݉�퍉�۪�yU��w�PE���^�#���U�I�ڼOJ��f�6|�p��D�$$�Ţ#�F��z�ᬵz�l6��35y_�槼��+G��%�,�B{�q�t_0{������CElᑊ����p=��W�p(oQ�R�W����<�Rߺk;<�
1ԻWv%,
���ë��
���轇��֡DV�[�g]Z>�Ǒʍ+R��Q�m\d0���t��ju�1/��	�|0+�Q�*v���#e�~���.~C����?Vk�>D�|���_Q�+u;=��7'tҽc��Ǣ@�K��6	�5)Y ��Kt6-�<�J?�j�ۭ���&��(��R����N���c5�/)����h<Yl��K�?���-C�}^Ads��z��a;�r�'�B�j�L%c���L��.��Ђ�p;�Z}������PJV���\_���xF�սܒ�%��iSr˳���F�ԝת�TO&;�R�]|�'�;���Z�G�,���JY-�D��	��B&|[�U_�?�ߨ�p1I�Ӝ����G�C��`�ĝ��$�L�=C�{<��^|u؟�����#J�o����gPu@�V�����oLQ?����G���JR��#	��*q{s�)챛��_��۬£q�+8w��h|iӼ.�0����}���˃b�ּD��xr�̦����U�X��a����,�i�W(b���_��`��R&M�u�̇˿������6�iѭ*�\,�:U@��fi,,��|��_tZ����2�L���5�,�+!��T9�MZ�"`�.-�r0���.�ﵽ<��/���T���}�yE��[����S��^���Nut>O�ӹ`�<e��<��[��_��g��j�=�G�Ŷ��w�X�#���ڒ^�ӀGz��M��=��ߛ����]�Z��Epǟ�eʢ%쎵�H��n�)rǓ�׆��&(��e$i�:r��*������cy�,�]���-�D�OSh�y.V?08�͞`�;�p��&�\�n�zx2��A�T�'�1��ڸ�W��[1{��D%����*��������U$݌�:���))z;��v�
��g�Me��#2���ҊΨ�݃.(J&��)h�k��~�wj
o�FT����\<�m�ё��\f4���r�b �>D�B�6�S��W�d1�=Tv(�k��t����)�fU�F�Fd�@_�y���E��o��i?$�C�?��0�k(��H�+�Z���C����`��l�+�V��r��=�B�26C����[�sGg=�x�`��-ބ��zv��'E��oLV�̗c��Gs�}��4���9$�'E�j����a;��~:2-�� n����<�XE��2@���xK\�-�3*�)e���uS�EW���2���,ۓ7�S���Nw�;�M��3���s���pfЙ�S��n�N�)fF\�/ا�����V�p���"v���56������߫9^�kˤ�`���-fN�W�%H4��x˷r(s[�b��L�T߅ǯ�����)�q���_)���5�-$���	��.�@���:�㸲����K��t���C�J���i�F�i��ڛŴ�Q�����"�zLS�6���¯�œ9P�������[s;�!��^?�\|����@�[0G�E��j��~���[	�S��!���m����(�숯�BK�J��5"�Y�A�‿��],�6w�W��t����EBi���>�ܯ5Z1Yy裭�i�,�5��.�\ķ�ht�O�R�0i�d �%P4�XOz<pњ�U��Xl��_z�b�#O�.QP,��J��ȷ=�̖�Ҭ����)��{:�����r*������S^����
c`����s�py��&�UP��ȨV}����A����-��e���m�AI3�*���sn|_�/�S��B��44�˭��3'��:�P�e���@�ҋ'�"�lJ�<�n��B���#��+~�gm5&@,�F���|�Yg%�$&M��1�5�	�� ��ۯx��Ԍ�7Y���I/���I�yG�k�j�2j"Asf�GǑ������:L��z]��ZO�i>Z4F�V�=�*�m�\������;fd��#\Ɲ�up��®��^�b7O�6�Uq�bH�|ym�W�L������9V�nr����,?)P�ʬܘ2�`�Th����1lRNx��?���H����:��yJ�,���:��3�4�'����Q�@-�nA;$��!ޠ3��XsŌ���o��7?�m�y
��ۤt��w'B8"�%`!�v\ R/X�A«:�u.-�t��l��dilG����c��xT	[c�������Pl�v�2�X�/e/�����X��he��1�2k�s*��g��[�k�����`P��s��jl>y��h�� U�1o�*�d� lg(��K�<�a%k{�1���Q��u�ނ.H��F�9��j����=��L�hr�n���G�	���H�Q�����y +^���A_�@�A���A� '�\n�)D�](�WHO���_�!�ٴ�E��\�O��$1Fb���u�����+Y���fs�{�T �ŝ�c�����)�i��|���ٳ�nI�P�IH���/����E*��[>6�u
,�D�H�7��5)Xv���K��	Or.��X�^ʔ����pH"�g:�:_��4K��{��&e�����~��b����;'�j��/Rz]?�e>ju�w��:����GK�s�xU;�Y�<�$V��Y��%��NQS�������^%x�ppJ'�9�z������7_k���HjJ���҂3U�`N�u�8^
�2'��S�X�������\�@Ѥ$)R�_�}Ҍ��L2�����}@�g{����N���A@g�x�%�܉ق��*���.���Nt=��*��f� ]�)����Aas��M��T+�Q��f�������ŀd��g{MF����0���iR�Irt5}e�	�s=/3]+Z�-;���\�I��l��IY'+�_W/�uǨ�]y���m��e[�J�Ǧ����T�/�@�86Rh*p�X��WO�MѸ�>%DA>�7y@�v��:�᝸���gK�x2�Te)��O ��6Ks�Rʶ�7�4H��77׾	�+��\Q/CUM�}#A�'͚�u6b���,�}h�ۯ���ū����9�!
�ٵlRȝ4��-X����L�BƸ!����X)����%�ߠ��W� qfM�Y�%%����v�9��om��Z|G��'�r���#�J�l�F���	Kܓ)���4���g��R��d�>��[:��|;0`Oůg�N��Ӥ�=��&S�����e�]��+�'� �!QUuW`��(��zG�G0D�ǧ_�y������o�|%�Y��d��v=��>�H'�[�J{4e�1���~���'L:7�ǅv�!�N�D^Jh;���#�*X5 ��!�/�����ίW��$��V�d�Pg��N0����y���fx��o/ ����.Dߺ� �{_.5K�!^�b�$l����˛:΅9�$����t�7o�Vdև�L+��f�����H�w5��4n)#��Om,�(Ѓ��M��: ��4ɤ��K��՗�.���ȃ��W�sP�7�@c���;��q�E{i �ͧ@E�"�U��}$��섎�V$��.�����MM�|FB��\G]|�,��DcѴ�����$�_�D�e�dʭ/���G���y���m3�T���]W�1��B'm �24�Ǥ8���V���.J�ጣ�x�`���ӗb�0�>���F�f�t���i���i� ��fz��ZkWIg�2�(�le���xxdphNd�	�YmE����}�R���vm	G>�T�~����x6��6*�6V��ҏ~W
�M	hB-x�T]��2�r�LO�U��Q�����"��.s���P�t^G� ��ejA����Y��zZrq�d��������0'�K��Mp��{(#S5���9Տ�u�l��wb�駈��-�Ȅ�;��1+e3����3��<�=�kB5B^eH9ī�]QGc����X�J]¦3������A�}��!m�W�����h�BO<�ٻPg���E���.��z�3�/pp<ۺ