��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�!��
��%Y l�׾����|R�b�@�n�?O$��5��z����reWL����L�Q l'�� ��a��%5��6���.�gi�`h(+)��g���L1�W���&pŶ�ϧq�ž �E� 3؈�L���_��[_���� �v���l-�.�l���q�clKR��)��>�r�D9�ҭ?CT�u��Z�ʁ��<	�I�*�@*��s�mG���'�F՟y#'�`Nq��:�\-�7�nQsu�	���s�_-��䞏���&i�j�`��+a�ܷ�֯jaXY�.��o�~�,�;� ����]�j	��\�/bj',v�%���oX! !�N������8��X��/�Ʀ$G���6Tۯ$68ȍ�L�>z	� 1�� $�nS�&Wz�"ia�t.(��i|�9b0+��A��i��j���LUdT�µ�44-j���-�oa ۆ�����1�d�dzlj�'��M/�������h�WB�r�������c<��b��;(���&�e�2�ʃ�Ƭ˾�z�X�'��b/�0���i$�<��i��*�N�AG�j��i�Т��s<t�[�.nF#c�SP��֣1��tp�'aջ׋y���i�΄ؚ~�*]��U�d��eV&���H��3��9*��M���ܯ�䒷F�X�w�>W�Ŵ���A�IX;��#�ֱ��^=��lנ}bV�� �3����8o�����BZ��@5ZN"'�%^	�,lT0����K�L��Q$�3���}A����]n��ko�9%�i�� �@���v8y?�����2g:a��6�����"$�b3�@(
S0�@��T��i�$�A�<d�y�*H� z�=UFXĩ�RH��ZD�xÿrA��<�(HU��> ��"���4g�愑�m����</�î�`�",�K��Bk7��܍?�#�W}q&G��E��˱��"0Ej����0_�83�OM�@�o�hD�-�m#����ˆCi�IP�%=�a�m;Z5>������ߙ�T��� |��8n�6>���n��%wC&V.� ��ѣd@K��ޗ�~l��p�~!m4�LoPRjc	 +RE���'��d6�6��N\ún�j8D%؃7.��}�)lr�O�+�� e�z@(�S4�A�!sȲ�z6B��k���������i:�`,J�|�e�h�ɏ�6��y1�e�C�9�=3�_|�0iu�G������3�k�N���㜍��L��N��-y�.�	/j����9]��h\����@�|����������40x����d�����E|�zu�lH�O�+u}	ʬ���_�n6�ޅ �o.�i�.!�;v=�xGgw`�|���"ȸ���=�e5X�o�~%�}�֐UJ|6����$'�d�C����z��&vh���[p�/s(+�i��n�2���O���qH�>�4�HҞ9�Z�a��7,�k
|4Uj�n��Ul�w�$td�"d���0�V�װ������RR��&�I3�� Y�1d�'h�5(����G-�?`i�$}:��p^�_Q뼾缛�����` �����-��Ԍ���w��O�<P
�a��'�VSI@M�0�g������ي�;�]09b��3,����a����n�^��W^[�7d���������V=��?��)7�O�_H���h�z���%��T�W(�Ura���l ��W
`��1��:���sׇ�߾lt�0�fg;�X��XT���-�6��w�jͬ࠙�u��(�u+�+����&O��N��x��7Bׁ��=#�ܫ�=�v��qQw������V7<Z�<�����W!��' )�h�!Q�,���8c�{5p��2\K/�Gxπl�Ϛᶧ5M.M��'� �v"�g��h[�t��0��ݻ�m��?��r�9o>i>~&0�{�G;(G��+���i�=�xQZitą��$k˹�'D�֟����|�G]b$v�������6$��@�Z��N�Xۆڇ����r����~B�wR�@Cs�c���R�j���@�Z�<m3�,=�5�����A�|��w��܅�S#� �( 3��Nn�c�����N1hp����䀦�*ش����O��k����L�>�j�Q�ʢ��I]Om��x(�]Rf)��h�'�b6_�x�0�O�/��"��K��-%z�w��"��ř������
o�r�+�Ǧ������t��u�&ZщGڔ���a��Z�dq�+x�?��(�\�f����f��իB5�Vg������12�k��Y����h�B�p5��Y�E�4��*�|2�m�iK�����0V��Q$k��E��IŒHڸDJ�.�P�����ּ�Z��/<�9�I�eݷhs�^�w�B�$_�E^6!�۱B���-�K煚�"Z�E�ۣȓ���e��{��z.������2z�g��e%|w�?�А��)�_�w�,�����\�V\#�]�M��P��ozB���FG�fټ�?�ܞ��BK(X�w�M���]r!_.���7�By� �~�H#YEܪE��p䝯(�2(s4�6��[�Z5�W�l��v+�	�AG��&�C���,%	rH0"�+�fJ���B����KF0>���\s�X��U#ai �W�wP��QY4}L����ᔚ▝�0���҇ԋ��Y��~Hб�L���Xg���R�[�'GaXBS�XBT@pe�<�/T�u}kg���(��B�~�����.I�{�ܖ˴Y��]0�\�V��p�"�X�-�?��������{\m!m�=hп<7-5C�yk7}@�3�庱�Հj��ׁ��}�S>w��M�|  �̟0�_a�q�/`��Bmg�k]�@��sX���HRu$��At$VՉy\n4U�
۪*8�2�b��u�� R�������t4�?AQ�ט\ã�iӢn�0ʢm6������!�L���➷��4l�,�69��pƓ�6ƻ^�y.j"	���xJ�cD�Eb�w���T��c���,FoB^0�J�#��Hm�n	�o��Mbm�^p�ڥھ(��x��)�����3[���u�;�%Û@�س�9�?T�����D\o~<�Q[�=F��EK����Ew�����D�*QS�����GL�Q~W�e������l������_LS$L�\�.ώ��eSd��O�O�z�V�f#�\��Y}S��z�>�Wg$��4h�"iqb���8;�z���i3��Ә����0�J@��)�F��Cf�vo'i+`pP��s�'��@�� >���$i�V)�c�,������[$��I���������7�Jg�'ǣ����x��e�ݾU���ӂ*�D��?��8��3o��87�0��/��iN���G�1�z��d7��]Zh��W�t�=�!&*E�EdǪ- �C"@���K�֧���d��3J���-t�����f�mw
�� �K��tm���`�Z�î�H�Vt���������n>&&�������M�PA�j��uF�h-���Y��A�(��[�s^���h�M�lo�veC#��.?-"RV5��8�J�*�uHJAB�c�8��2Ve"&�(�"�O\���	�B���G�1���c~nd\��J��̅���HkS����a��3�6U@;Jh>ݒ���u*���k����n�eM�,-��� ��8��~$H��^mO�<
.�K�H{�2�j��1��9�o�Y�+��(m���ɭ�gM���J������~���i���4��� �9����*�V�$�xʯ�l�,V�kD7�Vɤ���������/�ZӉeE��oQ|xxI�^�����o,�u���O���m���ˍ�;�Ӝ�\P�Gl�{5b�Z9-����h0q I뻣ڢ�e��z�c��|[��8BQ��	Pva�N]�.W���x��G��2r�!	�r_�6w�]��W�I��f�%�汰0e�ˎ�h3���d����c��
��)�d8|����"	�>B6�(h���T}��X�Ae*˵�$���Z��"M`�5@�Z/G�K����w{ɆVa��sbz�x�}�R�ρ�*�Y�0�t�Pq�<́���6�T� ܎��ඉgʝ�dB/Z�Bauw��D]�҈�A|$Cd#y�U���H|}�6��9'��#���>N���M��;;��Oq֭p?�/p���(7����v�L�]�z��C��TJO��nLF]�4h��1��o`�a\��ᛯ��ȳ�y:$1=���da*u�����~DɞS�ts�}�:Š}���?Z2o����/��;��&a�YP��������GY2�W�v�֡�x��_�J>P"�ݯ8�6smC�g����f��N2�ֲXjd+2Y\1�Kx*+ܜ=�o��*�r�E���2QN݌��Kr@�E�$O<ls�~�x����;�z�-{k��^|���b4���OWi�?Rٔ���/cV���h:�׻�'�{��N�k�PX�&��u<E�e��kY�����Ìp�˾��aB�T얛�՟��Qo�W�Ӱ
�(Y!n��`)T蜺w{��Hm�M�����S�����}�\A�Qq�?�q��ñ��m�DkȽ�R��E?��f6wQ���v��?��TRݜ=�F��
��n�tڔ�w-�w��Z�SpB�x왴I�T�E��϶�Y��G`�v�1�/��.Ͱ��P�>�N���'�<C��H��Z�3�U��\gRg㍮�)t�a���tG�����8�I���;�u�݈s6g�~I����A��)J`��a�ۗ-�2pߒg�6MC�}��w�����#�Et���� S3f`U�E�̚_�L>��En	|��l��u��JMI��gۻ��Q�_b����
y�k>�}��&���g���_�Bf�"	��Z!C3i��wV`g�&Ic��x����(�(s�4�J���)YC,��P��vH�_�w��^S��+�����)���;��M@%��"���f�n�U7}�nzQ]`�w���n���$u�&$�J:z�\G�D��"a�����E�0���u:3�O��[E�����v�j������m#	�o�uŒyX���G��>���:���6�o�l�1�7�A���E�s�X�)�������`p��GE��Yz��CW�I(��^����U��s��%˘�!0��̽V3?s��U<�!/�erh�q���$)��a�59"=FU�O����R�ަaZp��8R/�*N�4�d��p��\
ޓ�Ęe�O<Lf藟��G��DD.�1a���VDh���
�w�!�Y�2���x��]#En�|xʟS�5/�u0�$'&^՜��C�7c6����7ko�_M82�>\,���}<�'^�Q����X�E��2�\r ��Q����᭗�|��[ğ�b`c�6�K�x3T߰(�M�Z��O}ρ��b�@V-i����Bt���M�7���G���?�5P��%4*s��Ն���eXp묵�zAr�, 5106}�D[&�oLK�e�ҭ��̣��>}bi�e������
�Ǖ('�E�1�|��`%rg�.�{%D�� �.��*8�N~����`5bH3�Pq�{Nz��VG*r�jM�p��p��S��5�2��M�L	�t {��"�R}C�������0b���ʣaӪ�C�!Ư��J��̳�l�����~��{��CG��)µ�E�f�QP*�����-��4^ŧ��Ԙs��?@������yʁG�`��-ͦ)n(�5�	}�h����9Tn�+C��=ؾ�!��9ײ ��)��A5�g��n�:0�E(!E���P|b2T묊*�Q��*Ef��xirH��ܢH�xp7�U5��"r�ڏx�	F��c�s5-�#*�~��1ż������Ü����adw،"w�����R-���V���q�F�M��#�?��Vp�=��@�6�� {�����������v��NM�.��6wj$�+;��޿H�*/>`��,䀘C����*h�������8��C2�L���S�T�fqw����=�.���&�җk�cQ������x4��ô�����M����㣜װM��[G�0�IK�3�#>l����p�\w����w��D~��fqb�������a+