��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�KW�UHս�K�7b�^��<{�+LP���E�[��,LUU7��o�9Gj]>�U7��w��L�s3~/�E�����Z���1�"�pK���;L�P�����^��c�f��5�-���j�x:�Ӝ�,o������zi��jWvs����hT�)h�����Ƭ2��|�l���XW��PV�cJB���"�1�)��F4�P��,9��r_�o���!,�!������ʼN�BӸ~���;$��,=��[�u����s�U08��
dѕ��6������Z��gLU�ˎU��ϧwO���DM/�.��j�X�;W�Y]H� ��9ߪ��c�X�Su�K�����C�UJ�?̃��XE�+�}��	���[���C�V��z��!VXNF*�.@uL��Ms �$���t����^�xG�Тhţ�����+x�p=���I(y�D�#���o/��I\����fGuO��Ũ��fA\!0m�Ģc��&d��VN��3����A&���e�m+}N5�+�ut0'�`�$���_��������k�U3�헳�M��䞵�ң�:� �l	6a=���)�`�2�~���]�tݙ���,���;�2f�r>�&�AJŨ!���B��&xL�:��[�m=�,;��*Wɕ�l�m��Һ���/�p.�_��p�&��Z���2:>��yI�f]+J_[�3��NmK��$�oN)0|8�~�f=���똅׍r�:0�αݓFy�u��.��_�D�,�m�9C�`�QA&��ٯ��+����Ќi��̹=/o���uK�:��)�N��f^���c�^7�L&��<y�CM�X[�_�%Ah�[�*>L���Ɗ+��\���`'��o�x4�:����dd��ş�)''c�ܹ(�i\�qep�7ɀY�u��������Ǐ�o㸦0�]Ѓ!\��H�BMpm��5�Hdf@�Q������#��/%�s�����U>d�F����)�et�z�Ő����7W�VNo*<"mՆ֓8Z__��Gz����[�h�����LQ�4�������)��Rt��}�IPss�9��Z�9�9�_�*UZ�5���E�1]����@����
N
���ݾz�Gꤤ��R�0��F���vgz���7��b�@O<=�~nr)��qR�����V��]�����=�bX��?H<�:����2G]�Ҩ�։��rT��
�{��2D?��W����ֵ�%�i�3�_~�H���h�:���M*���G����V��
י��~d��nqɎ��f*�}p�x���� ��xvN;�Z+A�S����؟��q9��n޴��vfu��=\��Q}(c�r���!=�^
����M�� N�h��>�`�<��1VT����|b^|c����!�+��z�7{F5�ձ�aB�-I�nR�0��J[���b�OJ�4���>f��轄>>N��aC]k��sҧ�o�CW ��q��$�4Y#�r��F("�:���v�f�X%�k�	IX�F.�����/7;?�t�N��jb�K*I֦D��o� �Zџbcy��6�4I��}*���Q��wU|��Z�kh��mOxf��!��BPJJ$�����������k 1y򂴿��@$�j��)�<��J��>6��,�s�q�=��Um��6H��Y�"
?�\J�Ș�q�+��a.t�����qD\�1���d�p�s��B��Y��_�	aX_�g
�P�2Z����7)��k�6��X�Z����_^�-�#�`o��#�k�������u|S�^���N
��g�-�}��F�ۯG&Ů������+{�:��Y���K���N9�S��\m^|��<���X�)׉�[`7���d���q���G�U�v�5j)'\B\��V}=r7�	+~�s1�6EP��ЂZ��K�!�����愨3���囨��G�xɕ�34p��*�"�ps��]��ʴ@u�7dȣʐ	��[*�A�Ӓ9(
OQ�O�,�R������c#�gԣ.��Z-B����!{'=0�{M; �(�<�I]c?����7�Ð�5E�L4#ĉY?��_�.�H��N*�_�O7�2���T~1,�K�� f�߾�`�<)8l�q?[v:I�u�
� {��fO^q=���C@��G*���zDu�z��A[��>f�t��W� ���r��d3�C�-�t�d��՘و��W����җ�Җ�<i�7���1�UJ�*��^R��)��=v Jh����@���/���kH���ؼѴN����ʐ�w$��.RЉo�y�fq��T;���	��J�Z�s ����9�Nk�J�<��Y�u!z�jQބ�b�e��:�����g��K䒛8�2�װ�X��E F;�U3F�[�,0�eO�9�RE����HW�f���0�����_�6��f�ۦ��m�p1�y,����{�ޚ��|Ծ���ō�k�o�^�}q�m�_��Z-
II��F�	䶫�����h�ֵ�����V�����$��'�#n�V/�L�&ISZ��J���ha��C�\���;R��c�hx�3|��\�'��7=�[����aE���k8!��l��3[(_�]�Z�N�֞��Ȕ������J8�Y���quȶ$o��j�o���C-�1��`�%�*�:;�G=�xǽ�W��QD��}{��f	<�Yak0������Z�vr�q�m~��coCnh�S���\�d��4���3�#�<C��<�:&����m
�yiiv�Q,şl��Z�J�f��O���wD-���p�;P	υrK��D�>
N�����[=PkR��.�BO%r�����cw��\�Ӧ�����	�r�X[���S�}��\ޥ��c*RMk����b�U��$���;,)�U����T����}����/�Ŭ)����bZ/�?i���`q�3�Bc'�l��V�>z��5�jj��cx������>=T�3p����c6B���~�đ�+�.�U������=���K��]��@��^�69��*�l�����J��P�׽�S����[�
o���֕�(����m����z�"��Wy�>�vA!l�k����ZSmv��l9]M*ͷ�?�3�V�rգ�gC�2 �N�]�� o�D{MEy�8<���(�^�-�鎁�Q�X)m?��<���|o��!�aHY�G@�4�~�j,������	EƎ�U�N*��]��t��/�����0Nq� p98�ϩ��p���e�zO̸+0�ւ�ڊ:Gt
>�w;ъ2����qN��m���������=�����i��v��\�/��f �T�T>h4W�C�z�2�����,��7:-!��tX���#�|�HV��Kc6-��QυZg*�1g>o��y+�L�`Ɇ �Դ~f~����LA:*8�������aa��B�$�>mM@�}^83��u�N�W��v�
�+�W$2�0s'�{��T�ZTJ`Ov�?��#��?�����B�+�����0��;��'Ȳ
ݧ4G�Y���`��e{��D`��F��a�2֝���S��l�� ʨq�#l�w�w"��yQR�zF%�������x'�L���o�y6-Li�H����&���6�[�wH�Io ��.��݄lyy�O,0I;{ڗk������D)�HnȈ׭B� ��Ӡ!N��ĕg����_���]��]U��
E�farZ��D���lcXO,����:uH ���zߨ:߮���_�!/��P��%�p��YQb9D�Τ��kv�ն��u�T�Lx��9F܋n�׏����Y=�J�-���?P�(��K�y�*=0� A�U*e�����	��O��&�ȟ3λr,��Bp+ʅ��mF\�.<&$�%��)1�Ӕ�7�%����S�4�)y��=�w�@R��������Q]y4�c9]bbTy�~2���S��!�3��eU�� |Hۙ���M0���Äb�G�xk��*�0���zR��b����d�'.B�UM��ϋ�pi�0�i��6e�iҀ\2�&sJuz��bH�=�W����Ƚ���{�g>7��wm&��9�b���±y�����jov{0f���5���{�V�*1U����1�<��,�63�|��7���/���G(C��0�T���!��)J��T�����9������`�����J�:���x䣺�]'z�� ���������ڧ'�u`������眉��%�C��պ�y���N3���+�h��~txCݏ%�5Uu(T EJE,�^B�7��
3� h�Z7���&|�iC��m�dc ����蚼�*�6�<�*VM:���T������r20e���(���_r������/vYM}U�IӴO���'~�W�(�s�e}��z�I13`�&r1�+l�l�]f�G��*�H�GT>�mʹ���S)�Zw����L}gNz�>!�f3��9���v�����S�W����B,|��V������9_��Y�}8R�T�X�b�GZ0��M�~z%$@ ә���雃�Ņ�s�<����g���J�9�w�m%�m��48p��Ȩ��+֝=�5�=�tH��8G�����'ҍ=��:��A�B/n/�&�q�>�fk32��~[���V���U����bMΒ_��1�)�@�N:�������=��8�RR:�`�O�#��� WE\%)�B K1�L�J,�����bPy�}B8��@W��w��&����1��%q���y�]!�xж�7J�ض�(�����Я5-���NX�Ac����d=ж�q)Ӯ��p2f,&�JE�u�a��hfG����{6� �ɞO��a��������nj��� -QzKaEʩ{�ަ𘒏��->�w���5`Z}@;�ae� �7bD�!l��@�e~>9��}�1��u��-���jC���j�f��>�A �P�m=k�jRB� �M�r�S��c���u�&��'��E��l����}���� ����Q��5�e���X$�5׍$�+'��MD�a�o?�Z�U3��Q�)D��.P�xD����P��Qܢ�@+5=��N��5rBhCd�[�bm͹~I��6G=F�T˱�m�a��L��zk,��?��N�ǔ�%�`!�{ ��t}�۸�ODR��������^eiȫ.G��/\ވ`Ρ&��=��U=p6}�P�IY*��e�̆U��W�����G��~���9���%d�n?���B`�oG{~HM�X��V���FL���O�:!~�"\<��i�:�̂��$�;�kPgy���yY~�]5��-���w�L �<&.�vu�w��fP�WY�����L�ֿ�a6�/WC_���_4Z9V�Q����Q�V��'�"@X�����w���8~�il��Y�~� �@MG9q�O�l�����\��z���7K�r��Ps��\�t��c-���1�;�{$���m���LJ�##	@��+�����3O)���!����h8:�V���wF������=�#�<�Hw�@(�}����	c�Tz~�K��v?�R݅��f,�M�ڙ�9����R�an��Q�G �����\I�/#6�>c��W�0�>���\�#�mߺt8^���o)�����h>��Ck-7����S5@�`Y��c�27cqqM���!MIy�w�I\�j{^q8�Z}�B�(��'7��)�5��CCt��_��3������������,��fؽ9"wS�K�-A�d�B����%�o�ث��)M9�@�a�:��sm���`r��)ΐa�T��4��U;|� �od�� :9��I�͏HH�R[�>��o6�x����D��O�L���l�s�`^F
r0�wr�Iu�@��d%C��J�k�y%�S��:h@�5�ǡk�@�25������S�v��֬8 Ra�Ti�3U���T[�-A&9j�K�5N��1L]���apr�q�n���U�d�AUY�1�(��@J���-�jQ��e����`{},�S�A��h��b����l�-�Zڨ>��G��n55�ۂL��|}��P�-#�{�S�h��e+���]��&��֊TU�&� �3_�)12���}��JR �x��s��y �L��J���7f� ڢ�])�� !�ϡ|Mc8����r�Z�A"z����dR�Q�(��|�JIl-a`�^�m�%s��/Q^7�؜��Qf�Z�6�����F�/<�/��c�a�T3)X�Ԯ�����K��V?�qj�D�?)�R��W��j�i�@�%�(���Bp:@�l"V����^{v�8��΍̄��x��C!�v>�����>�71<�%G�g�>��i��Hy����e�R�/�ԼÙ�tVZc�� ��C+nE ى�Jx �A�S�HY�j9NQ�aYY�R�fF���϶,����^�hJ��T�N�w�~�\\h�:� �v��g��S�ʦ?1�|pϳ��-w���ܦs<9y��y K�2�;�>Qِw��a_�]h�ʟ�ї�ۙ;iV�Dz{˰����~�7e�S��["������Qq���DR ��PB��0��n���z��%ך 0_iS�:�S�Y��R !AƆ/�$�Z���69�S�{[����y!9.҂P�qk�M�`H�H$C`d_�&�X8��"��ئ|<MMpFܷ��(L,��Yк`�e*N��a�ČG+���u�}�����	?�z��-�ahm���7͵���A�"/d�mϑ��;�W=ƁS"�+��߇��,R�T�!WcX1���D�e���uwk��TBuY�Xp�Ig�фu�W����o\����$Y;���<)!D� R�Uf���B���*9�p�|���]͆�B��r>�E4�0�ga�i�CW�e�d��@�f�ߊ2<4N2i�Ѡ��C/<)t�J@ �,��-x�YC7�O�|��XF\O�d��;�? LH��j�〱Ri�%��qM� �k�<$/���F�|̴>���aY����Q��,bԁ�_�\6��׸/�W����7��e�AqB�bO��gև��JL{�9�hrc�����K�7�tF�C�l��h��>�]6�Y �vB�Ra�J�D��O�����d�h��'����T���<Yd�7΅u@î�(��ecGM؋��R&9d O�� ��>�o�뮙���u�5³��ײ�Wx�y>��+�9d�A6d®ȷ�|z��cs�o�Ra�8,����?wv�zZ����ns�t�ylF趬� 
h�5�U�-:3avQ:�c����Y~�@=�>~���<�}�7G��
�iz���xB�Ģ&�-����6���&�J��㢲U�^���*�j1&; ;�3ˠ�q`d��Љ���M�A�(Z�8�`�d\�&B�WAv1 /qd�-�A���{�[	�S ���X�Ta+���
^�N��L���ﳪ0�c/�>�5kQ�t)I���p�lЭz��tP�p3�6��a�j|I�F��NL�F��-*&�	�,1]�|�����+�TeuC�5uY�@�rq��Xs�]�a�
�jxՓ��/g�Ja���pY��6o�����/nl$�f��P�����S��xv�ʃ��2���:pW�MX\�n��;������K- �C���5'o�o#�&1WtS�����%L��$���Q���!k��}0��:����N�xFzd�O}�q�y�%���n�I��<,N��-\��(�+w�|`��+3H�J(b��՝�G��	^_���zV�����2�x����j��FE�#�Mĳ#�������,߀���!|p��yə�``�j�%A����u��� Ai\��� m>ܪ�E�F�\"�li��Z�7 �H���I�R�+�g���(4|�p�p��Ѡ�J�940o��3\=�n?�?ipU��L+����Q�h����cfm��*��v����I��~Yj��SΩc|��o���HF�em 3U>�=���H_��
����C�&gG%�Hq����� �wP#��6OAd��'��I���)�����P4�IF���(D7fc��5/,�[�֒{����<���u\����J����-����>��-d�@���߾�+.\�J��e�A1�ԛ���Y���ZASbM��ƱA�#r��Eϸ�bm<zMt7@>Hk�.wK���Y������!��<������R�j��Z�l�p��k0iA�ϮRR�Mle���a촓�k�;8�J���]�.Lǭ��Q��}YO�G����2����d�T�Q&�a�d)Sb!��;IoG� ��b��0���ˆlӥ�*B3>@Ƚ��ќ�PJ �V��ĒЎ�a�zA���9	7Eqkk�i���O��h������=%}�/�"s�Ny��V�%����������������4���
$^A����T���j�_Ӽ.E5��W�ۆ�BG\�]+���dئ� �.Š/�â�ڙH�&u���.�S`v<���p��� ^c�|�Mo�%��ue��`7Ow��i�b[<��.�-&U���,��,�����8��ra�
B
���E�:�Ȁb�tl��3� ��vg�R<o��N�M��)�����pKW4DY,׭b�q׏bj� ��w�n����Թ%uG��GP����Oȟ�];��N��zJ��_��
i.����K�����^�g�]pI~���8��'�q���P�0]=���T�2]ق��>�?�{��d��X|!]�I�p?�`{)����a��4���[�d��k��<�'V��T�Ս��ˑܛ�Z�X8�^ر��gpD~�,��DL�[	��u���=qM7����A�/��5�����D��De����TI>�٧1����~�!Q%��m=U�;�N����-��p�q�J�@PK��W�����&h�Z`��b���8�c�>�� �ڼ>�Ԝ	ޕ������=qj-�xM��I�0V��/ w�^�����a^�!��d9G�mA������yBu���:�1F��F͖�M�Wǿ�w��eV�1	4�:��]���W�����KD��nio�hWBA��1VX�*�!�dq�$�U_]�5rk-���M�n%˷����I�v��zw\�ǂ��V����3��'�'��c�����{!�p �[���mԩ��ũy��3�Q`͡��� ���;�vV��G�b��O���>�
|��Iy�{���JQwZ �����j�&�a

c��X3�h�ՒV����I�'@���ϋ�7D0�2�֎�>���jMx!�y��7c%1��t�T%�Ŭل�g]D���`�����]F��c��}�`t�n)�u���(/7h�ڠ�U�b;�aԅ�\��c�2����N�����E`!��,4�О�a\����BM���(�qCn���`D��=�~-���♹�s!�Um���[�`,F���N�P����[S�g;��}Н�A,'�q	[�6^nPD��HW�#�����~d�<8������7t��Y�~�>���\����w��U��^��A�+G%v��JpL�Cc�y\�5S����b�mi�Q���� �������m�e�0qtO#�F⽩YL��l�vB�h���6Z�\U|��ԭ���N9��xԂu8OjGG>f��׿�W�E9���s�!�T�؀����H�$�H������b�wNCW;�[x�v2�N@~<�k>�Q+���gR�
ꭈ��'�8�k#h�j���ZΫ��-}�����({K�w�W'�S���H��StY��@�S�xuU���]�u�iZj߷�ėE�ů���;Fk��FmY&p���uw�"+|�.�?(.�O��njY߯�Y����NJqBz�� �Vb<?t�*I��ʨ)��X����j�o8��	O��Y�M���]�~��63�D�+�!���Sf���p��B9	z�aIF��lُ�Mj��&]:�!O}Vlqk��j�4hY��a�s�!�N���t)>��&�������c���R^�Ǒ!} �C�
�ؾN�g`CJ�q���M9f?�|W.�}�POR>2��zTQ�֎�W7uғp�Է�9�����Ӆ�淢����k!�N�/�m��֛z�������T��aIhm�;��s|`��dl�v^ F�t�V��T����<�eiIlA�~�>�2frE�<�Ea��T;GW .��Į-Y�L���XO��Ơ/�_wǁ���iySx���O��$qʷ�zN��4�@g��zaBs�R=��/ԾQ߁�^I�d��dY�&�y��]���[&D�Y�@͆�pj5����~����<^�O