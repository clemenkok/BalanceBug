��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�!��
��%Y l�׾�kqDL��y���O�ɀ���Z�J1m~+�O+��L*z��S-��
�-̕�+�%|Mѽ���M巙N���[���ݲ�W�od�D+�Nl��p�U�OQ -7���
��w/o��,A�wۭ���'��	c���*Xws5�@�����0�l1�	i�G#�¯f'�,YƆ��LP K���a��d�����X���`�չT�~A+�1|�W2Y���u_0����k�<6<ۊ��#M�����X1�(�^���iR�\ٗ|����zjsuH����~Q�@�3	=�/��z�u��:�w8	�d�֙��:c�3��U=ؽ&3�0�@�h3?��p���a{Θ��Fvnk=��^WZ�� .q,����km7i=�@������%7�=P{虞�y'{�@4��Pp����BhV1�d�3.艡�a�@�?o�F�_\q[�EĚ�L�y�˜�|�x��'/4� n�s�
�]!�G�Ɉ׫4��\�j�G�A�d�y{PN������)�
���4!���O�U9j���q���X�)G�	�'k���A�d������'���9au<���(�߿5��+��i��9����|�[_�

p��Xa�z�]C�r�(X]|��I>����U��.+x��>�$uHT�t�C��0/*E����J?�n�JH��Zlk�y�Ê`i+�����o�w�.��Xgh�>L�[ ��ṉ́vJt�����ṵN �c��*�Tg9�'�-�;Z��:;ދ����q��w�����k�<7�s������σ �Jn�$;�����D�z����Y]����q�+�eI%E�-�FO�λ� �灞���d�3��zfW2[��q	�>�SXQ�dާ�'�qԙ$���߀�q�j�Fo�Δm�u���I���*lw�v�o�cJt���E?_E̵*ֱ;��q�D<��q�mR�R�A��>�DG�����a�
v�	��5�o'G�>��3w4���m�7�5U�tӶ���s��� ��v��4:�s���!�����< bH��_/��A�������x����	��/�C��G)0�Z./�Y+�Lɕѹ��:��T��i�L59x���ʧ�r7�脥���7&��o9������RMz� ݹM�S|��br���s��~��W'��~�A=w�	�	�q�6���i�c�{r s����@4�u鉸ؿ��y��^~�H�p��>� .t����\�3���{��oX�ߌ��Acj"��?���uF:�c
�`���+�	em��kc���'�9�#ꈔ#�����p� T�`��D�H^Wؼ���4Z���6N��A�)�O^�9�G�� �̘d����d��Cs��&+���p�)'�m)���m�]�-�3v$_m��䮄h����M8����kp<1,,�G��	�ES�W�i�77;{������ ݘ/I��c�j-�k��6A���k�4�����p�=F��T_קJ�c�cc�]tBt�0U�1�u��U<]d>n�kʧ}RɗdsE�QW�b'"��s�b��@JћT *:D�j0i�$9qN�q�{J�b6SX*��;VҫZ��bǁ.pɎ�/������	�#�n�D)FU_����6�(zN6����1��l!���Ow�&�BZ� A��s��
+!��Xm �+�=�B {���L,s�ڝ�?�.U]v�WkoU�d����
�h3;ח&8���qO�eV	O��r�TX��VD<���.���M~���-������נ���~���d�B�]a<[Ci�$C]���N�҅벹��4��`�\e	x���c��6Z��7���CaT����)���T6�G��!���i�c�b���l���Q�Y�3Q[��u���|�H�UR�x��0x=>��"�J�E��[��VC?��G�NtUlw��9�b�W7��]����ޠ.��}�NОV�~���g�7�6�?4�)��M��d�-�4�mrg�j�\�kbǞ�g�E���ܚ1�E�@* �aY��|@��*^>~�h#�m���V7���5.T�Q��kR�|��UE�W����5v�����nO�tp��ӕ�x�a	5�`��[��Vy��&�t��!�KI/s�5�6'ǴQu�D�����,�1D±k� �	B,ף���<��Q�]7��!����8�����x*�ŗ��6|^_v�̚mkF&�W�������i/| �U��h��I�S��9w`�pG��i ���a����b'
i����l�dT8)+����ץ#H��p&"Ԧ��=���h���Ǹyɳ
�c�#�K���zD$0��ܞ�M��t�""9����zQ#�v���e%�Y�퀁��rc�iR;��K�^�a`b({Zg�Daw�#UhK|rBF�-ڨ�D��iq��P �`|[�U���?���8/h�
^��� �z\*"�Lݻ%����Y�)��)�TG�v�Ͻ��ߘ[�x2��
�Ro�DI�ga�WgT$�m(��E��O�Y$X?�qB�Uj���q���*X�Y$� �g�M�������_�S8�|˥5�C��}:t� R��wT���cؒ���ٌe������qO���e�J�8�P��>ݽ^2&ovg�űۑKzZ�q���>3?��N��������(��(�����k��B�+='�ڶ:�A�5�=)��P�V�)���	��}��W�q���3,���q�F�E�=�����É�-�^]��T��W�X���.��n�ՀB�D�2"����ؖ&�	�
Q� �m�0�"�:ƃ���;�����E=� y��h9#;���]�T�)���Iy(z5*�GL���U��ߊ����/S� �\�PA�0-��|y���_;J�Y������g�6�&f��2���d[ؽ!TS_��E��V�U ���� lp��9����]�a3�E!8$M�'��t^�hTUX��@$���F�kK^�ȶ�_
,�
�.��_����M�,��z���ӑ�=:/���r�E.����vZӼ{�J)D�`���U�xi�Q��&�XA[��S���.�i��h_#'��5�o.ΈC�Ϻ&H̛a�~����Y�3;%U)X�9ɬ:z#�����: �--����
���DtAB'��)�R�QH�@��V3?'`ٛ1��T�^�K�X�?&��~y�4�7|�(V
�i,�˭3y?����mZ���lRs�A��Egs��Եw ����Gert�)HX�.5��/�|��P
�h[	�d!�B�=�9�1�����C�G��{A�A����˒��u����u*��f{2�
����6a���D��
���R�3�z��� ���� x�};_F�9���8���2��m��й�],�>hX[4�
�w��]	G��~\OU+#4��n	zZ��2�؋�#.�O�~����AAm��U�W<[ä�o����0n@�Q;Lx���x���Ŧ��\`���b=�;h �]�4�Y���4�N3\�wN�ɗ
 �ʛ�s+B���z����=˵��F;d��*hp��|#G1�����,d,�f�eO3], \���4�Df5�è���H+�l6�dXq�k����j�9�Ē�Gfmu�7���Ȩ�I-ƃ;B�=��\0���3�THVT�w�Jİ�� �	�	\�3z��Q#j�B��<ą���<�o�iW��֣!��@+4�DqcQ+��F�D����O[���j�d�;�������dp��[}��)�:s�\l'�{D��ǓΚ[����_�t(55�	���ȴ`83�`Q��?��,_���Oky�(��"]8�PFJ�r�߲�����J�Ӓ���Ur[��7��?�z��a8y�ÀPZ��Se������:��,s��%�|��r4��A�cQ����\�c��BVuق-�ؠ!�]̭z��9Ų�
N��x�C*m�������p��@����ɥfڰ���['����^&!�xn�Q�#2���f�Z�k�2���H��-�;�tyr:D��e*![��q�lq�g�)F�9�u�F�����Q�X�9���YS�dxC�P����_��dS��qP�+��#��4`ah�/�K1���P����*1���-5c��ǧTý�˫���1�7�jUC�fI���݂
k�{����Qgv9�X���)��4�&�DW��%E ��<<[�W�Ծe������d6F���uE3�T�(x����>1]�72?���$8�D��+�؞�wO�yMJ2��r����Z���o?�������<�;D�CxG�x�����'A�+7�W�����G����@h2��ۺD.�s���c'd������;��O\�C�U �{��T� M�4]��_	��΂���-�ʓ!�Bqw3�v���Mp&�`?��q'כ�����[��a��x�/�$g'��Uc�#�\+����ݘ�9Oͪ��i�L �ز\x�j4CٳY�E{��߿�1�o��������A��
��;��R9p*辷��X�7�F�X��G;��~����3��F��/v��B�9�׍3�O����>��XMw	�
&��ɭ�.�]꣋A�� ��<�J��Fp�����2J6�G�.������"N���:a�#ڏ���]:eBj{��mj���|�:_�^����t6��n����܆o�p��NLR��
�;H�p�<��K�!��j?���z�W�������%[5��v1��s�Cl�����I��xӽ��H�Z����������Y�ؘ$Z��O�ԫ���#�<�n�	E��D��j*�7�y`�Z�aƷ�(��~�e�oE69�@hKd��bMP���ц�Y,�iKL��ӉX����fJ@��G�Ʌ���N^XZ��] �o� �i��(��qS�Eք�P�'�p"a��N��F)����,h�:��\E�`۝S:·D�ߍR����3�����2�o7$���.�i�S��Y�~�ͺ�j\sj���TMY��#m�KЋ�I�Rq�ˑ�Y�1W�Y/]x_,�--�0���.ZC�:7zp��󅙾�i�J�����EX2��G����L���J���#*��I��Е�U{��B�˂�|���^�LPU���ˢ��Y��|FϵҬ�*_ysw8�R�|	�H�p�t��6�����>(xdjQ��ͦP����M��+���P&&y���ܲ|�b�B��j�P�/���}
Ji��b���j|�$7�P��Kf� 듴��)�,C����$�Z��T�ohǜN�tVyƳ3`��C�f>�N�0uA+ ��Xk^�K�q�����.����(/$�Є���8h�����C� WrD��DP�z�6dni�.nQ#����~	��ػ]RR�~z�g��Q���[��}��e�@����zH�4@�����Ƿx��P�I��T�lI��Gt&aI"��Wm�dIj��mɄ��dU��� ����̄5X�˲�#HȾ8ɴ
Xd�\!X=�R�K1.�z�R���&�cJ׿����F���@�kz���sÆ^a� Ha��;���3	[�n2�T�A����YM>3'� X���u�������Հ� j���;�cu*�'�/��7�A���2��Q�����ᆰ�?�yf^�tp�8�Pq{��Jw
F��o.�R��7K ���l��8���)h>�@)����8�t�t�15E�o���~�����{��,��������h��M̹X�޴���_��OdY)��]���)-� >P�����hI8�j�-��r�e�����i��97��|�l�8b���Lz�K��+bh�<�N�G��V)d6���@��u�o,�؊���*���l�nv�b���d�/��������J���j|�x�G%��z�!�5%�t�P<N5s"��Lz��!���x�������͉0�G�'�K���~�6`�J�@�#7q qa��(�ʥ��"~�ȓh+�!~�F{GLW�{p�E������ج���Tl�ٓ��9���]��^N��H�M����A��c�;�ˮ#6��k�{MȜ�T�Y�7�5yWZ������b-�+!�mb�!J����>$�R��@�Z�g�>kvLњ̱lT�T��.�a}�ٱ���XOX��:<؉__/eݔ�����h�x�m�[�B#M�������{찃�&@6v���%�?K�����.YiTp���%����sD؄8��x������؈�hP^[SP�+�2�ƛ���l�Dk�6���o�)k�H�hu�_:
���?�H,�r����,��1�G
�Qh�}�K����T��ے5{��B̡�r�,b�GdQʧ{�-iB�>]a@4�46�tV��)���<PJ �c,͌��D�r@�)mU�7����w�_m=��4�byf� �I�����p�8e��$�93l"��r}+R�L@߶|�Dw�1ꁠ��sQ���f��ɐ���>Y�����|�گ�a4&E�}{�A�<�(���	���`��_8��ֆ����W@aK9P�nQi�=1���	\wm�y�%�T�;�2@��P��+�#d��u��&��Y����5��
Xz6�K3XQ���Yk@�����e��;Tʝ~���Up��ě�2�j�*�4�+�ܠ���AT;{Ռ�x�~1Z�؂��9k� �:6������������J��ɤ�,sy�t:�VX��x��YS�v�J~����X����ܷ��?���'����Z�4b�
P:A9ȷ[5�'%���]�����y�T����"B~v�<>k�nԦ�O�u��J 7J����bl�_K{������U� /6��.�%��w�}���L��F�*b����敱ٱ�L��̗P^�'#Y�<9��F�KYߊ�!��5X^�Y5E�
FM�H�,8�;�,BAq7��_@�i#���My�?���]��)\���'��33x�g�%5l�<-���
S����ek���|gǒ�u���z'[�݉P9���B#-H�˅Xz�Ӿ	�#��u�zI���45��O\+f\�׆�����O�x���fj�#;���+<��@���t�������j(a���R�m8$f`L�V]�І˹X �N�|�˴k�^��M�����[=B�4e�E��B�k�7}P;&�/g�(����	��ke��C�^���\�����p�I�Ճ*�'<��(����\瑅~\��� ��Z�Ȩ>,�a�qL��+�Y��)�#	��GXGx�y@��X�w �"�1�ʎy��5Vv�?�4�|��ZA�wk'B x}-I@O-Ť*^p���('�� D����ud�8�s�t�ds�a,t�`����{ֻOO��Oi,��'���\?��:��.�o3� &zh�������P����þ�������y����H�S�J\`�h�-�<��1u/���J�|����eV�.���=�5%�0�G;b�]|��S�t��;}���Uk�N7�3��[
.�y8В���[��x ��[�5��EF�Z+w��k����g/�v���zSTX��YC��_��%�cHx��8��,p;QKz��"=L����>9iϧ)���{��bH�N�V�7�}l�&�:�_���H��@.%�����4��<蝮0��y?�㔓yQ&yӜt"�����쌚!�̀�x���V���b����I��*��Q�{���b�#����)ߊ�Xjft��nΫ���,�ɧ��]�~RX�@��OX��%�� F ���%�����w�N�Q�G��Foq��;ُ
~x)H���T]j�a��OR�vc6�!(�j<2E�g�A����)#ix�tN��ۇe�y�ˆ��4���K�@m�
G���8��A�n��Hʎ\M��hǖ~V��C����h.�0��N3~��dY�qM��מ�W�e����<*�1�-�*�i�`����E��Cl��6�'zC�XKW�-4`5�ժI}K�Vr)朡�Y�.��	�����+�5�
㧶vkM4)�z�����B!�M������ ��{���yKl��єM�!C����`+��1q��(E]4 Z������׿�1o�cB=�rZ5�-��o���b�Dp�Da~Q���x`s;-��2؄�����j5ͦI�k�{Y�`k��[��C�e��w&�!յ	�P�E�)���" �Mn����q��ATv0�wVrB+�z2_�`k���O��ү�>��f#_��a�R�؇#���B���C��>��5C�U�OH���(�h��q���US��u�v$���$�,g,�,d|,�B�g��QY㕍:k2�������(w7�q�dNb�q�������V*����L{����ɳ_�nv�U~������M��T�5�P�5�L:5��U\qž�c��m�ȭ�ic��$��Ӿ���i�!f	k�EI	����"הN��(��ia�P�F�py��M
UW�y��'h�3)g�N��x��l�����"�+��xr�{�ݿuKN�bg`~�j
�0��C�%�fc�O^���K��,�]]"����J���:(���qr�M�фV�A5��}�d������p`�D��0Q�x#A�ؕ@�͟�u-�+���P��L{�^K��1�����%�=)÷��Z���1�¹:�! L��7�����]+ZWB�Rm�͝.���~����r7���hr��`�{>;�>M �^l
�\h�3���	�:��e�.��+��EDaJ|�I�:Z*F5���&�s�\���%D]��PS'߂@�N���,)��6����K{�����R�v4�E�]JYWͲ�N�I�F��Ґ���ir�1^��`-N~X�"�.������6B1ʏ *Kܴ��Q��-��XOw=���ᠧйT�=o�d&ˮ��Hym�%�FXsX�5�}�N�w�=���Ld0)�~D}�5xi�2�G�٪h�� D����3�������&&��b�b
JJ�v��o2g����?qW"�q��A@j��i��	�\k��/C�7�J��W��1Y��o:��9ҧR쭋���4Č�e=R���M1OӺ��'B����v�R��+Ș2m�]�b$Za[I�	T�e=��٨����y���l�r��+I��F�?���c�,Ηbմ�NIq}��G�����"�_���:��e \�i4�kfz�&��Xۑ��i&������Q[�-�l�O��N5�^|'�G4�� ����{�T�e���ռ�����'�Ⱥ'n��pW��j\&�]ԧ=�� @1��e�h(�����\�<��m)�`#eK�u�d��#f��1qb�8�Z�?����G(=���x,4��
�5y($���{E a���C���D
��nx˘����zCbh���-+��.�2�;��{�Q��Jх����r�H8�,��g
v@:S{��mbM6�[���)�m�I���s���N2�*�V���W�stC�m͙���D�\��܍k<�R-0�X���k1@��Fz��[4�{"