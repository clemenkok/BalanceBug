��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�!��
��%Y l�׾�m�F��������2�p�D������c|[�Ԗ�D�[5-#�ܰ|���:�mՔ����.x:��9�pgzij7�9���<M� �)��b�Q�o�28t`4�&Fl��ݚK���)��Qq�hh2��^�D.�~�E���I
'����]�dk~�t<�@����Vnn����o0oˬ/_�/6AQ�����JF�Sl-:?�,�v~n�����3;|�|�n���� $T�K:�2FI�u<]����Qu[�*�	:^�U��綾\��r��(PB����XTM?��7��Ɍ�t�!&����]f�@"Ƙ������뛕��0*g �# "p��.'i�D���!\��{^��h�b�L�����o�L��0RD�We�S!�vb�Y|��7��<� L�/X�Q!;[�&���)�����
���A�5\�#z���kW��3���Ћ�p��nB�z��!��ʪ�����B�a�X4{
���Y��Δ}Q�.6��ar�=�5��<ed	��F�d{�����������?U0KήËXhܣ㘧�M�J�}�>m�qO7{gZoM��t����\|]��̽�7�ӭ�ߦͰ��vVg�SU1��g�(���L̓����Y-�$�	�R��W�q2����GǼR)��'�)1��uv�M��0P�Ǘ�i�9O˫h�^��һ�<�l2��:�~Y`�#�����{�!���'���	=�vc��bDCe�~ ���_��g,����(Ag/��Db��������e'ЊIh�'�蠵�1�mćZ&�i~U۱��z�����a@�#�4��2~�|��gc־���U�cf�H�����n�� G+�X���($H�)�m١�[�Q���'K[�"���Q���qK;��/;��1�j��N�%�`��!̷�K��.X*�a��>V��`TiK��[�TK�x�l��q!��k��AidE1&#��>YPI�%ƶ�4-{�~<���H�Y�`��.�D*%8>W��I�����J{��Nho�MQ>x�鰶q�#��ѫ�H���]Kk��h�A����EL����p��&��%�j�|�3T�3�t�i�09�Z�O���O��`?8�+���z��-�0�j;�7�96��@ud�+sTߺ#O� ����������5�z��R ���;���Pj�����i%Q�ex�țh��C���J0OhN��K�ú�U�;�<�%v�����We�3��wV3w'��&��u��R�O��칛�$�C~�I�@]����
���ma��U=hRIٛ@�9DX H�/�J�e���v`��+4����~`;�+,������pJHLL_ZU�<��(z�	�>����f��1�[\~��\  �q �7��n��E�*����"2�F�Qi�.B1�~��A7�Yye����n��_��4�<(qkfεv��/F��c�{:��e��r����ʻ)�P*�#Y�J#�4��d`"�0����F�(��t�f���7�����`%��<"�4��D��:Z$��s�2���g����>C����>��M�),<W�Z!�[�`���aq
wvLtl�ꬮ�#;6�$���d�0�+�o����7�H����A�qi˯��L��p�~�k���j���ړ*{�Z,�<L~}[���)�T���W��zc^���r�>�">�x~9 6��IN�C��"y�k��F^"��_}3�qI�۱�o6N���4���7w���vjUt3����_� cV;�a6�8���2�F�?q�tȂ�!�g�
l���?ί�@��@L���5Tٚ
�xƺG����)�Iz���ܔ}��lfC񚹯h�n;��Z^�e� �J�)u�	ݕ�&�lV��X�^cRe��@t��0�`�f(������T	{"���a��w��J۶�I(�D�ۊ�.�:�ә6�˼jj���?7��K���Eu
��;l�j�cM�f�9.$(�W""���U�ly`t�F��QN����^�P��m�h�������hB�$�෵�<=hL?(m~�0UMrG������/��e-i}���X_G��,���c߉ 'y��M�u݌c��'q�̖�_x�h�o�Y�w8�FXV�&�;�5��b$���M'
eUJA	)����ݜ<�{'R��NB��{� Cg�eG�X�>�,U��Lt;�j�w���ᝐ�Y+{��ꫯ����u�
Y�@����ޟ�]�8��@�Q�<��-6ߗ�I������^�L���ꨶ����f<GX��Y�Tq�3b'�1Xx���L'�$`g^�&,����l8�W�ᶊ;�ʞF��*��������3{o�K'�I�5���*�U�����s�%y	���v��64�b�8l�A�
�z2𴧢|'����w���E/�d�$c���Ԥ��R�������l��	VSs]l�\����
���l�X�s��YDW�`=a8�?�vDBq!8fZ�@�=�K�y(���B̧�-]P�Q(����9 5�$��� e��O�����l������%Vx�7Kj��#Jt���'��Պ��X5 ���+օM�i��&��C�B�� Z��ᛒ�~'#�E�����'�=7�v� � �.�ӺBf6?aL��'pխ��Me~X5F?��Q�c��W�	:?�Ⴝ'+�si�X𴙖���h����&Mٵ~��G7���~�2���<��,�����v�,(�=�"���(e�g
d�'מ@��v~	��^�U��T{�J��O���| :�]���8 ܍e)�:īo^��g/�]u����&���(��=L�?|ѶL<�|�Ӫ��R�����H�[��M,�Hi�7��W"�1Ѻ�� �D��F��c웑��c��Ըq*��}N���}뻤G|�B�Ӳe{�7��V�o����^�%�M^�������	�Qs�FÍ�=�7���j�I�7r��r���a*��[��#**^���6�F��Zcoi�*cZX���R]d�!��k����{���Ե9��<�/Wqx�!�EY��i���!EF�D�, A�3�q��A���e�Ʌ������x�o�E���T�0e;q� `���ô��°g�Wn���rJ���c��m]|=���4�0��oeo\�L�ŃdNL!�ѡ���7����KyP5!{�y�;@/׾�=�U�ۯ���]�k�L�E�[��3G���ѶmŶ�s,�� wU5F�	��gw��7�Ɯ�O���=dnW��mr+5G��k�ʚ�������#7����� ���.����������[�@��Zd��ѷ:\�m�<�h�;Ů���o1I�PD�����[���uꈨ��^C��t�kBD�~�e�a�\eG2��>^ԅuy%O�e��#��;��wXw���@#1�q�+ �>5^�Z4:6v����V��}_Y�}&"���a�J�����lvK�W%�*� ��O��&8m�g38��X��%��k3jd�F��fj�����S	�t%�S��k�nbG���&�%�LhD�o:3�o���Zl�UO\��j~���� j"��]�琪�;7%��b����[D9n������S5�Y^^z���1<�U��am���gS9Ґ�^�Fn֛�pg���>�I�̙~A�K�a�T��裞'Q�P�NJ��S��)��,�Bs�M0`��CS�&(����+:�K=�nj:���N��`pTR�=*�&Ǐ�ȴw(Sf�:�0D1�z���8��?p��p�6�����G]���>��m�6a�U6m��&����X��=�vk��e��Tçh�ޯ٨���FmKȻ��#�oc���B����P�8����#j�һ@�@�Y(�������D�V�� ��1��.J�[�_9�ݟ{��=�!�=�B�#!_��a ��Sg1*��6�8~�z�L�&Ζ�(�����v�ޢ�A�5��w�����1�eƍ�K���,��q�x�>	It�0.;�G�%r��;�(*���ͪ�Gwn�,~q�ŋ1�l^�}��+a���S�z�q�VԿ�Იb���4���W8�6�Y|��>�����GQ)��K���P7�"�*��U�b�R�~V~��ᨇ�V�k�H�B�ų�M�$X9��s�/YT��4Q�}������E������Z�^K
�t'gE_s�X�˩e#4����H����;c%c�E�ۜ���ԅ�(yd������m1�܍�VB�,a���&}.�o��_n�l/�PU@}���k���B{)���[�+6��2��"9a���&�xb����ˏ���ת�z���5w��U����i��zv�u�<���4T����6�,� +��]�{^�`� lŲ{�'��nmj���L�ĠM��EU`<�s�5z��%wW�SQ/`��p��s��w��;y0�ۗ���B�A��"^W[����P
�z??W�#�2�H�����Kt�U:�����(���ĵ ����J�pr� 'fnz ����o�ЎaL����>Bc%#��M�T4V�6�\����=��2�K��64�L����?���J`�F���E ��aM^�����3��P��4_�2�Cmf�"�x�a\ܜ5��	ұˍ�S�Y�XVde�]}��@>����b�@�����1�Y�T#��^���E���sh��ZNhWN��4���C���9���(z�����6ܺ->�1�����K�~�`�!C�FMu�pe�WA��a��0{Y���Z�=���υ�,K�GZT!z�#�9b�*�L���iݞ��ҋ�7�ݲ���T�B=�2�������`��-�:���+2��gF�]�O4��4�G�9��_�&R����hKu�R�V@�z=-lhz����_��7�+�OJ���w�Lm��5�8�ؗ�])Z�m�� �av�(V��~��@�&m�I���[���1=k�Gʮ�u ���t�gh�a��8�k�� ���k�|��H߻����=5�Y�y�h�<�B�� 0�� 3v�E��$����&w�ju"2N��+�%�˷�\R�hu�$��59��[ީ�0�C�k��d8YV�Х�+�V�@󼙙��c-��sܨ���Ɖ���J���)�d8�2�x��9�d����8�'˪�Ҿ����������0�Qަ&�����=adѠ7���;�Jgt��f��rf״�y��ְ+�e�9���i�h��x���c�ͽY�D�@P����K��J"~-r]L�!H�r���ꢩ�vX~�ȹ0z�]	��dW��d���y��]�޻�*��+"<P��J�CKy;��Rf�`vi��l�<ݷ3R���k�cʢ��5����[T��9Ļ���/�4�����T�4�0�m����
vVǷl�2m�߼�;4��^};H���%���\�N�����!���Y-ĕ��r"�M� ��O���yEl�~X����`�L�|0�wa��z�ߪ�d=\�2�V�7qz�*��>��3������kyD$�&�K��ɑ�y4%§N�$zR&�o0���XCAbә�U�#��7?9�M��������w��s0������ut�\��na���?T<�)^�ߢ)Z��Ԋ=&}��o��	D��g��3����]p����:��Ө�D�¬k����c+{(���|7��&!��:��TS)2g�#P���.��l)�nD���gۖ�?�Qs�%T����&�*�5	ک������@-i�j)��;��'�Op|����� 7�K!����J碇Z)o�����J�ޣ7����$\��}>ళpR}(����9?���(_�@�	�vrY4�^3�����߮�cfY�E��q]D�AO�e3j�<�P��`%�g��m�¥�]Q2IY)�׸��8���y����O�H�8���C�j`�!�W��Sj^�ƌ�s�>ƭ�J��-�]2�C� M8�$�,�B$.���+X��1����O�S��de N���_��	��О�"@����o.�숒���:�����2~��TB�AD�k�O������J��8w����U����-x%mP�ť��U�n�'���՞�iͯ�b�d�Q��	�[�+P���=A���V'�<5�H�i�>��1�x���,��t��k&&#.�D2�ϬLb_��4�	��6�o�RR'-�١����h����K��;0��:�Ν����DK�����'�O�4/��B��9Q�͵vn���6���[	�!OK:�Oט��Q�[\] ��͕Rl��HB&��o#:��1l�y�nv�t8��W4���qHP���1��	�����qiQ7��� L ��>���������v�+v�h�#c�HY��ޏ���p�3k��bn�4�d�6^��{xh*NC���f��h%-�+���gJӅQC�m����⏢M�*�%gt���E�~�`J�2�
�F]����%���/Y�4i��<���FA�:Ʋ�%_o�"�Z�
�4�E��c`s�7�FK�Z�Ǡ^s&��5rtj���L�n�6��:n�:�_�};+�Y���e�Ux�N]�u���r3�ƙN�W=k �_��_a�0LH7(0��ԑsd�g�?�`���yKƶ]Dx6� �D����-~��0&�����P �K�P�<��R���%c-qπk� 8b��ڹ7��G=Kn܋�s��a�2�t�j)D׾0Tc�^C`tO"�0�S̳x
��9���D.[f�.��`X�psX(���9~�,�z9鋊�w�y�(��d|pmU4��w}��\8�<�hE�-CS֦�|����\4�v[�z`M�
ϔ��'=�JZ��s1��2a$����m�k{���]��g�
��\�{E�������$�</�Kp�pvҬ_�U�u�^%�
��JO,�p��}Fo���$�����ޅl1��H{�#z�C����r��=i���?�=3U�6���r��"�&W��J2�5D���Y<34X_�8�o$6	)����rBuC�{�/3�f- �~�LUTw�{�@��U�|�49�)��|������:FW��5��0Z���d\	�D%;�'�ԓ���Y�'߲��r8��{��^�#�,��<�ۣ�B|1�/N`_�7�,9۟�0�+�?#*�&�o�t���|}��_��_�(p�s(I��VP�艑T��z~:�S�}s�s����y�,�T۲���h٢��L�+���|SD�2��r-�*���.�F䍑���S��b���':�Dp"����o�2EL-�s������u�D�N�gh�lɩ����xR�;��s��;���ٱ�u;����O:����Ս|�wH�/�bg�$�����aǓ�ȵ�MD�M]"�k���j��O	��G8��+��)	ޒp*�Pz��W$�¿܎5Z���V�*�|�) ��-S�2�{�����vqlLߑ�2��*ἔ��������z��Z��*������"�2BW��ԉ.Ws@�Z�X���i�A��H?�US`�h��C��HP&-��r)�ק]��9�w�y(��ȣ�uH���-�F��K}��uI�_l1�%��!�T��H�U�Ry���D(�~�t�V�c�b�(<M�k_��5L�Ү�&E�琎wx,�o��>�9��8�<�o�V@�Q�h�����jq�d��B�yBH��M0j�
!��N��MӉ�`7]u%����R_�]��~�^b�P��r��&FJi�o�a��춠��	��ez�D�^�r�0��o���t��L���&ZR��2�)3����QQA���F�	��n��_8�3��ti�Ɵ�L�����u껠2K"x�7z�t�C�QS�G�X��o��dѹ4P2�K�e���!w~��'�5�dg��R���&�LΒ��%����+��JV^97����?�w��0���
E8�0������i�wĊk���3�x����و�p�ȾV�\0��y{�]pA�\��:���_��!�&æF=����i�l�0H�Kd��hy
ht��ԙ1�~��?ۣ�$��l}���[��,w}�EWB4`����w41p�Z	�ǧJ,��K��嬟�f�ACAZ%t���X_�-��a�SQ�������JqIe��)��-�LLi��QiF�֦��fF�7irh�(���)�d~1-Khڿ�C�W�I#��r�1i�LoX����E�!:Eau�i��Gu��͜���'KG��	)�=����F�����\�
QЌE�"��$2����͙��"ilh��W�_[b�[�9i�/��L����p�4X
���pt��Z�n�s�f@��#�]�6�u)E��[�t+��JJB�ѵ�t�sLxrܵ�UPA�&+�8nk/��������bBL�_C��y؉��m�{�0��K��� q긗Ҕ�!�Ɗ��C�;n[��O_��� f]B6:�}��A���h�34���I�@N�F|��Ьu�.�ɥ��2z��B����6lfX�G嚜RU�w!Rq��͸W7�eƮ2�&j�4����n;Wa��Z��֖��+�x}3r���fa,C�v���:��O�B:���XΏ����&`Z'd
T_L�SЇZzŁ����v�I]�{�� ,G���^@�W�R9��AS(�m�j(�΋�8�b$��7���p�w�Y>�Ɗ��_�����gO����뿨�N�j���.)�=|T��U�Ȁ�9�O�0�+]J�y�a^�e�SI<q�NP��Ra*&j��&��\g�qM�91��vN�1�¸���I��-e�o2L>�N?�E��R"j��E����q¶�?�	>�Ȟ�S@��Į��2�<��%6� !���C(�g&߼��+^ma4�eƼu��Hr-�6"���5���\�u}�{%[���,EK������y\2�C���NlA]���=[�h�{�3��<)��4q#k��t87�.��ȵ�I:�7�����eU��C |(L�@) i5!�è����xh�� yf�Ô�`���ϱ�Ѻ^������@OB[�q`E����B�}qe���:y�_��������wX�D�)y�u\�m�XЅ�}����9X��y�:Ÿ- �jW=���[݅�姀�~��R�!\�o��0:	 �Kn��J�[��{���~�~�^�d'�Є�a�+ņO ph����ɰ�e�jO�D�Z91�x����n[Y�iʠ�~��I,󵈾>���D���2�{�Ĭ��c��b1p���_��l]�L ׸ncAp�Yz��x�_���D�x-'T`��ƻ�2��O����������*�kXmp��[7��5�ݐ�@���/���,v'_Qy��^
���<c��h��q)�~P�N�Eo2P�:2��h����y��pK�j;!L�u����tUL~}�:�(�q`�4��u������vHL�+H�W�t�|��
N���ܡ��࠶���M?�1yd���{F[��=�u#�d*
d���HsE�㞣�*P��:��#�H,V��t'q�4���!�&����Ϯ��H�|��.��1>`�|J�S��t�6H=��U�9��C������g%�v���'��٪u�kl] �~ė���#�vqN�	��C�\�ݽcvxX�L�'.#�:�1�}+v�?��WQ8�"<������Eʲ��H��r�6! 5�(��g��`ciR�"�Gpl�o@��1+~����b�<����j�x?<��0>[|mJ�O��(��Ϋg��1T�ɿ:�0�����ȫ[$so�`5=E��4�&4�� I�y�#&]��K�.?��t��V%T��X({�R�����ף��Ă�t��	'a��9�2������!l���c ��+N��KM�A1䄷��g���[ v�Yc���	���1p�'_��y:���u�FΠ��G�X������4��J��q�FU���9�����Y�.Й�����}��e���d0�e�\�1�cϊ5�Hd6)C����U�0P��/eoy���0i��2u�Z����n��b,y߼�A��Q-��bj}hC�YR��_�)4+��?��.>��cݲt�j�%��^a>࠵�%`��ö����`^G:ۜ-��a�nPuf���:�R��l�;W�+l����=�j���2~��tI67Ð*A�Ꮙ�_�V/���w����U�Ů��>D#˵�R$?����K�Z����S���1����R~I!L�P)�c��C�b\�_��TX>�H�}ֈ2v����d��FF��su)C �|�>�i
��>�+~I{�=<t�<ڂ�!v���a0&^>���Ч3�D�,�G�9����P��lg�s���+�71		�g��$-�O}�p�L����)����	đ�6ԟBb�(�c�����?>�0�	�	,��-�	|3)^J7�I�)k��-�s5WOk�A�¡U;m`�4�S9������т|N��ϕ����g$���.+�V�}�I�L�w�?\Rt�._W�%�s�G�.�;P�\zl�n����15�R��.���+~�qOY_�*�l ��������_D7�t��b��K�	�ٛ�i�jL��ҙ�aj�AP:�
��£e�3�@?*>U��ty��{���O��m"���`S����5�yb�ZI\4l, ����zQݢ�e��:�?!ך�t;��O� sE~�@��[�q1��rr0�1m���(���X|�ox���
�7
͉��fNbs���w�D��ЃL@»�1���K����r��	Ķ��m==<���Y@�(?7(�[7��$����gh��S`�i�!T�7t���~�21�����;�`]�É��Q��M�9�̔��}�.���fJs���ɹ��w�Y��ژcF��h@M.�I�FL�}����#>�%�쒁�K%/��v��݌M�@zQ���
k=��.��g�U�߹۝
�@�?�����;��E7��s�Q�I���!s�8��&�B�4�{lY�e��c���ȹ�;��|�%��σy�r�'�u6���Pz���3U��jp1$�i�|�o�?��8�#$��/0Z�tv}yuLW��I&�>�.D����2N�T]��VI���<M��.�89ޞ��g�g~J��� ����}!�nD�R���KQ
M �е���ɺ� (�V(�6�_L�3�u�ك�\�{��e���D��16���8y8��R?b��������O"QpS�v|�<�@�臃C�u��,+���INq�>{��9�v�#�͘��OڍT'V��3��&�+o��j׫;�+��CKe����*:�a&���47� .��:�,t��xL�E�$���Հ���"���7�;֚��w�l�1���
�Tr�g�m�����n�3�e���2_����J#	�jkt|X�)�!l��L�8���:���沮ݓ��#LlN��y���k�믄3Ϣg_}!�Vޜ�����g�6�p���7�n=w�F�Ƕ�ʚ}v��}��dY�u�Ϧ�%���CAA���ʄ�Q�y�y�i�\5�<��N��-Y,�7I��7J�:?5:�U��$�	�P�3�5�v"^҆��H 3BS{r��Z��'�يIh��Fh�|��Q�;�~u�NE)�[
��QU�er�}���@9��ƛ���Ѡ4q�����	3���M*	���LQg�ⲿ�q��4��d=���������\�3�gÎ��/m�q�\_������mߵ��*��Mፅ� qpO����Q�fMv֨��/�8!@j_8���uOhe���ϊ�۳�i�J��)�����[�ڲ,��D��T|vYu�+�6j����G���(y3��\���X�3w��?�u�5�u��UzKZ�E�|�'���#V����!�;��Swv-����hs��b�x�f(@N��d�L�F����Z��W��-��:����
��K��:�_}��\��@k�i�,hV\A�pf�A֣I�6GJ{�����AĹ� �{�ջ��+j��]	�������O)��ɟP�GQbFZ�{a�
w9�v�vH)2�Ue*Ft"1��1G��辫E���� ��u��duSNg4��˰�k_˂���~eZ��9�axq-�G�X@��dƾ�6(|���:�L��P�t��)P�)
/Z+��Z����rS]J��m#`�z�E�pz	�c ���Y��ʥ�L)6ON�{�-
"����fx����~��X���)�!��)��K���А&t��;�m)J�w�rB�5{�8e�4�w�O1U/�*^{�EH�Vm��Ê��u����&��9AkͶwL�κ���ߵ�PS8��S	$!�LK�Xe1�ܸ��#n$�[��x�Ore0�J�ꎖӟ��BK��֢��f�"3�i�|Ug���N4�����>�fɼԇ����7mJ���S��$���ӗ����p��8�Y�xV�IWXW���y�>��sO�ݫ��'��ⷷ�r�P6u��hu�)�d Z$�v��q�1��j��p�]c��莽�˽�i���X�?X=t�N�i� �$���R��ߧ�Ln��/j�vAB��U H�d�/F^&������n�=�Xj����Mj�/�(���K��R)/��]Y	�	�s���L�^9=��ύ�_�/z�i�9�	i��g#�:8m�@1FE���>E={��]Z���oU�x��R~�^)7-u��5�L�zXz�sL���"&�=�{��d���0 ]	s��ፕ��ǫ��V�Li����Q����M�x�0gq۞�0�c�e�E��(�C�7��><�vr?;Q�$�'9���T#�:>^����t�.]&G.����.n��00/�%�4��E/��H��[�Sb`1���]iX�ֻFO*����aG��;�?�u&h#� 9�ݶR�k���C2�Or��M�tS.�HH�~����>$
���z���O-����YZ*ߢz?��8�%�"��R|�:�Ό9��K�+^��;�qJG	ޭ��/``>P�@Z�`���l�7Gw�Fϼ�6�܅;���آ�c��I�:x�JmR��+�[�-HT�oo[��R�2���)>�8Z�V3t0W{Ϣ���e9���`NTk "��Y^�5
�{Е�S�i-"�#+2�moKx��R��u�x�w؛-$;���b�B��r�Q�3������^۝����,��)�i���9኶ �y����|���YU���ymrM���1X�F�n��J�B=H�W�GV4������݌9�E��?بC��K3��Y���1I6a�`H��Ypħ��'���7���8��_|O����U[ڙa��6����ƥU<���JEw��[\ʚ.�a�c�b��=lp���sZ��0���l�� EC���-��t���
~͚��җ>Ћ�\�2J�%1�aX#����8�s*�n2�m;�	y��>�m�k:�3u��枺��BTƘ�"l�O���3�ޖb�}�v^Kb(�Me��>喝\��h\�s:�LZR�6S6nK���[����v~7SS"��A1�VEG{���Z�a� 8�H���3����	g7m)�s��7��`�:��p�lQ��e�$2փ�@U���O��`s�K���(�
�<�����~>�L�>CW��KA�*���
�����x�?��+N� mEy����oteH����'b+p�b��[��|��V�r��՞���r��!O���;��y�S�[~�Ī��<K�>B��	�B7�\: @���CZJ�d��ڝ�#��p=�V�����!6�,/��#F�Y�4�@?���$�薞�Y��p��е0W� ��n���2PX�s�8�0׍�kI���0�(9�dG���2|o4�I�$h�0�1��Ð� ��#��%T 2s1ޚ@�z����/���(U[D��p-��]*q��?j7��M� w�40{�ok�͋8����$�ɊEݔz�p� �fj�N@����"��"��$M��)vJ��Y��vh7���������eafz�?a	E�Q:���m:�I6̶p �u�bv���+�S!F:�t�L��Ʃ�x����$�<�e8�,?�È���chO�m�yJ��P;zl��I2D!i�������=j%$v�2���uJ�g�d���S~P��R�����f'�ukc�bt����������	�ֆW#�aY���wt���ONX�(u�1��� 5�@�H&�L�ZN|8���r�k�����(n��t�5�a�}��p]��9;�� �&��|O�0<9�֡�:d���q���D�t���!�-p�\��G��Z4P��}4/Y�}�u�T2�ߌ
�3m<���Wk+r�mr��Nn��O'�n����I@6�]�gBG�F��_��y@��@��;�9��jD*�wX5Cc8�$�c>��d�e �3�T�\�!⣿Ҏ� 9���4��FB��*�������_�u>���ǬX��ӝ,x���U:��X�Ij*�iڅ��!�'�GU������2{]9}������c�XJ
V-���ꔬSO�\�������~-�+Q�.쨿�����H��A��O��5���aQ��'7��AX�5�EJ�ޗ�I�����ֺ5���Q�2�X4rOl�p	3m�[�밒��E��d\�ď�mѯ���w@����@�O��0_�{�;��ĺ]��,P6�Q(�IF��˛��"�a<zC��\F���� ��>4�"���6���-�deX�&�7ݡԳ��o�%��Lq]=C`�l��E��
�;�H�6jB)�C��0N�JG3/ƽ3����XW�k���k5��C��A��v��':n�^���9"S�%2�s���M�fX����.�T>�2��q�Gg�o����ʓ�6&W�y0nWS�Z�.T�i�#k-�Ng*T}�H]��	��������X���>B�'��F�:�0�	a�S>�*��6?)�[F4Q��2��c%HkR,�.��Z���O��W����tSe}ʣ�nޞ	 ����_�H�ٯ�6�P��c$u/��	͛�r>��a�B�[ʏc0W�<c�~C(n5F��B�5�g�L�uҊԄ!�`�(�&�X��F���O�N��?z���<@�﷎����&9g��A��p�9yGO��/q����i���/#��ŕ���G�z<?Ka<����k2�}��}����꣒tc�-����[���IuMrg$�/��L_O6��4|i�}���u�j��2�i��y��A�ǅqW��\ޮ�7l�}`��d>�����~b'ndlWyZD9�b=��2_M��; ����j#�\:�7W/��3�ܶ:�F�pɤ��:���VJ
��� y�8�ƿĘF�%9Û��M[����DI0׍�?i����}(�QD�/	�x�XMh�l[�W���3�	ё+�P���K�ָ��a�q��>%�x��,�+�Q���L�M��Ρ���㹛�����/�^�W�*o+'�7���:g؄�r4��LD~�9�j�(�?j�	�$���(e�d���U��-`��dߤ��6qS��K �5!�sc�3�n�kAp��ckX�12 +�*�_�����Hn�	�lT	�*�N|�
s�4?��7m��{Y�|D���I�m���3�L�h�-�����!���R:�ހ�C���Zd1�Ge�gK[����? ���z���恵�-4�ّ��6�9Դ�6��/�
0���J9UU�Y?���>��ŉ�j�%��Ȑ�����6R���V�P���qc���(�I�ޘkA��7A$��]���c��5�w��ۗ]�	�E�(��;�ur���b�����Y����Pb�	���B�"sP2f�"IX���6/�vl`>��V~���}t�$�Mײ�(W��F�~��y��!�h�ڒ.#�PUw��>ϰ[�!��My��>Oh�?�� ���xT�N� 10G�:w\��Є��i�am������ϊi4���i�ci�$��e�5"��.7K�@��T�`�E������ܸ]&��@�fJ_ȔF؈#o9�ga���A�T=p�\�^�M��[]}�h��]���k
���+����l�����aɝxj�J�Ө��Q\H�e�0���Ջ<x�$�^c�	i!5��ѩ�.M̸@fd_�s`Pj\��m[t��0b��G9��/�X���wO껡/Y(��j��C
9��������H.�Fv�D%����J
0L���fR��SSb#yeLo�D��g5�4d����}wV��/�ʂr��̽���S�V�C�w�j�f8��cJ;�s����x��d�`��I_��Ʀ[>4W��R!�"!�S���'�NCB#��R��e8@a�`�d�3�t=¶K��l&S��;��eQ�w��[ٴ�(��z5S^���29	W�Y`�Y�#fQY�!�lY��&U�w�LXe�M�\|�4�oBO�=��Ś�`�p0���3��BF���Ytưt�G"���GoF��iӻ�W�:<��m���ca$q0�O� ��JI��3��� bYj�
4z�B<�>���a�{�l8�9h��ۂcC�5�-��(Y3 �o˾Mwx���P�I��M�?CXv������z&�b'�-�멺�$��7��_#aA��q���F5{����0�k����v羦�4K5�8_w&0& �	-��i�䑴�¯��w44o`������oP�3�i�,z���q�B���п:��$_+X'>gP�Q���-�h�?e��n�8����.H��w�{G�h��j_'�!���DW����']���Ꟙ��>�9�����4��ǋ�7���� �-��]b1�T/�����|s�|�r�ā��tH�3{�J�/��o��ms�z�dyU��fݼRp 6��o��A��X���`��<tǔa圢C��lފ�� � d�C�(ԹX�]�WAl��E-ҳ�zI�N��  �|`3C��ȆU4˦�&�D ��>4c���gP
����3Q��d�r��WW*k�n`����3:����ӧ��pY�/�!�~>�vm����kB���~D�"�i���+ÝG]�������z���A�l������
���?��~I٭lp�\V�C�=6�i����߃lX�����re��Y����p9ڐ`�^�苡%���%�4�:��Q%���e���O�	8�+��(�+�u;ɵ]j����,n;;b߬��S0N9\�+*����^pP�+�b�3Ɇ��;�ə ,�ܸ����)kw��,��d�MK�*�Gnh#���l;�"GK�%����a�2�\�JR�}��oVն�q����L�Ǽ�!M�A�nִc�h5oJ
��y�ғ{crճ��PН�u�&��NWm�� ~��eI�|}������@Rp�u���Y0'�^N��ި]�V�*���<�PdT5z����Eg��hɈ<�%,:�8��G�u�G��+�{QE����E��:?ڵ�o:@��wZ2?3b㌒�0&V5�,�E��0�̦����f�a�^i�mF��]��a���JF`�(G�2��O��8J�����/�N�,H30�C�r=�Ո�Q���5o�?�{���ca��5�5��!�)�l]�4��y����YAa�5XS^�}>ڵz4\����H�:��S�5�1\�ƸC�~]n	s����x��W��F`w6/6jF���ү�B-f��b��Ww��瓴���G0�=&eɂ��J�hSJ�8����T&T�l�!t?]dV���?4>��I�� �pie��g�/*n�Ԫ�b㐳���P���C��/�2g�W��sF�dm��IV���A�p]�y ����uR�"��w �#<5s�J���.N݉;�KF��E��
�F���J]�� ���l�? �e���Et�(�>��6���g�o����m���N4W�٘�Qm[Z2�5X�N'�D-��ˉm=������	9��Z���É���Z�z�)n�D��J$�	� )��mQ@��"VO?��*�D憾�bt�4!�Q0}�p7e5/+tzj>D ��i��pP/�!E���	�/.�M�Q�cX�4����Y�4z�6�)H��p-ef"v�r;go�^��K<�� �0)˅o2�V��,;��v���2��P���@�Q$JZ���Ȱ�zi�&�X�soe������O�����ظ���
~_���.[-:��-g�T�cwV��7T|M{�iQ�F�YȈׄ�\���UMǠkc7L�
�������^56?N&b��"��Q{t(G�si��~�"���7*("�� U�,�W�L�)H?^7��'-���m�^ �-7���-#{�}Z�B�ѣ�I�o�[�D���8'��ܭ�ɩ]RS�(��1��an����8h����˓��A�D����V���S_\G��@�����@���@�n ��9��mmʈ|\���a!cV��"F���0G]^�قإ����ٸ��LT�`���!g�LA*1ߨ�۞5wI�m0o��#"�>WbS��HIgL�
��p:$��,�2	={B��h�H�Ͻ���G��kvk�k���i��ٖeϨ�|G�-=�z�]��׻��/�5%�(Di��2+���5�� G�Sp�#dnIr�2k#l�͜�zp���Sǽq)�S��QtА]WQ~��B�s�k����YsF"�m|�Z�{�B�L��^�,�]-e�6q1
�����6���e��nnh#p!�C*���8���\���i]���-(i�ص�����r /C�N�>p����5���ꁒ��ֽՅ�5_���5���|L)U��虚�}����b�:W=5A���l�oIQ;�iF�>����%��|�Nc�܅�	Jj#��*@�4LIl�8�@����f?Rz��mJZ:�[-�x�Q�)�!-�(��(��t˦I�C^1�T7�� ���N]����*�v��8'^�Xv�|�:�����Ѷ��t� 0�+�_�g���L*5���?~)�=�kg�r�i$����j��V�ᨂ:���J�J��ɕf�VTۡ����k�O�1n�55�6�;�=tK�u̕�	���t$�^��5P�Q�|��Z�t��xrL���0͖��فM��ә�[&���cҨ��4q�R(�]�>,�o6����5&�@�0!���b8���a��L��ݷ�Ɨ�mw���&��,8'�(�2g��\s*���ig�Q�R���j���R[�u��C�l-�y��q��z��; �ݸN=W�<�����N�']���ћ��_�sǱÏ|��
J�q�%#�	�|Yڊ�7ͣ��x>f���qω^��f�s)#��)S/L!�4�[Q\w�\�
d�X�%`�-���� ��4\�I[Dڏ:���ܭ�)�;Oq��5h�x�ҊH���^$�LƤʪ�%�1.�.��?���V����x��[���H�>���ܞ�^:� ��¨7$ےAzn7,�E�i��3<�6iɌQ�_N�ő�����;V���É���)����_��:���z��ܐ�[0H0Te��76�q�lri� �y�^sn�+�?��'��j�W>kĀ��,��_y��8���e��Q� �wޞ����\�E�� ��b)I�&�j ,ӭ��7���aP@y@ZC����G=�t�HW������1�b�������� 
��d�qz�����\�$h��dOV���G�q��6he:0ы׌_�@%�B|-*u��jG�D!�E��q�h���)���[F��6�9���}�s�=��?����g��û�3ND��)W�
?�ܩ:���Z�i�4��r��)-�v4�V�ޡ�|�	"8̣Ŵ�"X�٢^�����e��[F�r�v�e幝��Ɋ�u2w#��f���ip�1�g����B��Zks9H��21���`�U�~�,�W�Ll��R~��)S]�Z��o�)f�4����&��'�UD-�"I���4zL���"OG��'w��8�5n��v��n�9BhC�ڥ�8l#�N޵JG�!&-���#j�����xRd�RI��p�;I�+�l�8��� ��31�xJX���c�'*Ů��Z8�[�k*Fa�������5:7=؇]�L`M�>�U�'�2�=W�\%�e��N.��÷>����A��@�Hu�t�w���6ӧ�*�s�j|Iہ����E��r �0M�<�/GS�5�|�攔�B|��n�V��a�ٝQ6��l>�{ྣG��"�=`�pV����>�{'���+):�b�'`�����
�!���φ�����w/
�q�>�Ǟ������
��To���瘩ݟ>�cn �^�A���:�o���ό��o $݉q��vk�������V�b� ��t	<�l�qe]~7/���j��'�\���jϮn���)��HN�8����*f��Ec��9Z�Ӑ�Nȟ��u5䝀d�r�8�|�D���S8Q�e��c������щ���}$��7�}�w��u��-VN�",�W�����Z�r����>wU�^\���݈&F�ǀ��P(��n �.4�+�֚ �%#�m�w(��Vs:0�E�.�����P?H]I��iZ&�y�O���1�^6�\G Y/V#�h�~����tnvf�pe°�Ј �@R�65����-�$c�c��^-�=�M�!�����v%[��yn�K�Y�:M��s`A���\a�W䰋�kq�$�L��=��1̛�-���BA{{�e	@owד!��!Z��0�����W�	 �%G�M��dMb�Sg	�%H��	�?&W!�����!gg)�{�Y��X�i�	�=8��Fkѧ�`�N�-��_}�E�e%e��{w0�Ũ�獌V�������3Cnd'h���߮bk�ue�����˭����nǟ��G~�..�z����_Dy]�T��d�![��@�;��l**���Y�j�sT}e_4bl/Um�Ԭ�j�(��Q7���D��[����x�utk1v���*ph�B�h�hD��P��%� :����Z}�Gɇa88-Z������sTuXj���몭&�T�4����~�IE�/�^���">���N��V�o�^ּ�^�O�WL:
�B���<�Ū/c V����I��m��.���� 
���|y�b�O��rL5@�!e�����+��A�cm�P6������	�����DR
ڢl�ǅ!�� 9EXR� �e�fK���!�[�1(��@�����$��D
^�d{���+k�����)|xTwmWG �K���{���^�Y됄��Ha��
n���&�sI���=�B��Us��������A��x��W�b����
Apn�(KyT#NMd$D:��@{��8������4$��Te̗��xe���4��MI	��^��A�а����5�ᶊ�1����Ch�Dj#KK�K���U��a����u:�P��|8b���8t�2����+T}b�����6�[��1��[1W��l�?�����a�a�,��>O(�w3�;vd����T#3�k��?��d�3�i("����K����!��IgW��C���7��U�k�ܨp`��O�YCGC�dGk�� ��{�(�2�����=�8�������])�ԃ*�.����cn^�'��YJ�*Űh��p��i���c)�)�D����_��eܐ Z(*�H��r��x\v�V���n9��Byg|F�-�;�oA�CM�Y�#^�xԪf � �s�m��'�P�L��'6
7@ >�j��&x���d�#���<����i�BJ�"GS���!;�"����V���ޡq����e-v���0��vQ>r���	��)l_Kz}l/&� ��ӾŊ��n�p;`�z�vo����żp������O-��a�~�e�g�Ċ+�y��l8�\����;chd�߈}�YrySj�Vr��r���,*�P�&�hT��F^e�p�,[S�t�A*��Ja�����_=�h��O�,D�0wS�%���ć]l�u�B������\G4O��B#��e���.��K�X��r��Q�>A,�O��m��,Z�*>.R���~�3zCm��N����V������Bt�5�%���.��hutIe/dk8��K�n�υ�CI�8+N�)�0�7���Њ�{J՟fMN�ea��c"����Ë������'�3֑1�(�T�\/R������e��P����SF�����$��Ѣ��'ڦ.:������X�Ow�?*�-/W�ۏ��0A�n�~:;:th�LL�?�4�`L@A7�<Q�!r'�"JݕV�<l6iªc�r��6�9�w>q�3JAiPF��q��A�b�{Sy��(�`�b��~5����",��(4¨�l�����=��Ws�O���B��#�>������i�G��i��>�:S	��!9'�H�<�o�s{��9��Ct���I�Żu�G�ƸRǖ��}�0	fp��<-k^۱�t�l��f��y��²�Ԑ+�m'#&O1h �]}^~�>�̬cQ6�gה�%��3���?{s��԰�`#���>ƃ ��k�T�v��S��%�@Gd�/qq��7�<]��b�];H.]�1*C�ʏ~�����g�G�|r��O��؁��wÕ{&�3HKN ���l������V�ҭ���AP�9�<m=�*�q�\e�&B��;g���E�jg�S��k�<٪�0�5�8[@Ż};O"���`��b���s`��n�]�gi��ӱȰг�X�7(�+��Bj?迃8��(�W�*�1|���1�G�qm?�R��`�c'��>(�!.��74&�'=8�3���j�&bY Nqt_5�Gf!���a��:�Td@���~��|CW�� �0=�<���o�E�:�͵�	K��|.ޯ8���Ai�p��g�[��#��a����E��o��u��o��)�/wb�g*]Tқ.�b��.�(�����MqR���A�/N��v��-�Aj�jUR�%����6�P�D:�^1T�~~ԟ��Z 3�@�5�x��o��ZP�s����?���M�~7��W=?e��"?�o9��0�lC��� ��K�nۀ���0��{q�Ύ�v^wPƟ��gx���<8�<7�Ns~�5��+ORs���y�l�'�{2����;����'��L%���o���0����٬��6�ǫ��cO��2�%R���}Nyu��/��
l{������i�!O72���{��)��챽Wc��9�A�$_�I�K��C���%�g�v��F��.}sr������{e+�Ϧ[�!����HN��e��-�w��r�ryt��Ww[�!	]T��n0�ts�>��ew)̤%��s���xH) \n�}UN#���$���� ��XuK,Ë�e�σ7|�0ĉ3>�)a��ZE��q��R����&<��ш^�d��|�|7R=יSs��խ�GǺ�4<2�nNE�G�
9���bY�:@�b���|W��Q��@��(��S{���7�H�qm���G	�:r*�mQ@�p��Y��_�П�
o�Λ��E�b����I�N��ϮO�{�mNNxB��o�@��%*Q,��g$����a �5}GH�	qM��AG�w�ᇮ��]dNQ C��*���j����;��EmɰM91Wx����$�.F�������:��\��o����y��-ot�o2'�AAfQ�G�T��xd�.�g�g�DK�n�����A�:07���9rHvE5�Ŕak������$: �s�h�z�4�K�4j]8X���9��#���<~�����q��;#KG�4l�a�ֺ�]G�I
�)C:��߳�@>���,�6�����$���I�������c2e�TN(�/��&�K[�ufqx:���a�7��$�\��=�ɛ�=Et��|m��\�L1W=��3�p���y)-�e|Β�h`|����)j�Vb���v���f��{$|��3-|o,�����a7�*g[<��" P>�\�N�Ê��+ԭ~`��u�}v)���%�⹌ⴛ���k�� �>���P�*�-��e^`
�@d�oG�X÷�i��]��Ѿ��t�\��T�.�b��&�do��-X�Lo��}&[̮��=� � ��4b2��$�q���@�Q?{l�q�V�z�>u��)|��=	��2�8�I^���X�����e@|�A�Z��6��
^�f�1T�z�����騪�>ܺC���'���3[��#�O�:�½_8q��z�g�G���EA��"���6aَ�l*rX��^" �5�D�.�\�H�̻&%"�S�AE�򫼑�T�Im�*�ubN`����pX�v�_ؠ��u�W��M�Bat���8	�z3���%1`�?a3�`�Y]�!,M�z_v�`Db,�	e^5m��ȬRt7�c�/�le����xeB��z�J���;�� ᕽq=m:�#>=����Z�{�w�i��H�A�v���:���V���ź<�p��};���	w=	����:
��R��V�� ٿZ�k����6��׿�J�F޹x���˧��3��_�9���" �Zq?�f��h�͔� ;����SNG$���[��8{5���N;jR����ȁ���eg��������pH�\������O�fރ�����I|q�ka�&�p�2��=y�j�^��bj#�B�㣈��1�Ʀ����Ȱ��t�P��t�k�|�&�c�u%���w��g���|-��V�Ϡ�+��,C��h��A�%�JR���P/�i�K2(�È?�{�4�1�j(���s?U�{MҨJy����� ��.)9��N4�P!�F�ίK�0���F�
s�(
+����#�j`l|cUtu�.id��/$�����~��0������-~F���?ʂ����Cdm�;��UG��'�1�<?8%)����W����\d��G)��Lc�t_���h���5i����m�}jG�<���*�>�����+6�S��4f����AE�i��x1��k�����@ަ��U�)m�ƞER�wfv��?�gL�W�{�,M��ف�;�{����@�`�}�4�����p�R �����;O��t
ז�M�^:��̊&��Vd���YY�ݛq�>y�W-:��ϔ�	�)�v��}�3P�{��zhf�;G"H��������6�<��5�d�߇AC3?�EUGß�-
py� A�.�G��P&q0�t:�5�g�c��[��#��k��}U���l�CЛP�8w��P��ڢY�짬f����E�0�4�Ϩ�yz�{�����j��
Ch�M����k��:O�@:�����F_H�|���U��ݴ� ]���(qث|��(�L`���J��;�\w�Ae	�����^��t�P��S�[�:D���ձg�Kh��9X�<	��%�c~��u�Z�pPg�IF>���{�����_��2w�*���&þ��3m~O��#���m����>���^»�?Oc�g��E��
-ڜ ����NZt!L���]ê����M�����5[%�|_���|)pL=2[��c�&�=�{���(�s(�o���-B8"������X�G,C����`�bs\T��
�'�y/?cY�,����yGH_J8w�\�ug�mA|�����Q��� �=Z���Y�gI���]9��K�O��g�<Dj�� �l�fzz���,���S,��$�-��<7���X�C�R���7d� �L1T�[��vcT��z�����H	c�>o����~�B��$9�M��:Yq-�H�������_�.ѡ��jZ $�|��zP�ƶ�"fݴ{d�\�0�~e�Dy`�тl%վ��*&�����;�$��"!Ckq�����fw䜉|̔"g6F'u���<r/����������@H��LK�dA�,nz��U�����m!�%���;sJ����q�#1�e��cE#MoD\}����]��Ie�'��H����g�Lϼ�K������>��ӵ�<Bg����Kr0�_d�M��A�_��M�6��f�G��:�EY�8%7���<eS�aQ�42q53�t27���1▣~��1�T�a��N6�S[����6�^�&��h��m���X�䅗ra'3!s�N����mE�&}�r7�)~�?쩱�&!�c=�Tx��a���q�`������tR��kw}�::,����٬�a��G��Ȑ������J̍���?�[�{�)�hr#Kq&�����&�<n��v�Ҟ�"?vtP�.�R�?�L����s�*�V���g�
r\WҪ�
�/�[�* ΍��GװIP��+�\Ǖv��3��/JG��l:��	>v��@�R��9�.�tZIL��:
Sc�^`!j�𸶑�0W�Ȏ��u�4E��,�Xd�|:�gu����5b.�Gk�w]�T�4҄��\g0hg9��앛y���"����N�'��fI�����0@c�ά��0<[w�{��k��Q8�h�-�J>*�؄l�¶'�" �2p׎�%SW�ک�=�� ;���H�z����6�S$m�D70�e	-:�!�T*l��r�<�\�$����TI�*9D�=����� ��ʾ�o���/�����#Ƿ�q��8f}+�[<����D�2���y?�!���!&�fb��mKl❅��Iv��W�,�rK��6*��e���;��E���^���ߠ.��%,�?mo���)�D֡1� Ҵ�N�Z7H5�~Cj?&F��T�,�RRdM�/��\/�4�������O3���)�T&4���/��:KT�尨��>eQ^Z}�����Pms/p���};�H�uګG�gCkz�؀��FOTRn9�뿬(��u��n���iC&�bc�	��#4Fe��|��n`Ņ/�tI�L*��j��/}��!���E'K����Z8{"N�H������	W� gp�e�)X�;`�b���D�x9���B�t�'�dsw��7�v�iYܐ���Wzo��u/�_��e Y�AԎ�Y�-�8;ҁ����ʴ�$����_�k��zYݿ�.������α�5���q�!���f�$����q��X���FS+S��d��Њ�Q�a��� Z��.���]�;HF���������*x�lx�`��6�D�HJ��vX��!��톺LNH�ëz�ς���
��.�^������ޮ�+s'�.���):���3����?��7�����Hz�0���q��;y~��s�24�1_��B;s�Y�[K(�Z��֡cIf(�3���C铁[����C��� ��Ag��z4R��/�WSC�z�t��7�"Roh[K�U;)�0"sW�Jn����q|�ݾ0Z���X�:s7�&1�]�4l�"_���E�(y��זĽ�xJ>����y�t���OI9�>?H�`Z��ut%|�*V��~�/�gD9�~5se�5*�����vv�)*f�j@?�&���u��=�t��x>�Q`[�D*���I-6y������xw�O�A�����j�tfȤ�o���U5�}���<�ĶE��a$��<�?�ǹ�gG!�%�)EE5�3c|/o���+b�1�Y���ѹD�NOa��b���evIw��R�T%�Q��#�	��yפ|�͓0
N�|�C����x�Q�~�����YL�x�*>��KV�DHwyp\���\�D�g�N
�)E�ƃ@����Hi-���y��Hq�2��(���=�x�j�SFY����F��Sc��Y;��k6�L��� ���|MJ�I��0���U��4�����E'�O>���1gT�׶^dGA<��\I��8�\������69�*?��`����p�g�^V�j��9Y�bsMS�.kǢ߭q�:*P>����<P�=R�4���x�ǈx�S�F`���E[o�a��_qX�Fلʔ�ewa��%j�_9/���.�~cF��U8F�=��^����� �U~>诚A�2^�!)0Z�<xBǍ�8��b���p�5�?��0�+j���y9�n?��R*9\7J[T[��
W,-Rz&iH�NUO�)�$WS��Ω��l�a�*�!�,Oq7�ĳ��uZ�E��*8#��D�!̖�g����t�EQ��\��n��?4���so�6e�tK�>�G�2�@K���j��_�<�M��Z��ע>�oaC 5��8��ظL*��`�D�".���]d�%�P0��T0�H�"�8n�7~,��/L��J�Jg�B�DBdTRl��$b��%����,�����-���+$��0(�+S���{�	U����V�(�GkVW�"�|̧3L��H|�������[��.e1/��~۹�@��ƕڦ{#8&�c�Q1E���IY��j�+�20'Ș`����3���r�j��;��L��n���S��2�y�V+
oM%gҍO3��AX	`�4d4�HXc)���5sR�3વ��"D�u )�Q��sױ��d�QB�ʻ8�5R�L}�/��d��I��4����_1�c��TO��.9F�+��HjQ����̈́��'���]8�3t�N���mbԙ"�����[YQղ|��M��'H��6K�v�x�W=SJ�9�0���n,���B�̇�y��"9�M�ዌշ�]J���yv�q�=2	Ɣ�D�H�8 g���*�޵�tC�]h0�	�B�_O%�x��-Q�Q>���D(i\�Ls��K|�˃���%�!�Yȁ��e�͑	�J�(�h菄���&�V�-13>#[n�Q�Ц�Dy GP0��kp�-��G��o~��|8�.Y4.5�+<ź�� ��B�ɐ^U��WZ���(3H�zϴʅۙ!���(�oTn�*��b:��;���4�A�=���C�x���u���gN��d��@2t�� �׊���{��*#���_!�_��C�?����,�cJ�ai��m� �x{k��p�B�������5��3D1.�_IA�hߪ��0�U�4PO��w+5�<5ȷ�F�o���<,��g*:�u���L�^$viNϽ)���v��#:�߇�#��C���[]���7m��D�}�Y��O-^���ܤ�Q���[�brzr�6>;�&��S�dx���iK����Y�I��G�am�Y�K���k�F��o��-�����U��`�}��1ܒ���tECg,�֩�	B�2h�':��(;�c"V�~�'$-"K�[se��Y�a͕R����]��S��6�������!{A�HS�_fL���A�w^xW��V�;�&��gW��Z꿈ws:T譗��/\�J1U��C8�������f/=�+	�����%��#���b.2�!