// D8M_QSYS.v

// Generated using ACDS version 15.0 145

`timescale 1 ps / 1 ps
module D8M_QSYS (
		input  wire        alt_vip_itc_0_clocked_video_vid_clk,         //       alt_vip_itc_0_clocked_video.vid_clk
		output wire [23:0] alt_vip_itc_0_clocked_video_vid_data,        //                                  .vid_data
		output wire        alt_vip_itc_0_clocked_video_underflow,       //                                  .underflow
		output wire        alt_vip_itc_0_clocked_video_vid_datavalid,   //                                  .vid_datavalid
		output wire        alt_vip_itc_0_clocked_video_vid_v_sync,      //                                  .vid_v_sync
		output wire        alt_vip_itc_0_clocked_video_vid_h_sync,      //                                  .vid_h_sync
		output wire        alt_vip_itc_0_clocked_video_vid_f,           //                                  .vid_f
		output wire        alt_vip_itc_0_clocked_video_vid_h,           //                                  .vid_h
		output wire        alt_vip_itc_0_clocked_video_vid_v,           //                                  .vid_v
		input  wire        external_clk50_clk,                          //                    external_clk50.clk
		input  wire        external_reset_reset_n,                      //                    external_reset.reset_n
		input  wire        hdmi_tx_int_n_external_connection_export,    // hdmi_tx_int_n_external_connection.export
		inout  wire        i2c_opencores_camera_export_scl_pad_io,      //       i2c_opencores_camera_export.scl_pad_io
		inout  wire        i2c_opencores_camera_export_sda_pad_io,      //                                  .sda_pad_io
		inout  wire        i2c_opencores_mipi_export_scl_pad_io,        //         i2c_opencores_mipi_export.scl_pad_io
		inout  wire        i2c_opencores_mipi_export_sda_pad_io,        //                                  .sda_pad_io
		output wire        i2c_scl_external_connection_export,          //       i2c_scl_external_connection.export
		inout  wire        i2c_sda_external_connection_export,          //       i2c_sda_external_connection.export
		input  wire [3:0]  key_external_connection_export,              //           key_external_connection.export
		input  wire        mem_if_lpddr2_emif_pll_ref_clk_clk,          //    mem_if_lpddr2_emif_pll_ref_clk.clk
		output wire        mem_if_lpddr2_emif_status_local_init_done,   //         mem_if_lpddr2_emif_status.local_init_done
		output wire        mem_if_lpddr2_emif_status_local_cal_success, //                                  .local_cal_success
		output wire        mem_if_lpddr2_emif_status_local_cal_fail,    //                                  .local_cal_fail
		output wire [9:0]  memory_mem_ca,                               //                            memory.mem_ca
		output wire [0:0]  memory_mem_ck,                               //                                  .mem_ck
		output wire [0:0]  memory_mem_ck_n,                             //                                  .mem_ck_n
		output wire [0:0]  memory_mem_cke,                              //                                  .mem_cke
		output wire [0:0]  memory_mem_cs_n,                             //                                  .mem_cs_n
		output wire [3:0]  memory_mem_dm,                               //                                  .mem_dm
		inout  wire [31:0] memory_mem_dq,                               //                                  .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                              //                                  .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                            //                                  .mem_dqs_n
		output wire        mipi_pwdn_n_external_connection_export,      //   mipi_pwdn_n_external_connection.export
		output wire        mipi_reset_n_external_connection_export,     //  mipi_reset_n_external_connection.export
		input  wire        oct_rzqin,                                   //                               oct.rzqin
		inout  wire        terasic_auto_focus_0_conduit_vcm_i2c_sda,    //      terasic_auto_focus_0_conduit.vcm_i2c_sda
		input  wire        terasic_auto_focus_0_conduit_clk50,          //                                  .clk50
		inout  wire        terasic_auto_focus_0_conduit_vcm_i2c_scl,    //                                  .vcm_i2c_scl
		input  wire [11:0] terasic_camera_0_conduit_end_D,              //      terasic_camera_0_conduit_end.D
		input  wire        terasic_camera_0_conduit_end_FVAL,           //                                  .FVAL
		input  wire        terasic_camera_0_conduit_end_LVAL,           //                                  .LVAL
		input  wire        terasic_camera_0_conduit_end_PIXCLK          //                                  .PIXCLK
	);

	wire          terasic_camera_0_avalon_streaming_source_valid;                    // TERASIC_CAMERA_0:st_valid -> alt_vip_vfb_0:din_valid
	wire   [23:0] terasic_camera_0_avalon_streaming_source_data;                     // TERASIC_CAMERA_0:st_data -> alt_vip_vfb_0:din_data
	wire          terasic_camera_0_avalon_streaming_source_ready;                    // alt_vip_vfb_0:din_ready -> TERASIC_CAMERA_0:st_ready
	wire          terasic_camera_0_avalon_streaming_source_startofpacket;            // TERASIC_CAMERA_0:st_sop -> alt_vip_vfb_0:din_startofpacket
	wire          terasic_camera_0_avalon_streaming_source_endofpacket;              // TERASIC_CAMERA_0:st_eop -> alt_vip_vfb_0:din_endofpacket
	wire          alt_vip_vfb_0_dout_valid;                                          // alt_vip_vfb_0:dout_valid -> TERASIC_AUTO_FOCUS_0:sink_valid
	wire   [23:0] alt_vip_vfb_0_dout_data;                                           // alt_vip_vfb_0:dout_data -> TERASIC_AUTO_FOCUS_0:sink_data
	wire          alt_vip_vfb_0_dout_ready;                                          // TERASIC_AUTO_FOCUS_0:sink_ready -> alt_vip_vfb_0:dout_ready
	wire          alt_vip_vfb_0_dout_startofpacket;                                  // alt_vip_vfb_0:dout_startofpacket -> TERASIC_AUTO_FOCUS_0:sink_sop
	wire          alt_vip_vfb_0_dout_endofpacket;                                    // alt_vip_vfb_0:dout_endofpacket -> TERASIC_AUTO_FOCUS_0:sink_eop
	wire          terasic_auto_focus_0_dout_valid;                                   // TERASIC_AUTO_FOCUS_0:source_valid -> alt_vip_itc_0:is_valid
	wire   [23:0] terasic_auto_focus_0_dout_data;                                    // TERASIC_AUTO_FOCUS_0:source_data -> alt_vip_itc_0:is_data
	wire          terasic_auto_focus_0_dout_ready;                                   // alt_vip_itc_0:is_ready -> TERASIC_AUTO_FOCUS_0:source_ready
	wire          terasic_auto_focus_0_dout_startofpacket;                           // TERASIC_AUTO_FOCUS_0:source_sop -> alt_vip_itc_0:is_sop
	wire          terasic_auto_focus_0_dout_endofpacket;                             // TERASIC_AUTO_FOCUS_0:source_eop -> alt_vip_itc_0:is_eop
	wire          mem_if_lpddr2_emif_afi_clk_clk;                                    // mem_if_lpddr2_emif:afi_clk -> [TERASIC_AUTO_FOCUS_0:clk, TERASIC_CAMERA_0:clk, alt_vip_itc_0:is_clk, alt_vip_vfb_0:clock, mm_interconnect_0:mem_if_lpddr2_emif_afi_clk_clk, mm_interconnect_1:mem_if_lpddr2_emif_afi_clk_clk, rst_controller:clk]
	wire   [31:0] nios2_qsys_data_master_readdata;                                   // mm_interconnect_0:nios2_qsys_data_master_readdata -> nios2_qsys:d_readdata
	wire          nios2_qsys_data_master_waitrequest;                                // mm_interconnect_0:nios2_qsys_data_master_waitrequest -> nios2_qsys:d_waitrequest
	wire          nios2_qsys_data_master_debugaccess;                                // nios2_qsys:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_qsys_data_master_debugaccess
	wire   [19:0] nios2_qsys_data_master_address;                                    // nios2_qsys:d_address -> mm_interconnect_0:nios2_qsys_data_master_address
	wire    [3:0] nios2_qsys_data_master_byteenable;                                 // nios2_qsys:d_byteenable -> mm_interconnect_0:nios2_qsys_data_master_byteenable
	wire          nios2_qsys_data_master_read;                                       // nios2_qsys:d_read -> mm_interconnect_0:nios2_qsys_data_master_read
	wire          nios2_qsys_data_master_readdatavalid;                              // mm_interconnect_0:nios2_qsys_data_master_readdatavalid -> nios2_qsys:d_readdatavalid
	wire          nios2_qsys_data_master_write;                                      // nios2_qsys:d_write -> mm_interconnect_0:nios2_qsys_data_master_write
	wire   [31:0] nios2_qsys_data_master_writedata;                                  // nios2_qsys:d_writedata -> mm_interconnect_0:nios2_qsys_data_master_writedata
	wire   [31:0] nios2_qsys_instruction_master_readdata;                            // mm_interconnect_0:nios2_qsys_instruction_master_readdata -> nios2_qsys:i_readdata
	wire          nios2_qsys_instruction_master_waitrequest;                         // mm_interconnect_0:nios2_qsys_instruction_master_waitrequest -> nios2_qsys:i_waitrequest
	wire   [19:0] nios2_qsys_instruction_master_address;                             // nios2_qsys:i_address -> mm_interconnect_0:nios2_qsys_instruction_master_address
	wire          nios2_qsys_instruction_master_read;                                // nios2_qsys:i_read -> mm_interconnect_0:nios2_qsys_instruction_master_read
	wire          nios2_qsys_instruction_master_readdatavalid;                       // mm_interconnect_0:nios2_qsys_instruction_master_readdatavalid -> nios2_qsys:i_readdatavalid
	wire          mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;          // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire   [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;            // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire          mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;         // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire    [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;             // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire          mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;                // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire          mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;               // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire   [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;           // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire          mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_chipselect;  // mm_interconnect_0:i2c_opencores_camera_avalon_slave_0_chipselect -> i2c_opencores_camera:wb_stb_i
	wire    [7:0] mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_readdata;    // i2c_opencores_camera:wb_dat_o -> mm_interconnect_0:i2c_opencores_camera_avalon_slave_0_readdata
	wire          mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_waitrequest; // i2c_opencores_camera:wb_ack_o -> mm_interconnect_0:i2c_opencores_camera_avalon_slave_0_waitrequest
	wire    [2:0] mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_address;     // mm_interconnect_0:i2c_opencores_camera_avalon_slave_0_address -> i2c_opencores_camera:wb_adr_i
	wire          mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_write;       // mm_interconnect_0:i2c_opencores_camera_avalon_slave_0_write -> i2c_opencores_camera:wb_we_i
	wire    [7:0] mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_writedata;   // mm_interconnect_0:i2c_opencores_camera_avalon_slave_0_writedata -> i2c_opencores_camera:wb_dat_i
	wire          mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_chipselect;    // mm_interconnect_0:i2c_opencores_mipi_avalon_slave_0_chipselect -> i2c_opencores_mipi:wb_stb_i
	wire    [7:0] mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_readdata;      // i2c_opencores_mipi:wb_dat_o -> mm_interconnect_0:i2c_opencores_mipi_avalon_slave_0_readdata
	wire          mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_waitrequest;   // i2c_opencores_mipi:wb_ack_o -> mm_interconnect_0:i2c_opencores_mipi_avalon_slave_0_waitrequest
	wire    [2:0] mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_address;       // mm_interconnect_0:i2c_opencores_mipi_avalon_slave_0_address -> i2c_opencores_mipi:wb_adr_i
	wire          mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_write;         // mm_interconnect_0:i2c_opencores_mipi_avalon_slave_0_write -> i2c_opencores_mipi:wb_we_i
	wire    [7:0] mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_writedata;     // mm_interconnect_0:i2c_opencores_mipi_avalon_slave_0_writedata -> i2c_opencores_mipi:wb_dat_i
	wire   [31:0] mm_interconnect_0_sysid_qsys_control_slave_readdata;               // sysid_qsys:readdata -> mm_interconnect_0:sysid_qsys_control_slave_readdata
	wire    [0:0] mm_interconnect_0_sysid_qsys_control_slave_address;                // mm_interconnect_0:sysid_qsys_control_slave_address -> sysid_qsys:address
	wire   [31:0] mm_interconnect_0_nios2_qsys_jtag_debug_module_readdata;           // nios2_qsys:jtag_debug_module_readdata -> mm_interconnect_0:nios2_qsys_jtag_debug_module_readdata
	wire          mm_interconnect_0_nios2_qsys_jtag_debug_module_waitrequest;        // nios2_qsys:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_qsys_jtag_debug_module_waitrequest
	wire          mm_interconnect_0_nios2_qsys_jtag_debug_module_debugaccess;        // mm_interconnect_0:nios2_qsys_jtag_debug_module_debugaccess -> nios2_qsys:jtag_debug_module_debugaccess
	wire    [8:0] mm_interconnect_0_nios2_qsys_jtag_debug_module_address;            // mm_interconnect_0:nios2_qsys_jtag_debug_module_address -> nios2_qsys:jtag_debug_module_address
	wire          mm_interconnect_0_nios2_qsys_jtag_debug_module_read;               // mm_interconnect_0:nios2_qsys_jtag_debug_module_read -> nios2_qsys:jtag_debug_module_read
	wire    [3:0] mm_interconnect_0_nios2_qsys_jtag_debug_module_byteenable;         // mm_interconnect_0:nios2_qsys_jtag_debug_module_byteenable -> nios2_qsys:jtag_debug_module_byteenable
	wire          mm_interconnect_0_nios2_qsys_jtag_debug_module_write;              // mm_interconnect_0:nios2_qsys_jtag_debug_module_write -> nios2_qsys:jtag_debug_module_write
	wire   [31:0] mm_interconnect_0_nios2_qsys_jtag_debug_module_writedata;          // mm_interconnect_0:nios2_qsys_jtag_debug_module_writedata -> nios2_qsys:jtag_debug_module_writedata
	wire          mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_chipselect;         // mm_interconnect_0:TERASIC_AUTO_FOCUS_0_mm_ctrl_chipselect -> TERASIC_AUTO_FOCUS_0:s_chipselect
	wire   [31:0] mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_readdata;           // TERASIC_AUTO_FOCUS_0:s_readdata -> mm_interconnect_0:TERASIC_AUTO_FOCUS_0_mm_ctrl_readdata
	wire    [2:0] mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_address;            // mm_interconnect_0:TERASIC_AUTO_FOCUS_0_mm_ctrl_address -> TERASIC_AUTO_FOCUS_0:s_address
	wire          mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_read;               // mm_interconnect_0:TERASIC_AUTO_FOCUS_0_mm_ctrl_read -> TERASIC_AUTO_FOCUS_0:s_read
	wire          mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_write;              // mm_interconnect_0:TERASIC_AUTO_FOCUS_0_mm_ctrl_write -> TERASIC_AUTO_FOCUS_0:s_write
	wire   [31:0] mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_writedata;          // mm_interconnect_0:TERASIC_AUTO_FOCUS_0_mm_ctrl_writedata -> TERASIC_AUTO_FOCUS_0:s_writedata
	wire          mm_interconnect_0_onchip_memory2_s1_chipselect;                    // mm_interconnect_0:onchip_memory2_s1_chipselect -> onchip_memory2:chipselect
	wire   [31:0] mm_interconnect_0_onchip_memory2_s1_readdata;                      // onchip_memory2:readdata -> mm_interconnect_0:onchip_memory2_s1_readdata
	wire   [15:0] mm_interconnect_0_onchip_memory2_s1_address;                       // mm_interconnect_0:onchip_memory2_s1_address -> onchip_memory2:address
	wire    [3:0] mm_interconnect_0_onchip_memory2_s1_byteenable;                    // mm_interconnect_0:onchip_memory2_s1_byteenable -> onchip_memory2:byteenable
	wire          mm_interconnect_0_onchip_memory2_s1_write;                         // mm_interconnect_0:onchip_memory2_s1_write -> onchip_memory2:write
	wire   [31:0] mm_interconnect_0_onchip_memory2_s1_writedata;                     // mm_interconnect_0:onchip_memory2_s1_writedata -> onchip_memory2:writedata
	wire          mm_interconnect_0_onchip_memory2_s1_clken;                         // mm_interconnect_0:onchip_memory2_s1_clken -> onchip_memory2:clken
	wire          mm_interconnect_0_timer_s1_chipselect;                             // mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	wire   [15:0] mm_interconnect_0_timer_s1_readdata;                               // timer:readdata -> mm_interconnect_0:timer_s1_readdata
	wire    [2:0] mm_interconnect_0_timer_s1_address;                                // mm_interconnect_0:timer_s1_address -> timer:address
	wire          mm_interconnect_0_timer_s1_write;                                  // mm_interconnect_0:timer_s1_write -> timer:write_n
	wire   [15:0] mm_interconnect_0_timer_s1_writedata;                              // mm_interconnect_0:timer_s1_writedata -> timer:writedata
	wire          mm_interconnect_0_i2c_sda_s1_chipselect;                           // mm_interconnect_0:i2c_sda_s1_chipselect -> i2c_sda:chipselect
	wire   [31:0] mm_interconnect_0_i2c_sda_s1_readdata;                             // i2c_sda:readdata -> mm_interconnect_0:i2c_sda_s1_readdata
	wire    [1:0] mm_interconnect_0_i2c_sda_s1_address;                              // mm_interconnect_0:i2c_sda_s1_address -> i2c_sda:address
	wire          mm_interconnect_0_i2c_sda_s1_write;                                // mm_interconnect_0:i2c_sda_s1_write -> i2c_sda:write_n
	wire   [31:0] mm_interconnect_0_i2c_sda_s1_writedata;                            // mm_interconnect_0:i2c_sda_s1_writedata -> i2c_sda:writedata
	wire          mm_interconnect_0_i2c_scl_s1_chipselect;                           // mm_interconnect_0:i2c_scl_s1_chipselect -> i2c_scl:chipselect
	wire   [31:0] mm_interconnect_0_i2c_scl_s1_readdata;                             // i2c_scl:readdata -> mm_interconnect_0:i2c_scl_s1_readdata
	wire    [1:0] mm_interconnect_0_i2c_scl_s1_address;                              // mm_interconnect_0:i2c_scl_s1_address -> i2c_scl:address
	wire          mm_interconnect_0_i2c_scl_s1_write;                                // mm_interconnect_0:i2c_scl_s1_write -> i2c_scl:write_n
	wire   [31:0] mm_interconnect_0_i2c_scl_s1_writedata;                            // mm_interconnect_0:i2c_scl_s1_writedata -> i2c_scl:writedata
	wire          mm_interconnect_0_hdmi_tx_int_n_s1_chipselect;                     // mm_interconnect_0:hdmi_tx_int_n_s1_chipselect -> hdmi_tx_int_n:chipselect
	wire   [31:0] mm_interconnect_0_hdmi_tx_int_n_s1_readdata;                       // hdmi_tx_int_n:readdata -> mm_interconnect_0:hdmi_tx_int_n_s1_readdata
	wire    [1:0] mm_interconnect_0_hdmi_tx_int_n_s1_address;                        // mm_interconnect_0:hdmi_tx_int_n_s1_address -> hdmi_tx_int_n:address
	wire          mm_interconnect_0_hdmi_tx_int_n_s1_write;                          // mm_interconnect_0:hdmi_tx_int_n_s1_write -> hdmi_tx_int_n:write_n
	wire   [31:0] mm_interconnect_0_hdmi_tx_int_n_s1_writedata;                      // mm_interconnect_0:hdmi_tx_int_n_s1_writedata -> hdmi_tx_int_n:writedata
	wire          mm_interconnect_0_mipi_pwdn_n_s1_chipselect;                       // mm_interconnect_0:mipi_pwdn_n_s1_chipselect -> mipi_pwdn_n:chipselect
	wire   [31:0] mm_interconnect_0_mipi_pwdn_n_s1_readdata;                         // mipi_pwdn_n:readdata -> mm_interconnect_0:mipi_pwdn_n_s1_readdata
	wire    [1:0] mm_interconnect_0_mipi_pwdn_n_s1_address;                          // mm_interconnect_0:mipi_pwdn_n_s1_address -> mipi_pwdn_n:address
	wire          mm_interconnect_0_mipi_pwdn_n_s1_write;                            // mm_interconnect_0:mipi_pwdn_n_s1_write -> mipi_pwdn_n:write_n
	wire   [31:0] mm_interconnect_0_mipi_pwdn_n_s1_writedata;                        // mm_interconnect_0:mipi_pwdn_n_s1_writedata -> mipi_pwdn_n:writedata
	wire          mm_interconnect_0_mipi_reset_n_s1_chipselect;                      // mm_interconnect_0:mipi_reset_n_s1_chipselect -> mipi_reset_n:chipselect
	wire   [31:0] mm_interconnect_0_mipi_reset_n_s1_readdata;                        // mipi_reset_n:readdata -> mm_interconnect_0:mipi_reset_n_s1_readdata
	wire    [1:0] mm_interconnect_0_mipi_reset_n_s1_address;                         // mm_interconnect_0:mipi_reset_n_s1_address -> mipi_reset_n:address
	wire          mm_interconnect_0_mipi_reset_n_s1_write;                           // mm_interconnect_0:mipi_reset_n_s1_write -> mipi_reset_n:write_n
	wire   [31:0] mm_interconnect_0_mipi_reset_n_s1_writedata;                       // mm_interconnect_0:mipi_reset_n_s1_writedata -> mipi_reset_n:writedata
	wire   [31:0] mm_interconnect_0_key_s1_readdata;                                 // key:readdata -> mm_interconnect_0:key_s1_readdata
	wire    [1:0] mm_interconnect_0_key_s1_address;                                  // mm_interconnect_0:key_s1_address -> key:address
	wire          alt_vip_vfb_0_read_master_waitrequest;                             // mm_interconnect_1:alt_vip_vfb_0_read_master_waitrequest -> alt_vip_vfb_0:read_master_av_waitrequest
	wire  [127:0] alt_vip_vfb_0_read_master_readdata;                                // mm_interconnect_1:alt_vip_vfb_0_read_master_readdata -> alt_vip_vfb_0:read_master_av_readdata
	wire   [31:0] alt_vip_vfb_0_read_master_address;                                 // alt_vip_vfb_0:read_master_av_address -> mm_interconnect_1:alt_vip_vfb_0_read_master_address
	wire          alt_vip_vfb_0_read_master_read;                                    // alt_vip_vfb_0:read_master_av_read -> mm_interconnect_1:alt_vip_vfb_0_read_master_read
	wire          alt_vip_vfb_0_read_master_readdatavalid;                           // mm_interconnect_1:alt_vip_vfb_0_read_master_readdatavalid -> alt_vip_vfb_0:read_master_av_readdatavalid
	wire    [2:0] alt_vip_vfb_0_read_master_burstcount;                              // alt_vip_vfb_0:read_master_av_burstcount -> mm_interconnect_1:alt_vip_vfb_0_read_master_burstcount
	wire          alt_vip_vfb_0_write_master_waitrequest;                            // mm_interconnect_1:alt_vip_vfb_0_write_master_waitrequest -> alt_vip_vfb_0:write_master_av_waitrequest
	wire   [31:0] alt_vip_vfb_0_write_master_address;                                // alt_vip_vfb_0:write_master_av_address -> mm_interconnect_1:alt_vip_vfb_0_write_master_address
	wire          alt_vip_vfb_0_write_master_write;                                  // alt_vip_vfb_0:write_master_av_write -> mm_interconnect_1:alt_vip_vfb_0_write_master_write
	wire  [127:0] alt_vip_vfb_0_write_master_writedata;                              // alt_vip_vfb_0:write_master_av_writedata -> mm_interconnect_1:alt_vip_vfb_0_write_master_writedata
	wire    [2:0] alt_vip_vfb_0_write_master_burstcount;                             // alt_vip_vfb_0:write_master_av_burstcount -> mm_interconnect_1:alt_vip_vfb_0_write_master_burstcount
	wire          mm_interconnect_1_mem_if_lpddr2_emif_avl_beginbursttransfer;       // mm_interconnect_1:mem_if_lpddr2_emif_avl_beginbursttransfer -> mem_if_lpddr2_emif:avl_burstbegin
	wire  [127:0] mm_interconnect_1_mem_if_lpddr2_emif_avl_readdata;                 // mem_if_lpddr2_emif:avl_rdata -> mm_interconnect_1:mem_if_lpddr2_emif_avl_readdata
	wire          mm_interconnect_1_mem_if_lpddr2_emif_avl_waitrequest;              // mem_if_lpddr2_emif:avl_ready -> mm_interconnect_1:mem_if_lpddr2_emif_avl_waitrequest
	wire   [21:0] mm_interconnect_1_mem_if_lpddr2_emif_avl_address;                  // mm_interconnect_1:mem_if_lpddr2_emif_avl_address -> mem_if_lpddr2_emif:avl_addr
	wire          mm_interconnect_1_mem_if_lpddr2_emif_avl_read;                     // mm_interconnect_1:mem_if_lpddr2_emif_avl_read -> mem_if_lpddr2_emif:avl_read_req
	wire   [15:0] mm_interconnect_1_mem_if_lpddr2_emif_avl_byteenable;               // mm_interconnect_1:mem_if_lpddr2_emif_avl_byteenable -> mem_if_lpddr2_emif:avl_be
	wire          mm_interconnect_1_mem_if_lpddr2_emif_avl_readdatavalid;            // mem_if_lpddr2_emif:avl_rdata_valid -> mm_interconnect_1:mem_if_lpddr2_emif_avl_readdatavalid
	wire          mm_interconnect_1_mem_if_lpddr2_emif_avl_write;                    // mm_interconnect_1:mem_if_lpddr2_emif_avl_write -> mem_if_lpddr2_emif:avl_write_req
	wire  [127:0] mm_interconnect_1_mem_if_lpddr2_emif_avl_writedata;                // mm_interconnect_1:mem_if_lpddr2_emif_avl_writedata -> mem_if_lpddr2_emif:avl_wdata
	wire    [5:0] mm_interconnect_1_mem_if_lpddr2_emif_avl_burstcount;               // mm_interconnect_1:mem_if_lpddr2_emif_avl_burstcount -> mem_if_lpddr2_emif:avl_size
	wire          irq_mapper_receiver0_irq;                                          // i2c_opencores_mipi:wb_inta_o -> irq_mapper:receiver0_irq
	wire          irq_mapper_receiver1_irq;                                          // i2c_opencores_camera:wb_inta_o -> irq_mapper:receiver1_irq
	wire          irq_mapper_receiver2_irq;                                          // timer:irq -> irq_mapper:receiver2_irq
	wire          irq_mapper_receiver3_irq;                                          // jtag_uart:av_irq -> irq_mapper:receiver3_irq
	wire          irq_mapper_receiver4_irq;                                          // hdmi_tx_int_n:irq -> irq_mapper:receiver4_irq
	wire   [31:0] nios2_qsys_d_irq_irq;                                              // irq_mapper:sender_irq -> nios2_qsys:d_irq
	wire          rst_controller_reset_out_reset;                                    // rst_controller:reset_out -> [TERASIC_AUTO_FOCUS_0:reset_n, TERASIC_CAMERA_0:reset_n, alt_vip_itc_0:rst, alt_vip_vfb_0:reset, mm_interconnect_0:TERASIC_AUTO_FOCUS_0_reset_reset_bridge_in_reset_reset, mm_interconnect_1:alt_vip_vfb_0_reset_reset_bridge_in_reset_reset, mm_interconnect_1:mem_if_lpddr2_emif_soft_reset_reset_bridge_in_reset_reset]
	wire          rst_controller_001_reset_out_reset;                                // rst_controller_001:reset_out -> [hdmi_tx_int_n:reset_n, i2c_opencores_camera:wb_rst_i, i2c_opencores_mipi:wb_rst_i, i2c_scl:reset_n, i2c_sda:reset_n, jtag_uart:rst_n, key:reset_n, mipi_pwdn_n:reset_n, mipi_reset_n:reset_n, mm_interconnect_0:jtag_uart_reset_reset_bridge_in_reset_reset, onchip_memory2:reset, rst_translator:in_reset, sysid_qsys:reset_n, timer:reset_n]
	wire          rst_controller_001_reset_out_reset_req;                            // rst_controller_001:reset_req -> [onchip_memory2:reset_req, rst_translator:reset_req_in]
	wire          rst_controller_002_reset_out_reset;                                // rst_controller_002:reset_out -> [irq_mapper:reset, mm_interconnect_0:nios2_qsys_reset_n_reset_bridge_in_reset_reset, nios2_qsys:reset_n]
	wire          rst_controller_002_reset_out_reset_req;                            // rst_controller_002:reset_req -> [nios2_qsys:reset_req, rst_translator_001:reset_req_in]
	wire          nios2_qsys_jtag_debug_module_reset_reset;                          // nios2_qsys:jtag_debug_module_resetrequest -> rst_controller_002:reset_in1

	TERASIC_AUTO_FOCUS #(
		.VIDEO_W (1920),
		.VIDEO_H (1080)
	) terasic_auto_focus_0 (
		.clk          (mem_if_lpddr2_emif_afi_clk_clk),                            //   clock.clk
		.reset_n      (~rst_controller_reset_out_reset),                           //   reset.reset_n
		.s_chipselect (mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_chipselect), // mm_ctrl.chipselect
		.s_read       (mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_read),       //        .read
		.s_write      (mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_write),      //        .write
		.s_readdata   (mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_readdata),   //        .readdata
		.s_writedata  (mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_writedata),  //        .writedata
		.s_address    (mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_address),    //        .address
		.sink_data    (alt_vip_vfb_0_dout_data),                                   //     din.data
		.sink_valid   (alt_vip_vfb_0_dout_valid),                                  //        .valid
		.sink_ready   (alt_vip_vfb_0_dout_ready),                                  //        .ready
		.sink_sop     (alt_vip_vfb_0_dout_startofpacket),                          //        .startofpacket
		.sink_eop     (alt_vip_vfb_0_dout_endofpacket),                            //        .endofpacket
		.source_data  (terasic_auto_focus_0_dout_data),                            //    dout.data
		.source_valid (terasic_auto_focus_0_dout_valid),                           //        .valid
		.source_ready (terasic_auto_focus_0_dout_ready),                           //        .ready
		.source_sop   (terasic_auto_focus_0_dout_startofpacket),                   //        .startofpacket
		.source_eop   (terasic_auto_focus_0_dout_endofpacket),                     //        .endofpacket
		.vcm_i2c_sda  (terasic_auto_focus_0_conduit_vcm_i2c_sda),                  // Conduit.vcm_i2c_sda
		.clk50        (terasic_auto_focus_0_conduit_clk50),                        //        .clk50
		.vcm_i2c_scl  (terasic_auto_focus_0_conduit_vcm_i2c_scl)                   //        .vcm_i2c_scl
	);

	TERASIC_CAMERA #(
		.VIDEO_W (1920),
		.VIDEO_H (1080)
	) terasic_camera_0 (
		.clk           (mem_if_lpddr2_emif_afi_clk_clk),                         //             clock_reset.clk
		.reset_n       (~rst_controller_reset_out_reset),                        //       clock_reset_reset.reset_n
		.CAMERA_D      (terasic_camera_0_conduit_end_D),                         //             conduit_end.export
		.CAMERA_FVAL   (terasic_camera_0_conduit_end_FVAL),                      //                        .export
		.CAMERA_LVAL   (terasic_camera_0_conduit_end_LVAL),                      //                        .export
		.CAMERA_PIXCLK (terasic_camera_0_conduit_end_PIXCLK),                    //                        .export
		.st_data       (terasic_camera_0_avalon_streaming_source_data),          // avalon_streaming_source.data
		.st_sop        (terasic_camera_0_avalon_streaming_source_startofpacket), //                        .startofpacket
		.st_eop        (terasic_camera_0_avalon_streaming_source_endofpacket),   //                        .endofpacket
		.st_ready      (terasic_camera_0_avalon_streaming_source_ready),         //                        .ready
		.st_valid      (terasic_camera_0_avalon_streaming_source_valid)          //                        .valid
	);

	alt_vipitc131_IS2Vid #(
		.NUMBER_OF_COLOUR_PLANES       (3),
		.COLOUR_PLANES_ARE_IN_PARALLEL (1),
		.BPS                           (8),
		.INTERLACED                    (0),
		.H_ACTIVE_PIXELS               (1920),
		.V_ACTIVE_LINES                (1080),
		.ACCEPT_COLOURS_IN_SEQ         (0),
		.FIFO_DEPTH                    (3840),
		.CLOCKS_ARE_SAME               (0),
		.USE_CONTROL                   (0),
		.NO_OF_MODES                   (1),
		.THRESHOLD                     (1919),
		.STD_WIDTH                     (1),
		.GENERATE_SYNC                 (0),
		.USE_EMBEDDED_SYNCS            (0),
		.AP_LINE                       (0),
		.V_BLANK                       (0),
		.H_BLANK                       (0),
		.H_SYNC_LENGTH                 (44),
		.H_FRONT_PORCH                 (88),
		.H_BACK_PORCH                  (148),
		.V_SYNC_LENGTH                 (5),
		.V_FRONT_PORCH                 (4),
		.V_BACK_PORCH                  (36),
		.F_RISING_EDGE                 (0),
		.F_FALLING_EDGE                (0),
		.FIELD0_V_RISING_EDGE          (0),
		.FIELD0_V_BLANK                (0),
		.FIELD0_V_SYNC_LENGTH          (0),
		.FIELD0_V_FRONT_PORCH          (0),
		.FIELD0_V_BACK_PORCH           (0),
		.ANC_LINE                      (0),
		.FIELD0_ANC_LINE               (0)
	) alt_vip_itc_0 (
		.is_clk        (mem_if_lpddr2_emif_afi_clk_clk),            //       is_clk_rst.clk
		.rst           (rst_controller_reset_out_reset),            // is_clk_rst_reset.reset
		.is_data       (terasic_auto_focus_0_dout_data),            //              din.data
		.is_valid      (terasic_auto_focus_0_dout_valid),           //                 .valid
		.is_ready      (terasic_auto_focus_0_dout_ready),           //                 .ready
		.is_sop        (terasic_auto_focus_0_dout_startofpacket),   //                 .startofpacket
		.is_eop        (terasic_auto_focus_0_dout_endofpacket),     //                 .endofpacket
		.vid_clk       (alt_vip_itc_0_clocked_video_vid_clk),       //    clocked_video.export
		.vid_data      (alt_vip_itc_0_clocked_video_vid_data),      //                 .export
		.underflow     (alt_vip_itc_0_clocked_video_underflow),     //                 .export
		.vid_datavalid (alt_vip_itc_0_clocked_video_vid_datavalid), //                 .export
		.vid_v_sync    (alt_vip_itc_0_clocked_video_vid_v_sync),    //                 .export
		.vid_h_sync    (alt_vip_itc_0_clocked_video_vid_h_sync),    //                 .export
		.vid_f         (alt_vip_itc_0_clocked_video_vid_f),         //                 .export
		.vid_h         (alt_vip_itc_0_clocked_video_vid_h),         //                 .export
		.vid_v         (alt_vip_itc_0_clocked_video_vid_v)          //                 .export
	);

	D8M_QSYS_alt_vip_vfb_0 alt_vip_vfb_0 (
		.clock                        (mem_if_lpddr2_emif_afi_clk_clk),                         //        clock.clk
		.reset                        (rst_controller_reset_out_reset),                         //        reset.reset
		.din_ready                    (terasic_camera_0_avalon_streaming_source_ready),         //          din.ready
		.din_valid                    (terasic_camera_0_avalon_streaming_source_valid),         //             .valid
		.din_data                     (terasic_camera_0_avalon_streaming_source_data),          //             .data
		.din_startofpacket            (terasic_camera_0_avalon_streaming_source_startofpacket), //             .startofpacket
		.din_endofpacket              (terasic_camera_0_avalon_streaming_source_endofpacket),   //             .endofpacket
		.dout_ready                   (alt_vip_vfb_0_dout_ready),                               //         dout.ready
		.dout_valid                   (alt_vip_vfb_0_dout_valid),                               //             .valid
		.dout_data                    (alt_vip_vfb_0_dout_data),                                //             .data
		.dout_startofpacket           (alt_vip_vfb_0_dout_startofpacket),                       //             .startofpacket
		.dout_endofpacket             (alt_vip_vfb_0_dout_endofpacket),                         //             .endofpacket
		.read_master_av_address       (alt_vip_vfb_0_read_master_address),                      //  read_master.address
		.read_master_av_read          (alt_vip_vfb_0_read_master_read),                         //             .read
		.read_master_av_waitrequest   (alt_vip_vfb_0_read_master_waitrequest),                  //             .waitrequest
		.read_master_av_readdatavalid (alt_vip_vfb_0_read_master_readdatavalid),                //             .readdatavalid
		.read_master_av_readdata      (alt_vip_vfb_0_read_master_readdata),                     //             .readdata
		.read_master_av_burstcount    (alt_vip_vfb_0_read_master_burstcount),                   //             .burstcount
		.write_master_av_address      (alt_vip_vfb_0_write_master_address),                     // write_master.address
		.write_master_av_write        (alt_vip_vfb_0_write_master_write),                       //             .write
		.write_master_av_writedata    (alt_vip_vfb_0_write_master_writedata),                   //             .writedata
		.write_master_av_waitrequest  (alt_vip_vfb_0_write_master_waitrequest),                 //             .waitrequest
		.write_master_av_burstcount   (alt_vip_vfb_0_write_master_burstcount)                   //             .burstcount
	);

	D8M_QSYS_hdmi_tx_int_n hdmi_tx_int_n (
		.clk        (external_clk50_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_hdmi_tx_int_n_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hdmi_tx_int_n_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hdmi_tx_int_n_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hdmi_tx_int_n_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hdmi_tx_int_n_s1_readdata),   //                    .readdata
		.in_port    (hdmi_tx_int_n_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver4_irq)                       //                 irq.irq
	);

	i2c_opencores i2c_opencores_camera (
		.wb_clk_i   (external_clk50_clk),                                                //            clock.clk
		.wb_rst_i   (rst_controller_001_reset_out_reset),                                //      clock_reset.reset
		.scl_pad_io (i2c_opencores_camera_export_scl_pad_io),                            //           export.export
		.sda_pad_io (i2c_opencores_camera_export_sda_pad_io),                            //                 .export
		.wb_adr_i   (mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_address),     //   avalon_slave_0.address
		.wb_dat_i   (mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_writedata),   //                 .writedata
		.wb_dat_o   (mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_readdata),    //                 .readdata
		.wb_we_i    (mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_write),       //                 .write
		.wb_stb_i   (mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_chipselect),  //                 .chipselect
		.wb_ack_o   (mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_waitrequest), //                 .waitrequest_n
		.wb_inta_o  (irq_mapper_receiver1_irq)                                           // interrupt_sender.irq
	);

	i2c_opencores i2c_opencores_mipi (
		.wb_clk_i   (external_clk50_clk),                                              //            clock.clk
		.wb_rst_i   (rst_controller_001_reset_out_reset),                              //      clock_reset.reset
		.scl_pad_io (i2c_opencores_mipi_export_scl_pad_io),                            //           export.export
		.sda_pad_io (i2c_opencores_mipi_export_sda_pad_io),                            //                 .export
		.wb_adr_i   (mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_address),     //   avalon_slave_0.address
		.wb_dat_i   (mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_writedata),   //                 .writedata
		.wb_dat_o   (mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_readdata),    //                 .readdata
		.wb_we_i    (mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_write),       //                 .write
		.wb_stb_i   (mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_chipselect),  //                 .chipselect
		.wb_ack_o   (mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_waitrequest), //                 .waitrequest_n
		.wb_inta_o  (irq_mapper_receiver0_irq)                                         // interrupt_sender.irq
	);

	D8M_QSYS_i2c_scl i2c_scl (
		.clk        (external_clk50_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_i2c_scl_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_i2c_scl_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_i2c_scl_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_i2c_scl_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_i2c_scl_s1_readdata),   //                    .readdata
		.out_port   (i2c_scl_external_connection_export)       // external_connection.export
	);

	D8M_QSYS_i2c_sda i2c_sda (
		.clk        (external_clk50_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_i2c_sda_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_i2c_sda_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_i2c_sda_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_i2c_sda_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_i2c_sda_s1_readdata),   //                    .readdata
		.bidir_port (i2c_sda_external_connection_export)       // external_connection.export
	);

	D8M_QSYS_jtag_uart jtag_uart (
		.clk            (external_clk50_clk),                                        //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver3_irq)                                   //               irq.irq
	);

	D8M_QSYS_key key (
		.clk      (external_clk50_clk),                  //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset), //               reset.reset_n
		.address  (mm_interconnect_0_key_s1_address),    //                  s1.address
		.readdata (mm_interconnect_0_key_s1_readdata),   //                    .readdata
		.in_port  (key_external_connection_export)       // external_connection.export
	);

	D8M_QSYS_mem_if_lpddr2_emif mem_if_lpddr2_emif (
		.pll_ref_clk               (mem_if_lpddr2_emif_pll_ref_clk_clk),                          //      pll_ref_clk.clk
		.global_reset_n            (external_reset_reset_n),                                      //     global_reset.reset_n
		.soft_reset_n              (external_reset_reset_n),                                      //       soft_reset.reset_n
		.afi_clk                   (mem_if_lpddr2_emif_afi_clk_clk),                              //          afi_clk.clk
		.afi_half_clk              (),                                                            //     afi_half_clk.clk
		.afi_reset_n               (),                                                            //        afi_reset.reset_n
		.afi_reset_export_n        (),                                                            // afi_reset_export.reset_n
		.mem_ca                    (memory_mem_ca),                                               //           memory.mem_ca
		.mem_ck                    (memory_mem_ck),                                               //                 .mem_ck
		.mem_ck_n                  (memory_mem_ck_n),                                             //                 .mem_ck_n
		.mem_cke                   (memory_mem_cke),                                              //                 .mem_cke
		.mem_cs_n                  (memory_mem_cs_n),                                             //                 .mem_cs_n
		.mem_dm                    (memory_mem_dm),                                               //                 .mem_dm
		.mem_dq                    (memory_mem_dq),                                               //                 .mem_dq
		.mem_dqs                   (memory_mem_dqs),                                              //                 .mem_dqs
		.mem_dqs_n                 (memory_mem_dqs_n),                                            //                 .mem_dqs_n
		.avl_ready                 (mm_interconnect_1_mem_if_lpddr2_emif_avl_waitrequest),        //              avl.waitrequest_n
		.avl_burstbegin            (mm_interconnect_1_mem_if_lpddr2_emif_avl_beginbursttransfer), //                 .beginbursttransfer
		.avl_addr                  (mm_interconnect_1_mem_if_lpddr2_emif_avl_address),            //                 .address
		.avl_rdata_valid           (mm_interconnect_1_mem_if_lpddr2_emif_avl_readdatavalid),      //                 .readdatavalid
		.avl_rdata                 (mm_interconnect_1_mem_if_lpddr2_emif_avl_readdata),           //                 .readdata
		.avl_wdata                 (mm_interconnect_1_mem_if_lpddr2_emif_avl_writedata),          //                 .writedata
		.avl_be                    (mm_interconnect_1_mem_if_lpddr2_emif_avl_byteenable),         //                 .byteenable
		.avl_read_req              (mm_interconnect_1_mem_if_lpddr2_emif_avl_read),               //                 .read
		.avl_write_req             (mm_interconnect_1_mem_if_lpddr2_emif_avl_write),              //                 .write
		.avl_size                  (mm_interconnect_1_mem_if_lpddr2_emif_avl_burstcount),         //                 .burstcount
		.local_init_done           (mem_if_lpddr2_emif_status_local_init_done),                   //           status.local_init_done
		.local_cal_success         (mem_if_lpddr2_emif_status_local_cal_success),                 //                 .local_cal_success
		.local_cal_fail            (mem_if_lpddr2_emif_status_local_cal_fail),                    //                 .local_cal_fail
		.oct_rzqin                 (oct_rzqin),                                                   //              oct.rzqin
		.pll_mem_clk               (),                                                            //      pll_sharing.pll_mem_clk
		.pll_write_clk             (),                                                            //                 .pll_write_clk
		.pll_locked                (),                                                            //                 .pll_locked
		.pll_write_clk_pre_phy_clk (),                                                            //                 .pll_write_clk_pre_phy_clk
		.pll_addr_cmd_clk          (),                                                            //                 .pll_addr_cmd_clk
		.pll_avl_clk               (),                                                            //                 .pll_avl_clk
		.pll_config_clk            (),                                                            //                 .pll_config_clk
		.pll_mem_phy_clk           (),                                                            //                 .pll_mem_phy_clk
		.afi_phy_clk               (),                                                            //                 .afi_phy_clk
		.pll_avl_phy_clk           ()                                                             //                 .pll_avl_phy_clk
	);

	D8M_QSYS_mipi_pwdn_n mipi_pwdn_n (
		.clk        (external_clk50_clk),                          //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_mipi_pwdn_n_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_mipi_pwdn_n_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_mipi_pwdn_n_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_mipi_pwdn_n_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_mipi_pwdn_n_s1_readdata),   //                    .readdata
		.out_port   (mipi_pwdn_n_external_connection_export)       // external_connection.export
	);

	D8M_QSYS_mipi_pwdn_n mipi_reset_n (
		.clk        (external_clk50_clk),                           //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_mipi_reset_n_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_mipi_reset_n_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_mipi_reset_n_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_mipi_reset_n_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_mipi_reset_n_s1_readdata),   //                    .readdata
		.out_port   (mipi_reset_n_external_connection_export)       // external_connection.export
	);

	D8M_QSYS_nios2_qsys nios2_qsys (
		.clk                                   (external_clk50_clk),                                         //                       clk.clk
		.reset_n                               (~rst_controller_002_reset_out_reset),                        //                   reset_n.reset_n
		.reset_req                             (rst_controller_002_reset_out_reset_req),                     //                          .reset_req
		.d_address                             (nios2_qsys_data_master_address),                             //               data_master.address
		.d_byteenable                          (nios2_qsys_data_master_byteenable),                          //                          .byteenable
		.d_read                                (nios2_qsys_data_master_read),                                //                          .read
		.d_readdata                            (nios2_qsys_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (nios2_qsys_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (nios2_qsys_data_master_write),                               //                          .write
		.d_writedata                           (nios2_qsys_data_master_writedata),                           //                          .writedata
		.d_readdatavalid                       (nios2_qsys_data_master_readdatavalid),                       //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (nios2_qsys_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (nios2_qsys_instruction_master_address),                      //        instruction_master.address
		.i_read                                (nios2_qsys_instruction_master_read),                         //                          .read
		.i_readdata                            (nios2_qsys_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (nios2_qsys_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (nios2_qsys_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (nios2_qsys_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_qsys_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_nios2_qsys_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_nios2_qsys_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_nios2_qsys_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_nios2_qsys_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_nios2_qsys_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_nios2_qsys_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_nios2_qsys_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_nios2_qsys_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                            // custom_instruction_master.readra
	);

	D8M_QSYS_onchip_memory2 onchip_memory2 (
		.clk        (external_clk50_clk),                             //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),             // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req)          //       .reset_req
	);

	D8M_QSYS_sysid_qsys sysid_qsys (
		.clock    (external_clk50_clk),                                  //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                 //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_control_slave_address)   //              .address
	);

	D8M_QSYS_timer timer (
		.clk        (external_clk50_clk),                    //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),   // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)               //   irq.irq
	);

	D8M_QSYS_mm_interconnect_0 mm_interconnect_0 (
		.clk_50_clk_clk                                         (external_clk50_clk),                                                 //                                       clk_50_clk.clk
		.mem_if_lpddr2_emif_afi_clk_clk                         (mem_if_lpddr2_emif_afi_clk_clk),                                     //                       mem_if_lpddr2_emif_afi_clk.clk
		.jtag_uart_reset_reset_bridge_in_reset_reset            (rst_controller_001_reset_out_reset),                                 //            jtag_uart_reset_reset_bridge_in_reset.reset
		.nios2_qsys_reset_n_reset_bridge_in_reset_reset         (rst_controller_002_reset_out_reset),                                 //         nios2_qsys_reset_n_reset_bridge_in_reset.reset
		.TERASIC_AUTO_FOCUS_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                     // TERASIC_AUTO_FOCUS_0_reset_reset_bridge_in_reset.reset
		.nios2_qsys_data_master_address                         (nios2_qsys_data_master_address),                                     //                           nios2_qsys_data_master.address
		.nios2_qsys_data_master_waitrequest                     (nios2_qsys_data_master_waitrequest),                                 //                                                 .waitrequest
		.nios2_qsys_data_master_byteenable                      (nios2_qsys_data_master_byteenable),                                  //                                                 .byteenable
		.nios2_qsys_data_master_read                            (nios2_qsys_data_master_read),                                        //                                                 .read
		.nios2_qsys_data_master_readdata                        (nios2_qsys_data_master_readdata),                                    //                                                 .readdata
		.nios2_qsys_data_master_readdatavalid                   (nios2_qsys_data_master_readdatavalid),                               //                                                 .readdatavalid
		.nios2_qsys_data_master_write                           (nios2_qsys_data_master_write),                                       //                                                 .write
		.nios2_qsys_data_master_writedata                       (nios2_qsys_data_master_writedata),                                   //                                                 .writedata
		.nios2_qsys_data_master_debugaccess                     (nios2_qsys_data_master_debugaccess),                                 //                                                 .debugaccess
		.nios2_qsys_instruction_master_address                  (nios2_qsys_instruction_master_address),                              //                    nios2_qsys_instruction_master.address
		.nios2_qsys_instruction_master_waitrequest              (nios2_qsys_instruction_master_waitrequest),                          //                                                 .waitrequest
		.nios2_qsys_instruction_master_read                     (nios2_qsys_instruction_master_read),                                 //                                                 .read
		.nios2_qsys_instruction_master_readdata                 (nios2_qsys_instruction_master_readdata),                             //                                                 .readdata
		.nios2_qsys_instruction_master_readdatavalid            (nios2_qsys_instruction_master_readdatavalid),                        //                                                 .readdatavalid
		.hdmi_tx_int_n_s1_address                               (mm_interconnect_0_hdmi_tx_int_n_s1_address),                         //                                 hdmi_tx_int_n_s1.address
		.hdmi_tx_int_n_s1_write                                 (mm_interconnect_0_hdmi_tx_int_n_s1_write),                           //                                                 .write
		.hdmi_tx_int_n_s1_readdata                              (mm_interconnect_0_hdmi_tx_int_n_s1_readdata),                        //                                                 .readdata
		.hdmi_tx_int_n_s1_writedata                             (mm_interconnect_0_hdmi_tx_int_n_s1_writedata),                       //                                                 .writedata
		.hdmi_tx_int_n_s1_chipselect                            (mm_interconnect_0_hdmi_tx_int_n_s1_chipselect),                      //                                                 .chipselect
		.i2c_opencores_camera_avalon_slave_0_address            (mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_address),      //              i2c_opencores_camera_avalon_slave_0.address
		.i2c_opencores_camera_avalon_slave_0_write              (mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_write),        //                                                 .write
		.i2c_opencores_camera_avalon_slave_0_readdata           (mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_readdata),     //                                                 .readdata
		.i2c_opencores_camera_avalon_slave_0_writedata          (mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_writedata),    //                                                 .writedata
		.i2c_opencores_camera_avalon_slave_0_waitrequest        (~mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_waitrequest), //                                                 .waitrequest
		.i2c_opencores_camera_avalon_slave_0_chipselect         (mm_interconnect_0_i2c_opencores_camera_avalon_slave_0_chipselect),   //                                                 .chipselect
		.i2c_opencores_mipi_avalon_slave_0_address              (mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_address),        //                i2c_opencores_mipi_avalon_slave_0.address
		.i2c_opencores_mipi_avalon_slave_0_write                (mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_write),          //                                                 .write
		.i2c_opencores_mipi_avalon_slave_0_readdata             (mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_readdata),       //                                                 .readdata
		.i2c_opencores_mipi_avalon_slave_0_writedata            (mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_writedata),      //                                                 .writedata
		.i2c_opencores_mipi_avalon_slave_0_waitrequest          (~mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_waitrequest),   //                                                 .waitrequest
		.i2c_opencores_mipi_avalon_slave_0_chipselect           (mm_interconnect_0_i2c_opencores_mipi_avalon_slave_0_chipselect),     //                                                 .chipselect
		.i2c_scl_s1_address                                     (mm_interconnect_0_i2c_scl_s1_address),                               //                                       i2c_scl_s1.address
		.i2c_scl_s1_write                                       (mm_interconnect_0_i2c_scl_s1_write),                                 //                                                 .write
		.i2c_scl_s1_readdata                                    (mm_interconnect_0_i2c_scl_s1_readdata),                              //                                                 .readdata
		.i2c_scl_s1_writedata                                   (mm_interconnect_0_i2c_scl_s1_writedata),                             //                                                 .writedata
		.i2c_scl_s1_chipselect                                  (mm_interconnect_0_i2c_scl_s1_chipselect),                            //                                                 .chipselect
		.i2c_sda_s1_address                                     (mm_interconnect_0_i2c_sda_s1_address),                               //                                       i2c_sda_s1.address
		.i2c_sda_s1_write                                       (mm_interconnect_0_i2c_sda_s1_write),                                 //                                                 .write
		.i2c_sda_s1_readdata                                    (mm_interconnect_0_i2c_sda_s1_readdata),                              //                                                 .readdata
		.i2c_sda_s1_writedata                                   (mm_interconnect_0_i2c_sda_s1_writedata),                             //                                                 .writedata
		.i2c_sda_s1_chipselect                                  (mm_interconnect_0_i2c_sda_s1_chipselect),                            //                                                 .chipselect
		.jtag_uart_avalon_jtag_slave_address                    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),              //                      jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),                //                                                 .write
		.jtag_uart_avalon_jtag_slave_read                       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),                 //                                                 .read
		.jtag_uart_avalon_jtag_slave_readdata                   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),             //                                                 .readdata
		.jtag_uart_avalon_jtag_slave_writedata                  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),            //                                                 .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),          //                                                 .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                 (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),           //                                                 .chipselect
		.key_s1_address                                         (mm_interconnect_0_key_s1_address),                                   //                                           key_s1.address
		.key_s1_readdata                                        (mm_interconnect_0_key_s1_readdata),                                  //                                                 .readdata
		.mipi_pwdn_n_s1_address                                 (mm_interconnect_0_mipi_pwdn_n_s1_address),                           //                                   mipi_pwdn_n_s1.address
		.mipi_pwdn_n_s1_write                                   (mm_interconnect_0_mipi_pwdn_n_s1_write),                             //                                                 .write
		.mipi_pwdn_n_s1_readdata                                (mm_interconnect_0_mipi_pwdn_n_s1_readdata),                          //                                                 .readdata
		.mipi_pwdn_n_s1_writedata                               (mm_interconnect_0_mipi_pwdn_n_s1_writedata),                         //                                                 .writedata
		.mipi_pwdn_n_s1_chipselect                              (mm_interconnect_0_mipi_pwdn_n_s1_chipselect),                        //                                                 .chipselect
		.mipi_reset_n_s1_address                                (mm_interconnect_0_mipi_reset_n_s1_address),                          //                                  mipi_reset_n_s1.address
		.mipi_reset_n_s1_write                                  (mm_interconnect_0_mipi_reset_n_s1_write),                            //                                                 .write
		.mipi_reset_n_s1_readdata                               (mm_interconnect_0_mipi_reset_n_s1_readdata),                         //                                                 .readdata
		.mipi_reset_n_s1_writedata                              (mm_interconnect_0_mipi_reset_n_s1_writedata),                        //                                                 .writedata
		.mipi_reset_n_s1_chipselect                             (mm_interconnect_0_mipi_reset_n_s1_chipselect),                       //                                                 .chipselect
		.nios2_qsys_jtag_debug_module_address                   (mm_interconnect_0_nios2_qsys_jtag_debug_module_address),             //                     nios2_qsys_jtag_debug_module.address
		.nios2_qsys_jtag_debug_module_write                     (mm_interconnect_0_nios2_qsys_jtag_debug_module_write),               //                                                 .write
		.nios2_qsys_jtag_debug_module_read                      (mm_interconnect_0_nios2_qsys_jtag_debug_module_read),                //                                                 .read
		.nios2_qsys_jtag_debug_module_readdata                  (mm_interconnect_0_nios2_qsys_jtag_debug_module_readdata),            //                                                 .readdata
		.nios2_qsys_jtag_debug_module_writedata                 (mm_interconnect_0_nios2_qsys_jtag_debug_module_writedata),           //                                                 .writedata
		.nios2_qsys_jtag_debug_module_byteenable                (mm_interconnect_0_nios2_qsys_jtag_debug_module_byteenable),          //                                                 .byteenable
		.nios2_qsys_jtag_debug_module_waitrequest               (mm_interconnect_0_nios2_qsys_jtag_debug_module_waitrequest),         //                                                 .waitrequest
		.nios2_qsys_jtag_debug_module_debugaccess               (mm_interconnect_0_nios2_qsys_jtag_debug_module_debugaccess),         //                                                 .debugaccess
		.onchip_memory2_s1_address                              (mm_interconnect_0_onchip_memory2_s1_address),                        //                                onchip_memory2_s1.address
		.onchip_memory2_s1_write                                (mm_interconnect_0_onchip_memory2_s1_write),                          //                                                 .write
		.onchip_memory2_s1_readdata                             (mm_interconnect_0_onchip_memory2_s1_readdata),                       //                                                 .readdata
		.onchip_memory2_s1_writedata                            (mm_interconnect_0_onchip_memory2_s1_writedata),                      //                                                 .writedata
		.onchip_memory2_s1_byteenable                           (mm_interconnect_0_onchip_memory2_s1_byteenable),                     //                                                 .byteenable
		.onchip_memory2_s1_chipselect                           (mm_interconnect_0_onchip_memory2_s1_chipselect),                     //                                                 .chipselect
		.onchip_memory2_s1_clken                                (mm_interconnect_0_onchip_memory2_s1_clken),                          //                                                 .clken
		.sysid_qsys_control_slave_address                       (mm_interconnect_0_sysid_qsys_control_slave_address),                 //                         sysid_qsys_control_slave.address
		.sysid_qsys_control_slave_readdata                      (mm_interconnect_0_sysid_qsys_control_slave_readdata),                //                                                 .readdata
		.TERASIC_AUTO_FOCUS_0_mm_ctrl_address                   (mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_address),             //                     TERASIC_AUTO_FOCUS_0_mm_ctrl.address
		.TERASIC_AUTO_FOCUS_0_mm_ctrl_write                     (mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_write),               //                                                 .write
		.TERASIC_AUTO_FOCUS_0_mm_ctrl_read                      (mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_read),                //                                                 .read
		.TERASIC_AUTO_FOCUS_0_mm_ctrl_readdata                  (mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_readdata),            //                                                 .readdata
		.TERASIC_AUTO_FOCUS_0_mm_ctrl_writedata                 (mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_writedata),           //                                                 .writedata
		.TERASIC_AUTO_FOCUS_0_mm_ctrl_chipselect                (mm_interconnect_0_terasic_auto_focus_0_mm_ctrl_chipselect),          //                                                 .chipselect
		.timer_s1_address                                       (mm_interconnect_0_timer_s1_address),                                 //                                         timer_s1.address
		.timer_s1_write                                         (mm_interconnect_0_timer_s1_write),                                   //                                                 .write
		.timer_s1_readdata                                      (mm_interconnect_0_timer_s1_readdata),                                //                                                 .readdata
		.timer_s1_writedata                                     (mm_interconnect_0_timer_s1_writedata),                               //                                                 .writedata
		.timer_s1_chipselect                                    (mm_interconnect_0_timer_s1_chipselect)                               //                                                 .chipselect
	);

	D8M_QSYS_mm_interconnect_1 mm_interconnect_1 (
		.mem_if_lpddr2_emif_afi_clk_clk                            (mem_if_lpddr2_emif_afi_clk_clk),                              //                          mem_if_lpddr2_emif_afi_clk.clk
		.alt_vip_vfb_0_reset_reset_bridge_in_reset_reset           (rst_controller_reset_out_reset),                              //           alt_vip_vfb_0_reset_reset_bridge_in_reset.reset
		.mem_if_lpddr2_emif_soft_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                              // mem_if_lpddr2_emif_soft_reset_reset_bridge_in_reset.reset
		.alt_vip_vfb_0_read_master_address                         (alt_vip_vfb_0_read_master_address),                           //                           alt_vip_vfb_0_read_master.address
		.alt_vip_vfb_0_read_master_waitrequest                     (alt_vip_vfb_0_read_master_waitrequest),                       //                                                    .waitrequest
		.alt_vip_vfb_0_read_master_burstcount                      (alt_vip_vfb_0_read_master_burstcount),                        //                                                    .burstcount
		.alt_vip_vfb_0_read_master_read                            (alt_vip_vfb_0_read_master_read),                              //                                                    .read
		.alt_vip_vfb_0_read_master_readdata                        (alt_vip_vfb_0_read_master_readdata),                          //                                                    .readdata
		.alt_vip_vfb_0_read_master_readdatavalid                   (alt_vip_vfb_0_read_master_readdatavalid),                     //                                                    .readdatavalid
		.alt_vip_vfb_0_write_master_address                        (alt_vip_vfb_0_write_master_address),                          //                          alt_vip_vfb_0_write_master.address
		.alt_vip_vfb_0_write_master_waitrequest                    (alt_vip_vfb_0_write_master_waitrequest),                      //                                                    .waitrequest
		.alt_vip_vfb_0_write_master_burstcount                     (alt_vip_vfb_0_write_master_burstcount),                       //                                                    .burstcount
		.alt_vip_vfb_0_write_master_write                          (alt_vip_vfb_0_write_master_write),                            //                                                    .write
		.alt_vip_vfb_0_write_master_writedata                      (alt_vip_vfb_0_write_master_writedata),                        //                                                    .writedata
		.mem_if_lpddr2_emif_avl_address                            (mm_interconnect_1_mem_if_lpddr2_emif_avl_address),            //                              mem_if_lpddr2_emif_avl.address
		.mem_if_lpddr2_emif_avl_write                              (mm_interconnect_1_mem_if_lpddr2_emif_avl_write),              //                                                    .write
		.mem_if_lpddr2_emif_avl_read                               (mm_interconnect_1_mem_if_lpddr2_emif_avl_read),               //                                                    .read
		.mem_if_lpddr2_emif_avl_readdata                           (mm_interconnect_1_mem_if_lpddr2_emif_avl_readdata),           //                                                    .readdata
		.mem_if_lpddr2_emif_avl_writedata                          (mm_interconnect_1_mem_if_lpddr2_emif_avl_writedata),          //                                                    .writedata
		.mem_if_lpddr2_emif_avl_beginbursttransfer                 (mm_interconnect_1_mem_if_lpddr2_emif_avl_beginbursttransfer), //                                                    .beginbursttransfer
		.mem_if_lpddr2_emif_avl_burstcount                         (mm_interconnect_1_mem_if_lpddr2_emif_avl_burstcount),         //                                                    .burstcount
		.mem_if_lpddr2_emif_avl_byteenable                         (mm_interconnect_1_mem_if_lpddr2_emif_avl_byteenable),         //                                                    .byteenable
		.mem_if_lpddr2_emif_avl_readdatavalid                      (mm_interconnect_1_mem_if_lpddr2_emif_avl_readdatavalid),      //                                                    .readdatavalid
		.mem_if_lpddr2_emif_avl_waitrequest                        (~mm_interconnect_1_mem_if_lpddr2_emif_avl_waitrequest)        //                                                    .waitrequest
	);

	D8M_QSYS_irq_mapper irq_mapper (
		.clk           (external_clk50_clk),                 //       clk.clk
		.reset         (rst_controller_002_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),           // receiver4.irq
		.sender_irq    (nios2_qsys_d_irq_irq)                //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~external_reset_reset_n),        // reset_in0.reset
		.clk            (mem_if_lpddr2_emif_afi_clk_clk), //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~external_reset_reset_n),                // reset_in0.reset
		.clk            (external_clk50_clk),                     //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~external_reset_reset_n),                  // reset_in0.reset
		.reset_in1      (nios2_qsys_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (external_clk50_clk),                       //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),       // reset_out.reset
		.reset_req      (rst_controller_002_reset_out_reset_req),   //          .reset_req
		.reset_req_in0  (1'b0),                                     // (terminated)
		.reset_req_in1  (1'b0),                                     // (terminated)
		.reset_in2      (1'b0),                                     // (terminated)
		.reset_req_in2  (1'b0),                                     // (terminated)
		.reset_in3      (1'b0),                                     // (terminated)
		.reset_req_in3  (1'b0),                                     // (terminated)
		.reset_in4      (1'b0),                                     // (terminated)
		.reset_req_in4  (1'b0),                                     // (terminated)
		.reset_in5      (1'b0),                                     // (terminated)
		.reset_req_in5  (1'b0),                                     // (terminated)
		.reset_in6      (1'b0),                                     // (terminated)
		.reset_req_in6  (1'b0),                                     // (terminated)
		.reset_in7      (1'b0),                                     // (terminated)
		.reset_req_in7  (1'b0),                                     // (terminated)
		.reset_in8      (1'b0),                                     // (terminated)
		.reset_req_in8  (1'b0),                                     // (terminated)
		.reset_in9      (1'b0),                                     // (terminated)
		.reset_req_in9  (1'b0),                                     // (terminated)
		.reset_in10     (1'b0),                                     // (terminated)
		.reset_req_in10 (1'b0),                                     // (terminated)
		.reset_in11     (1'b0),                                     // (terminated)
		.reset_req_in11 (1'b0),                                     // (terminated)
		.reset_in12     (1'b0),                                     // (terminated)
		.reset_req_in12 (1'b0),                                     // (terminated)
		.reset_in13     (1'b0),                                     // (terminated)
		.reset_req_in13 (1'b0),                                     // (terminated)
		.reset_in14     (1'b0),                                     // (terminated)
		.reset_req_in14 (1'b0),                                     // (terminated)
		.reset_in15     (1'b0),                                     // (terminated)
		.reset_req_in15 (1'b0)                                      // (terminated)
	);

endmodule
