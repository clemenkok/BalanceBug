��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�!��
��%Y l�׾����|R�bD�E���y"���7�c�t#�l��I�k����;�6�����M�^�v���A�ko�aB��mMe�S�?U�{�S!=B����[[؊�W��5,�ɮ�-�g��Ok�w��1CieS�:hB��a����i���D�ٮK���zm"~<�E=�ܣB�r|��2��L^A��/���󥿛�9F�r��:٩m�}�I�C����F��ofSN����=,�s��|�M�?���E�+���d4�/1��&�tz�TА���}8=���)�*�i8M�[���i�ƵjhI���M7V<�<��S��r�d����_]D)�["\��2��E�&"��w���z�}s!��"��8'*a���J�tY�g,}���Y-y�@��FU%�ropW�.'�7{��+�-T�UV�F�>�?��,˅�L���VKmw�i�b���Ԥ�����q�йXu�f�%Wt7�H��x�kwbJ�o���������~-F4^L�!t2�#�������<�s�R�U�� @�m�?�Fft?>]eq�A7XH� Cq��k+���Ԓ���񅳢lM@\I�D;<8O����7q`/pyQ&�3b"�Q��z�w
�eS�$6�'�����ce|���O��3��#�f��SlK�@ϱ*0��*�]�*7�y�S�/鸘��p�'��e7ؖ�3�2�����"I�Čm/2�`�"��5�	�[#��+)|�G��G8��5���N�� �p���5]�eU�,�	�i��KӘ���vuɋ �I�>g�0A����Up��ʘ9�O6Qӛ��ia{bi�M�9�e	u���Eq?�d����ݚ�׮�=�i�Og^�Q7���^��{��Z�'z��$Hm<	�4:��51U�o���F`{H�������$jK���#y؈2D�&�2�7�1`(jl�2�i-iD��}w�'$#�A�8;u2',.MRH;8�B{��m�G����K��@\N}B<J©$�6�H��Kd�w�̕h6�U<��X��`�ɉ��Rꣷ�2\����^,.�4�VoC��7J�R[%l*�ps^�Tɩ�iZ[A��ӷ�Z���{�;�u��G����7��PO0K����_~�*���>!ח�E�����:�+��Y�"D�¯G��U��ʑ�,p�"������j짾�E�]z�qsuM��g��C6�/���2e��u)�#͔Y�������S�k��~1\��U��h�r���TT��?�rx��~��E_�������Z3�i�{��(v�{��w�\�(�@�e�Ñ������Q����+.(��ʹ�̷�}��e�Zyf������h$��X��<�l�)����k�~��M2���7�(U�^�e5�`�H5Bç�I#�X�|�:m�C�*����s~�����n�%Ww�h���Ƴ�EEz����Xi��a��Ն2�Qr�m?�z�áikWD��k�B�5��:�4�}�Qݔ?��de�5��k���\�J�2R�G�*�W8E~���#���"�VI���b�.-\>x.Xև���2$C��I%��r�]��,�1e,_���������>�Q�Cif6{�9����}��`=«�V��m���|���9f�o��$BSl���g ^)*K��y��^�b@���D��|��ES�bx4����[`� ��4b��s�-W1��sܫ��a���cCT`c�}�п|���ҧL�H�೔�#C�?M�w�x�.�nzI�_���D翸SN�����o$[�;�ҡ�����j@�?S���n�W�h��eZ�%)���J�X4,y$.�F�5� ?�_Q�c���r)lb�z�T ������'!_1��l~&_񻞦�~����+��#�Rc(�B��w�n�N�q!!�5^gV#2a������7�K�U�!�R�Q�L�!�x�EZ,[�y,Z6�YU˂���t*�?�OX����f=������dnB��+���P��9�B�p�)<|���u,I�n�	[t�$_�[����&�"xW̽��_I�<'���cs�}�6�ͩ��R����匽K�f6tĠ�P��\0���_�OM�h�&"H.�0s������.��^��\Z�iM������)�v��"�1��1 R�P��n����Q��{��=�״������f�[v��s�����,6�ʋj�if����Bj���J�C�=+M�U�
��۽��^�m5��b]#N�t\p��\Z��Σ�H�����8E�gd-#4,%����96���:��c�-wlY��԰G��U�;.�㍟�oUq��j0ʃ����A��n[����Y��p�,���\mq�uI��ov!W�1�"(r��W����o9�%������l�M�|�� /�rt�e��/�&FI~�����!7���`H�~"���p����QP!��;Y4^yY���
xsR��ffNht,�!�no�W�C)'�a;Q�:�6l���yͳ�i��₍�)�X��J��2(񹟌��<o��6�-G�_�*��J)��46O��=Ì8M�1h�����'Ɂ��&��@*�� ��'�bڕp9$x	܌�y��)�c����2��Y>{I�8ήb����)q�I4�=�[C��K`2j^9������������S�Z�"ퟯ�̱�M; 2�5C��dx� (�c��.�.`�,��1��7Pq��\%��&T��)AHc�h{5��72�yW��݈�ȩt��NQ+��4\��Mܟ��F[�Ti�O{@
���q8�^�L�}�j����D�V�hg�땸*�o%����V��}�2�՟fN��e�\��č�,e�JS8��SH	K�o:k�rc�ʶq�u������RM|Nfxc������S���k��x����>��`��\T����W6���U�Y��I�e0}�3��B���_p~�M�\4��u�WJ�:�"3):-AH�R�n(�
MtQ�����,���tQ!�����!Y�!O
����.��TE��:��-~'7&�*^�y������J�����Ϋ�:�`H��d�O���/�\�k�M>��kȡ82aQ���-��i�O�������?Ec~g��=�L0^؀8^���k�CΔ#��{�u�f;<�3�.(�7�s���b���۔���Ǽ�ZP�7�f�Č{;���Û��9�z��	O)��`&e��g���j�'�b:~C�:�$������6Z8����y�~��QI�@� �8SjBNc~=��?��Hޙ"]�|��[9`m��O�t�vpj��j,6=�
E��Ig���M<��T6�k�+�lL	n�� �!k���Sه�YBoJ�O�j};xa����6��������1Bg6�T:�M`Mo�`s���X��<�?����x���eQpVef�ȷ(�۱�dL�0���
l��K$�j�z�ԃ^��t
9��;ڝ]c|��=��6�3Z�F��2Bp^r�%���b���r� 6~�o�C�a�*�77�_Ch�w��%I�H۠�X;B�������t�Q�H�J�y��f/�7�^Dw�OW!\L�7���*x�F$~�3@��X���rq���/����
�ʸB�E�k5��k�$�H��<֣����p$7{�K&�S��b,�G޽�޶�"U�ib����3؏��e� ��O��Xe�m�[�Q�oRj{x�+�"F *=���1]p�`9�'��e �([�>S\����[��]ݾ�߇Aدv!��{�q��T2ϑ϶+a�?�E�pa:����jt���ʹ�t�b8�kT�����*�$N�
V&��e��d%T�C���a�>�9�kC�'�c\Z���=�"Dt�U=���n.=��B)����b'�/x�T�[Xv��m�#3��R���3]ڑ�p>�3'�[�>�d�=�����[�OC�Tq�v���=��ٔ���"⠓g'O�br-�[;��> �Z���O�&⺛��|����<	�g�����A�t�/l0��Q�w���[�����:�PG��@����a� �m�G:+H��N�D ԣXa���8p+�ļJCC��pl��DO�������o�!X�����_�1
!�ꭅV���^+"�\J����]3�����8�\�xӾɍ)<3��s��3�x�{AA�8�+2��'�WZ�#jVpU��ږ��5r[�� +"��S\���S�5JJ`�p��s�!g��gu�T����{g^�}!t��36�^"�Y(�P��}�`E^��5�Yö���|B"[��^;9����v4D���]7S��wi.ؚ��OS�y��2H�����s���'ž"�2�1�h�}8���a�]v(�^i�����?v�w��9�� ]i{�{04L�N�fD�;B�K��ˏE(,�n�r�r�\�� n�Xg�H�������px�e1�� ���t���&��]��������a�Ch�G��<�ۅ,�p�.�`}�>5K��6hd�*���@�7	��i᯴~�₰��q�vUI�ʬ�`^�Q'+��m��a���� �e轲�%���ʄU"5��@�ۤ�ԫ���~8��eR������R'=� �q�Ē1�CFV�ADf=��!�Sϊ��Xƻ�����Ϸ5��X�l7�UdwpF��%��f,-]ݔ����mk[I�����{��F�K�@�~�|�ږl0B}�<M�`����`��������bQ7C��7��b��|5_!��Bh�v[��h;�V_��#�����5�A��O}�-L�o�6�1��\���oe4�Q����{���p#c�����T�L����#b:������a>������(�E�>�kx�S���b�H�h���&�1����)�b�	�����!\X�"̡�jϜc�Ӡ���<�R%߶�k��g�ds�������4�P����tlG#� c��&Y���r c�ɢFK�aD�bd��3��>��lƺda{�o%��?����T�0�M��mn��I��vYG�6r��h�F�$�-��@@I���[���A�%Z�L���6����(�Y9�m�mlU�+ S��V�m>���������w�i���'����ൿ�1�,D�ߴ&���N��U�ˎ���V�o |�P���k�-�ZW��U�L���6	X�\�7�4K���<�lmX	+G^F5�wG�I>��I�f� �
�w� 4�C�;~����tX��Z��{`n�u��7��5��?(��B�����~�r7��H+'�(݉R3��@��Y�G���N��i�Uµ^K´� g�;T�� �6�@�[��t���{�IЌ���/���A�!���uA�Ф�������Qܷ���+��d�Dm9�b�Uc�]F4�2�d�#���sYHZ���4�r��~����_a^��:�4�w��9Ku���p��+����	�azfJT]_��{�z�5�&D7^	&�`�A�Y�O�U�c��l �&|˄���Ǜ��x�3����`�Ml�s��&�p{�4F0����i۽�mZ�,7eꄷR	R� �y0����46yEL��.�PY��B�<eP�;���"M[4&[������:� >�+��1�����7�S�t��@����Vk�i)���M�j_��P��N�!���n7������&gÀ�c���*��mlE���M�A����w��3^f��Nտ7�Eg[��x�0�^�.�ڧ�q�z!�#��?�A_:��N����ض�h�ɠ� h�ˮ�`��o6kP�&go���(��E>(����t��<�y��n�ֹ3P&�e�����$ɑ�/�?�?h�qj3W�g���B*��^���t���P+R����`�XE-��f�Ž!E��7<�RH�sq��{��fCr��^�����X�\9b�r���@{��gǄ+�즐�3��+���U+*�xW��|�I��`Wd-$�]����S���fTMo���f�$,�p�X�3|:=Z����2>C=����&:1i�)4�d��@Gh���Y����Cq��nq���#�3��@&�f��.�$랳(w,��FEw�F��Ћ�b[j�� _U�G�5Y�\!ĺ>���"��55T}	�L�B�z����nuCSP���Y�y�/ ��L��k~j��7�=�����9Z!�c�1Z�vb/��q]�#�+���^�fAyQ\��ӛ��T���$��[��)ɐ�_Ih�4X������;�rA��C�����_3/�&���{�~>Qj��T�5%o{����T���6��0��i���*'�������=��;�6�6?�kco-V�с]0T6I@+� ���� ��WM��o��'��,�d��es%�7��i�&�r�2�	ߒ�����:ä�HR��Tn�G�o���k�@��F�����H�"��P���g�@�
��* ��ꋶm]-k������[��lB��.��f����&~>Q����3jvB��+p�$TQ�"�ܲ.�p���W!����b�DG��ϮщL�V�k��I�Q�N�D����{{�^�d���L!B�hН��%n.����.����Ag������X��_�-��'i�ԭR\�*u��9����\�2��1O-L��J@� &�j��ס����ىk��S�l�|l��-Jz|�����ـ?b[/��ӰTTt�3V�����B�䳥�Hϣl�Qg�%5PF��I1��M�N%W$T�f�WLw�(Sk�J�?Z����qe�O�_�"����3�ƃ���]�d�K\fK�6q�� O1B�� OaHi��Wi0"hV��J!@m;d��<�[�e�j�f����*f�Y2�A��X���  �{�]�j��dPs�CÛ�7-���6A�r�E��ԒuYݗ:���,�����o֖(���������E9��v"wTF�=_-	λHqv�cu��ĴK�O�}o���D@``�Q{1N�s�f1=h���?ۘ�'&�Ǹh��P/����4u���kzG]���`�'����T,y&����[}��Q�-���ߤ�(����[�b�vԶ�$��-�2�O�y�[x|F�74�Q�}R<P��5��u)�y��#�P���.��=~2��OW��:�Y{'��o��2���V�s�w!��5X�@E�R�<R�3R����7B��ɋ���[3��Ty=ʲ��5{�?WN�ԭ�(�?YȐ:�	�Ϻ/����k���!fU�F���mg�,!@��O�y�_k/�x��z��M��9����(Hm�����8�(Uaw'�*���,��X���c�KR�@�w�e>yU1� ��؏�jz��-zͺa���D�\���e�u�2T������Bص
,�=j���<p�ʵ	��.n�}��6Y�SBc7"`>�PɀZ�D�������-|�4�`|��:L7�I/vo�������Λ�c����̌�g�W=�0�X	�Ŝ��ަ槺������cE` �� �;4ϙ��c-���ݿ�'�7�Ne
=C���!�g t#�Z&�t�r�V�G;[�jR/,���jO �XO�o���^��ح�w�XO=�*��b'o��c�I��6��`�*�êPo��vhsZk[iC��W�Mp@��o���`�YJ��TIP::ӡ�<��jN���b�~�"��)���Ob4��!Й�����=E�e�7HP�YS!@5��}����F$˙��e౾0rjFjV3�c1�rck VS�3X���0,����hc��tz#�]�.��+��UJ��(c��\��q��S���ן-l�='��i :�:f����c�t�RB�"�~R~H���}��g��1<X�a��^���u�p\��]\��2'��{k�)t�.����
J=�X��i�4��p%p�>�����!l8D�@/�덈�98����%�L�!d��x�%3ܺ��t�=40�[�<����5��7e9� '\�S�TR�=��d)rf�
���$�㞔�Pg��+az����S��̉�]�H-�c�'���ܮP����w��,b�c,��!�c��/��Ro�h`${�NN��O��1�2i`
`�jI�]��7�SΎ:_4S�I�T��j;�U�Qme�h�����Fߗ�ҧ�u��,�< A�R�@�����)\vxz�}hp3��ևzf	3?���w�F+?O�8a�ff�E���F�{��p\&ٻ#�s���j���p�tӖm!KW��!�j����.A(Y�N�)OSv�%���[w�sN���F��8,�Xq��N�S��Ҿ�i$��ay���j�5:��c=n%܁�l>�u�Ѩ|M.8g�v���yb�Q?���R���U�dX��s��ez��s]m��jMv���*��c��X�ҷX�꜕:�|[���mfWx�>�8�T!�ѻi�a=j\�c��M�����mnZ�����O)ߦm��V������˻Mtqʟ��Z���l�P��s�?��}ʉ��c�"(����,o�
�G��,I�\�-1fg�Ğ>N{�ܲ@�0���F���/��!/ {µ�	Vu�9Ь�^��s�q���P���`��q2�]8�d�G;F�)�!E�p'y����a�v�+,S�����2��=��Ix=k1��'�+ݩ��Q��Zp��n��Rtb҈�Lt(���|�U	�.���eĩǙ�0����twkv�o�t	���8+�ÄD����|}ʹ�^�Ûe����
L�U�X�֩��	�55����Jc��G	�f}�C�n`��Y�M�@�c�����G��Y�^|_,E�Ȋ�-�]my�WU��9�E���:��q{g��ul�-��Pd�����#7օ��U�_��'��v)D�H�ûϔ�֙�s����n!�XBj�'�B:����S�Mm$x�ummN0D^f�S��ё�R��Zۧ#Gޱ�Cm�������P��F1���#��=V|h�c?^=1Qo%՘z7+�s�������_E-Y�����o���%n9\dP��?��\��a�>�:Һy���_~&�ľ�嶅��Pa�^�l󝍮�@ĕl�j@,�1��N��P��Y�:�H}'�3C��t"W���ZKv���^TCy��m��˞�&�L��E�*]p�~����pC�]^�הo�����}:$YՏ"BKP�ӲĈye�v�<}[��mYS�4��ec���8(�Ѐ�(Z
��G��T�g/i��$e�k�����ԷD��2F �3u	2ȕ��+X�Ta��eGt2#z/�Π����ʨ<�׍:h�muo;�$�,���	�~¨���Oy����i`+��=)��a�@�o\d�;�.nP�����\��I���D~y�IcƂ�a ��d��`P�LF!1Mj��U�@hj����'�-�6<�g���=�^�� ��a��J4:��%N���8d�,�0(Hűg�&��男x_D��S&�����m����ec#G=Fw�#
�ҹ��c�@5&- +�ߋ%f��~x؞�&K�Z-xC�"�������`RM$%�Yȑ_b��2���]�x�x}���?}����#p����.s�BY���;BA�r

H�Mҁb�A�n@�)*����h�Jaݔ�״��%>�����E2�[��c@�lr��yS�E������L� ?c;~(Vrj����T�z/�.C����}`#����W�G�w�E�O|�R��J��Y@`B��U9+�w��$��r��pkF�,���X�4���+Q�?����䧌��v�>G���e9
���^#���Q���!m�X�}��>��^�m�+��E��5�qs Q}Hd�#WX����#��V�~�`�4ٔT5	��^�s$Zg�TR�<ϒ/���,#hϾ��3�uy^�E�-�=�0�Ri��f�����>�����5��{��Wqyv����Q�y�q�@h7����;��Z�w��X��67��� ߪ�?\�j=�)vF���9��	}B��Fy�%���7G�5��˜:��Pa�m�!J����2����X%�a�֙���T����Wk�F��H�\����6�td�!���[�=1�i���v'V���?�*�u{�5?���6��`4��3�K�"��K��$LE(,6[�0��\ścIkߎ��1�V���#y��PXu��8n
�>��$!E�ώ�����KS7���q{��U%;��}E�Fإ��mU�-ɾM��\ҧ��0
�dn8�@c�Ked�X[�7���;8��w�/e]+�$	�|����˓��#���<S��[J7��ofv�;�\��"k��T�&4�$�-���ӭ��rO�%��!zw��2�������>�#�,x����e���)8��!�&z�c7����5:�r1���MǓ�8���"D���L��+=�DZ�?e����}��϶R�q.���\��&c}�U��gBT�rq��W��
�!Z�C?��������]o7��;�ٌ
;�r�����̮�j�X��F�/m�nߍ�x"���t�9���[�����M/�y�����S�5^���l��?�aU𞪃�i'5Q�������tӒ�v�\]��t�nȎ�7fE�ƨכS�W���'��d�,U7��XVG�ڜ��jX���m�m/3X'/yJ��jiH�h�Y�oUAV�-��g�$��t{z�\bTb�~���αZV0
 ��~!
�,��q��t-Y�yjK�0�nsCNߝcD���S��r��[����